// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Apr 6 2019 11:52:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_drone,
    uart_drone_data_rdy_debug,
    uart_commands_input_debug,
    ppm_output,
    uart_input_pc,
    uart_drone_input_debug,
    drone_frame_decoder_data_rdy_debug,
    clk_system);

    input uart_input_drone;
    output uart_drone_data_rdy_debug;
    output uart_commands_input_debug;
    output ppm_output;
    input uart_input_pc;
    output uart_drone_input_debug;
    output drone_frame_decoder_data_rdy_debug;
    input clk_system;

    wire N__29944;
    wire N__29943;
    wire N__29942;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29924;
    wire N__29923;
    wire N__29922;
    wire N__29915;
    wire N__29914;
    wire N__29913;
    wire N__29906;
    wire N__29905;
    wire N__29904;
    wire N__29897;
    wire N__29896;
    wire N__29895;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29860;
    wire N__29857;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29849;
    wire N__29848;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29840;
    wire N__29839;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29782;
    wire N__29779;
    wire N__29774;
    wire N__29771;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29745;
    wire N__29734;
    wire N__29731;
    wire N__29730;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29659;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29618;
    wire N__29615;
    wire N__29614;
    wire N__29613;
    wire N__29610;
    wire N__29601;
    wire N__29600;
    wire N__29595;
    wire N__29592;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29588;
    wire N__29587;
    wire N__29584;
    wire N__29579;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29558;
    wire N__29553;
    wire N__29548;
    wire N__29545;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29506;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29482;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29470;
    wire N__29469;
    wire N__29464;
    wire N__29463;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29442;
    wire N__29437;
    wire N__29430;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29387;
    wire N__29386;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29381;
    wire N__29380;
    wire N__29379;
    wire N__29378;
    wire N__29377;
    wire N__29376;
    wire N__29375;
    wire N__29374;
    wire N__29373;
    wire N__29372;
    wire N__29371;
    wire N__29370;
    wire N__29369;
    wire N__29368;
    wire N__29367;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29363;
    wire N__29362;
    wire N__29361;
    wire N__29360;
    wire N__29359;
    wire N__29358;
    wire N__29357;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29353;
    wire N__29352;
    wire N__29351;
    wire N__29350;
    wire N__29349;
    wire N__29348;
    wire N__29347;
    wire N__29346;
    wire N__29345;
    wire N__29344;
    wire N__29343;
    wire N__29342;
    wire N__29341;
    wire N__29340;
    wire N__29339;
    wire N__29338;
    wire N__29337;
    wire N__29336;
    wire N__29335;
    wire N__29334;
    wire N__29333;
    wire N__29332;
    wire N__29331;
    wire N__29330;
    wire N__29329;
    wire N__29328;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29324;
    wire N__29323;
    wire N__29322;
    wire N__29321;
    wire N__29320;
    wire N__29319;
    wire N__29318;
    wire N__29317;
    wire N__29316;
    wire N__29315;
    wire N__29314;
    wire N__29313;
    wire N__29312;
    wire N__29311;
    wire N__29310;
    wire N__29309;
    wire N__29308;
    wire N__29307;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29303;
    wire N__29302;
    wire N__29301;
    wire N__29300;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29296;
    wire N__29295;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29291;
    wire N__29290;
    wire N__29289;
    wire N__29288;
    wire N__29287;
    wire N__29286;
    wire N__29285;
    wire N__29284;
    wire N__29283;
    wire N__29282;
    wire N__29281;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29277;
    wire N__29276;
    wire N__29275;
    wire N__29274;
    wire N__29273;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29265;
    wire N__29264;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29260;
    wire N__29259;
    wire N__29258;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28977;
    wire N__28976;
    wire N__28973;
    wire N__28972;
    wire N__28969;
    wire N__28968;
    wire N__28965;
    wire N__28964;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28953;
    wire N__28952;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28948;
    wire N__28947;
    wire N__28946;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28927;
    wire N__28926;
    wire N__28925;
    wire N__28924;
    wire N__28921;
    wire N__28916;
    wire N__28913;
    wire N__28908;
    wire N__28905;
    wire N__28900;
    wire N__28897;
    wire N__28892;
    wire N__28889;
    wire N__28878;
    wire N__28867;
    wire N__28862;
    wire N__28855;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28796;
    wire N__28795;
    wire N__28794;
    wire N__28793;
    wire N__28792;
    wire N__28791;
    wire N__28790;
    wire N__28789;
    wire N__28788;
    wire N__28787;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28780;
    wire N__28779;
    wire N__28778;
    wire N__28777;
    wire N__28776;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28772;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28765;
    wire N__28764;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28760;
    wire N__28759;
    wire N__28758;
    wire N__28757;
    wire N__28756;
    wire N__28755;
    wire N__28754;
    wire N__28753;
    wire N__28752;
    wire N__28751;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28747;
    wire N__28746;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28742;
    wire N__28741;
    wire N__28740;
    wire N__28739;
    wire N__28738;
    wire N__28737;
    wire N__28736;
    wire N__28735;
    wire N__28734;
    wire N__28733;
    wire N__28732;
    wire N__28731;
    wire N__28730;
    wire N__28729;
    wire N__28728;
    wire N__28727;
    wire N__28726;
    wire N__28725;
    wire N__28724;
    wire N__28723;
    wire N__28722;
    wire N__28721;
    wire N__28720;
    wire N__28719;
    wire N__28718;
    wire N__28717;
    wire N__28716;
    wire N__28715;
    wire N__28714;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28362;
    wire N__28361;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28355;
    wire N__28354;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28316;
    wire N__28313;
    wire N__28312;
    wire N__28311;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28307;
    wire N__28302;
    wire N__28299;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28260;
    wire N__28251;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28230;
    wire N__28229;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28221;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28195;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28168;
    wire N__28165;
    wire N__28154;
    wire N__28151;
    wire N__28146;
    wire N__28143;
    wire N__28138;
    wire N__28135;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28116;
    wire N__28115;
    wire N__28114;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28106;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28065;
    wire N__28064;
    wire N__28063;
    wire N__28060;
    wire N__28053;
    wire N__28050;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28021;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27981;
    wire N__27978;
    wire N__27977;
    wire N__27976;
    wire N__27973;
    wire N__27972;
    wire N__27969;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27891;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27883;
    wire N__27880;
    wire N__27875;
    wire N__27872;
    wire N__27871;
    wire N__27870;
    wire N__27869;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27853;
    wire N__27852;
    wire N__27849;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27826;
    wire N__27825;
    wire N__27820;
    wire N__27813;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27774;
    wire N__27771;
    wire N__27770;
    wire N__27769;
    wire N__27768;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27737;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27719;
    wire N__27718;
    wire N__27715;
    wire N__27714;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27679;
    wire N__27674;
    wire N__27669;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27648;
    wire N__27647;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27632;
    wire N__27627;
    wire N__27624;
    wire N__27623;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27606;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27577;
    wire N__27572;
    wire N__27569;
    wire N__27564;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27544;
    wire N__27535;
    wire N__27532;
    wire N__27531;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27497;
    wire N__27490;
    wire N__27489;
    wire N__27488;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27470;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27429;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27388;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27343;
    wire N__27338;
    wire N__27337;
    wire N__27334;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27307;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27273;
    wire N__27272;
    wire N__27271;
    wire N__27270;
    wire N__27269;
    wire N__27268;
    wire N__27267;
    wire N__27266;
    wire N__27265;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27209;
    wire N__27208;
    wire N__27207;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27189;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27161;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27124;
    wire N__27119;
    wire N__27116;
    wire N__27111;
    wire N__27108;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27059;
    wire N__27052;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27031;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27019;
    wire N__27018;
    wire N__27017;
    wire N__27014;
    wire N__27009;
    wire N__27004;
    wire N__27003;
    wire N__27002;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26990;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26973;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26952;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26907;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26886;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26871;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26811;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26794;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26782;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26774;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26697;
    wire N__26696;
    wire N__26695;
    wire N__26694;
    wire N__26693;
    wire N__26692;
    wire N__26691;
    wire N__26688;
    wire N__26687;
    wire N__26686;
    wire N__26685;
    wire N__26684;
    wire N__26683;
    wire N__26680;
    wire N__26679;
    wire N__26676;
    wire N__26671;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26657;
    wire N__26648;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26632;
    wire N__26627;
    wire N__26626;
    wire N__26625;
    wire N__26624;
    wire N__26623;
    wire N__26622;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26585;
    wire N__26578;
    wire N__26575;
    wire N__26568;
    wire N__26565;
    wire N__26560;
    wire N__26557;
    wire N__26552;
    wire N__26537;
    wire N__26534;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26516;
    wire N__26511;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26496;
    wire N__26495;
    wire N__26494;
    wire N__26491;
    wire N__26484;
    wire N__26479;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26379;
    wire N__26378;
    wire N__26377;
    wire N__26376;
    wire N__26375;
    wire N__26374;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26341;
    wire N__26340;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26334;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26313;
    wire N__26310;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26287;
    wire N__26278;
    wire N__26275;
    wire N__26274;
    wire N__26273;
    wire N__26272;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26247;
    wire N__26244;
    wire N__26243;
    wire N__26240;
    wire N__26233;
    wire N__26228;
    wire N__26223;
    wire N__26220;
    wire N__26215;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26193;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26175;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26163;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26116;
    wire N__26113;
    wire N__26112;
    wire N__26111;
    wire N__26110;
    wire N__26109;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26095;
    wire N__26094;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26077;
    wire N__26074;
    wire N__26073;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26058;
    wire N__26053;
    wire N__26048;
    wire N__26043;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25864;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25856;
    wire N__25853;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25811;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25794;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25767;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25746;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25683;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25659;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25638;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25617;
    wire N__25616;
    wire N__25613;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25598;
    wire N__25595;
    wire N__25588;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25579;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25567;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25552;
    wire N__25549;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25525;
    wire N__25524;
    wire N__25523;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25502;
    wire N__25499;
    wire N__25494;
    wire N__25489;
    wire N__25488;
    wire N__25483;
    wire N__25480;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25250;
    wire N__25243;
    wire N__25242;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25210;
    wire N__25209;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25155;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25066;
    wire N__25065;
    wire N__25062;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25050;
    wire N__25043;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25025;
    wire N__25020;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25005;
    wire N__25002;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24963;
    wire N__24962;
    wire N__24961;
    wire N__24960;
    wire N__24959;
    wire N__24956;
    wire N__24955;
    wire N__24954;
    wire N__24951;
    wire N__24950;
    wire N__24949;
    wire N__24948;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24913;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24904;
    wire N__24891;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24869;
    wire N__24868;
    wire N__24867;
    wire N__24866;
    wire N__24865;
    wire N__24864;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24843;
    wire N__24842;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24823;
    wire N__24820;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24779;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24754;
    wire N__24751;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24727;
    wire N__24714;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24685;
    wire N__24676;
    wire N__24675;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24660;
    wire N__24655;
    wire N__24652;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24634;
    wire N__24633;
    wire N__24628;
    wire N__24625;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24451;
    wire N__24448;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24393;
    wire N__24390;
    wire N__24385;
    wire N__24382;
    wire N__24381;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24333;
    wire N__24328;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24138;
    wire N__24133;
    wire N__24130;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24099;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24060;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24018;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23973;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23934;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23877;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23850;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23835;
    wire N__23832;
    wire N__23827;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23823;
    wire N__23822;
    wire N__23821;
    wire N__23814;
    wire N__23813;
    wire N__23812;
    wire N__23811;
    wire N__23810;
    wire N__23809;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23799;
    wire N__23798;
    wire N__23797;
    wire N__23796;
    wire N__23795;
    wire N__23794;
    wire N__23789;
    wire N__23788;
    wire N__23787;
    wire N__23786;
    wire N__23785;
    wire N__23784;
    wire N__23781;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23768;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23762;
    wire N__23761;
    wire N__23760;
    wire N__23757;
    wire N__23756;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23750;
    wire N__23749;
    wire N__23748;
    wire N__23745;
    wire N__23744;
    wire N__23737;
    wire N__23734;
    wire N__23733;
    wire N__23732;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23724;
    wire N__23717;
    wire N__23714;
    wire N__23703;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23687;
    wire N__23676;
    wire N__23669;
    wire N__23658;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23652;
    wire N__23651;
    wire N__23650;
    wire N__23647;
    wire N__23638;
    wire N__23635;
    wire N__23630;
    wire N__23629;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23605;
    wire N__23602;
    wire N__23601;
    wire N__23588;
    wire N__23575;
    wire N__23570;
    wire N__23561;
    wire N__23560;
    wire N__23559;
    wire N__23558;
    wire N__23557;
    wire N__23556;
    wire N__23553;
    wire N__23552;
    wire N__23549;
    wire N__23544;
    wire N__23535;
    wire N__23532;
    wire N__23527;
    wire N__23518;
    wire N__23509;
    wire N__23502;
    wire N__23485;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23470;
    wire N__23469;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23449;
    wire N__23448;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23404;
    wire N__23403;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23386;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23340;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23313;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23286;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23253;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23136;
    wire N__23135;
    wire N__23128;
    wire N__23127;
    wire N__23126;
    wire N__23125;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23101;
    wire N__23098;
    wire N__23097;
    wire N__23096;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23088;
    wire N__23083;
    wire N__23072;
    wire N__23069;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23053;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23015;
    wire N__23010;
    wire N__23007;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22939;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22914;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22897;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22876;
    wire N__22875;
    wire N__22874;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22858;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22851;
    wire N__22850;
    wire N__22849;
    wire N__22848;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22828;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22815;
    wire N__22810;
    wire N__22803;
    wire N__22800;
    wire N__22799;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22772;
    wire N__22769;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22758;
    wire N__22749;
    wire N__22746;
    wire N__22741;
    wire N__22738;
    wire N__22733;
    wire N__22730;
    wire N__22717;
    wire N__22714;
    wire N__22713;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22689;
    wire N__22684;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22662;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22591;
    wire N__22590;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22570;
    wire N__22569;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22338;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22309;
    wire N__22306;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22237;
    wire N__22232;
    wire N__22231;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22207;
    wire N__22204;
    wire N__22199;
    wire N__22194;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22173;
    wire N__22170;
    wire N__22169;
    wire N__22166;
    wire N__22165;
    wire N__22162;
    wire N__22155;
    wire N__22150;
    wire N__22149;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22117;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22102;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22084;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22060;
    wire N__22057;
    wire N__22056;
    wire N__22055;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22051;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22035;
    wire N__22030;
    wire N__22021;
    wire N__22020;
    wire N__22019;
    wire N__22016;
    wire N__22015;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21991;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21962;
    wire N__21959;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21928;
    wire N__21923;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21900;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21796;
    wire N__21795;
    wire N__21794;
    wire N__21793;
    wire N__21792;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21772;
    wire N__21765;
    wire N__21760;
    wire N__21757;
    wire N__21756;
    wire N__21755;
    wire N__21754;
    wire N__21751;
    wire N__21750;
    wire N__21749;
    wire N__21748;
    wire N__21747;
    wire N__21746;
    wire N__21743;
    wire N__21742;
    wire N__21741;
    wire N__21740;
    wire N__21739;
    wire N__21738;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21716;
    wire N__21713;
    wire N__21706;
    wire N__21701;
    wire N__21694;
    wire N__21691;
    wire N__21686;
    wire N__21683;
    wire N__21676;
    wire N__21673;
    wire N__21668;
    wire N__21665;
    wire N__21660;
    wire N__21655;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21619;
    wire N__21616;
    wire N__21611;
    wire N__21608;
    wire N__21603;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21565;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21557;
    wire N__21554;
    wire N__21553;
    wire N__21552;
    wire N__21547;
    wire N__21544;
    wire N__21539;
    wire N__21532;
    wire N__21531;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21487;
    wire N__21484;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21339;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21310;
    wire N__21309;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21255;
    wire N__21254;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21231;
    wire N__21230;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21191;
    wire N__21190;
    wire N__21187;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21147;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21132;
    wire N__21127;
    wire N__21124;
    wire N__21123;
    wire N__21122;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21106;
    wire N__21103;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21089;
    wire N__21084;
    wire N__21081;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21043;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20985;
    wire N__20980;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20962;
    wire N__20961;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20957;
    wire N__20952;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20944;
    wire N__20939;
    wire N__20938;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20861;
    wire N__20856;
    wire N__20849;
    wire N__20844;
    wire N__20839;
    wire N__20828;
    wire N__20825;
    wire N__20820;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20794;
    wire N__20793;
    wire N__20792;
    wire N__20791;
    wire N__20790;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20784;
    wire N__20783;
    wire N__20782;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20778;
    wire N__20777;
    wire N__20776;
    wire N__20775;
    wire N__20774;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20760;
    wire N__20759;
    wire N__20756;
    wire N__20747;
    wire N__20738;
    wire N__20731;
    wire N__20722;
    wire N__20715;
    wire N__20714;
    wire N__20713;
    wire N__20710;
    wire N__20703;
    wire N__20702;
    wire N__20699;
    wire N__20694;
    wire N__20693;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20668;
    wire N__20667;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20652;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20630;
    wire N__20619;
    wire N__20614;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20571;
    wire N__20570;
    wire N__20569;
    wire N__20568;
    wire N__20565;
    wire N__20560;
    wire N__20559;
    wire N__20556;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20546;
    wire N__20545;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20521;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20478;
    wire N__20475;
    wire N__20470;
    wire N__20467;
    wire N__20462;
    wire N__20455;
    wire N__20440;
    wire N__20439;
    wire N__20438;
    wire N__20435;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20412;
    wire N__20409;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20369;
    wire N__20366;
    wire N__20365;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20355;
    wire N__20352;
    wire N__20351;
    wire N__20346;
    wire N__20345;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20327;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20302;
    wire N__20293;
    wire N__20290;
    wire N__20285;
    wire N__20282;
    wire N__20277;
    wire N__20266;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20245;
    wire N__20244;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20229;
    wire N__20224;
    wire N__20221;
    wire N__20220;
    wire N__20219;
    wire N__20218;
    wire N__20215;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20150;
    wire N__20147;
    wire N__20142;
    wire N__20137;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20091;
    wire N__20088;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20073;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20063;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20041;
    wire N__20040;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20010;
    wire N__20009;
    wire N__20006;
    wire N__20005;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19988;
    wire N__19985;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19938;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19914;
    wire N__19913;
    wire N__19910;
    wire N__19905;
    wire N__19900;
    wire N__19897;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19817;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19801;
    wire N__19798;
    wire N__19797;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19725;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19710;
    wire N__19709;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19638;
    wire N__19637;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19615;
    wire N__19614;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19558;
    wire N__19557;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19536;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19513;
    wire N__19512;
    wire N__19511;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19505;
    wire N__19496;
    wire N__19493;
    wire N__19486;
    wire N__19483;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19466;
    wire N__19465;
    wire N__19458;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19438;
    wire N__19435;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19429;
    wire N__19428;
    wire N__19425;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19290;
    wire N__19289;
    wire N__19286;
    wire N__19279;
    wire N__19278;
    wire N__19275;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19233;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19180;
    wire N__19177;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19155;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19094;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19044;
    wire N__19039;
    wire N__19038;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19026;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18993;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18981;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18950;
    wire N__18947;
    wire N__18940;
    wire N__18937;
    wire N__18936;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18902;
    wire N__18895;
    wire N__18888;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18693;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18675;
    wire N__18670;
    wire N__18667;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18655;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18630;
    wire N__18629;
    wire N__18626;
    wire N__18621;
    wire N__18616;
    wire N__18613;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18605;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18571;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18563;
    wire N__18562;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18547;
    wire N__18542;
    wire N__18539;
    wire N__18538;
    wire N__18537;
    wire N__18532;
    wire N__18529;
    wire N__18524;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18486;
    wire N__18485;
    wire N__18484;
    wire N__18481;
    wire N__18474;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18457;
    wire N__18450;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18405;
    wire N__18404;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18244;
    wire N__18243;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18231;
    wire N__18228;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18211;
    wire N__18210;
    wire N__18209;
    wire N__18206;
    wire N__18205;
    wire N__18204;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18187;
    wire N__18184;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18166;
    wire N__18161;
    wire N__18158;
    wire N__18153;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18111;
    wire N__18110;
    wire N__18109;
    wire N__18108;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18094;
    wire N__18091;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18072;
    wire N__18067;
    wire N__18064;
    wire N__18063;
    wire N__18062;
    wire N__18055;
    wire N__18050;
    wire N__18049;
    wire N__18046;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18011;
    wire N__18010;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17988;
    wire N__17985;
    wire N__17980;
    wire N__17977;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17930;
    wire N__17923;
    wire N__17920;
    wire N__17919;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17904;
    wire N__17899;
    wire N__17898;
    wire N__17895;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17859;
    wire N__17858;
    wire N__17857;
    wire N__17852;
    wire N__17847;
    wire N__17844;
    wire N__17843;
    wire N__17842;
    wire N__17839;
    wire N__17836;
    wire N__17831;
    wire N__17824;
    wire N__17823;
    wire N__17820;
    wire N__17819;
    wire N__17818;
    wire N__17815;
    wire N__17810;
    wire N__17809;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17801;
    wire N__17798;
    wire N__17793;
    wire N__17788;
    wire N__17785;
    wire N__17780;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17569;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17536;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17516;
    wire N__17515;
    wire N__17510;
    wire N__17505;
    wire N__17502;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17480;
    wire N__17475;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17439;
    wire N__17438;
    wire N__17433;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17416;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17398;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17390;
    wire N__17389;
    wire N__17388;
    wire N__17387;
    wire N__17386;
    wire N__17381;
    wire N__17372;
    wire N__17371;
    wire N__17370;
    wire N__17367;
    wire N__17362;
    wire N__17357;
    wire N__17350;
    wire N__17349;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17341;
    wire N__17340;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17326;
    wire N__17323;
    wire N__17322;
    wire N__17321;
    wire N__17320;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17300;
    wire N__17295;
    wire N__17284;
    wire N__17283;
    wire N__17282;
    wire N__17281;
    wire N__17280;
    wire N__17279;
    wire N__17278;
    wire N__17277;
    wire N__17274;
    wire N__17273;
    wire N__17270;
    wire N__17265;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17249;
    wire N__17248;
    wire N__17245;
    wire N__17240;
    wire N__17235;
    wire N__17230;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17137;
    wire N__17136;
    wire N__17135;
    wire N__17132;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17116;
    wire N__17113;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17074;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17059;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17037;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17026;
    wire N__17025;
    wire N__17024;
    wire N__17019;
    wire N__17016;
    wire N__17011;
    wire N__17008;
    wire N__16999;
    wire N__16996;
    wire N__16995;
    wire N__16994;
    wire N__16993;
    wire N__16992;
    wire N__16991;
    wire N__16988;
    wire N__16987;
    wire N__16982;
    wire N__16975;
    wire N__16972;
    wire N__16971;
    wire N__16968;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16952;
    wire N__16945;
    wire N__16944;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16894;
    wire N__16893;
    wire N__16892;
    wire N__16891;
    wire N__16882;
    wire N__16879;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16837;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16825;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16778;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16766;
    wire N__16761;
    wire N__16756;
    wire N__16753;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16741;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16722;
    wire N__16719;
    wire N__16714;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16699;
    wire N__16696;
    wire N__16691;
    wire N__16688;
    wire N__16681;
    wire N__16678;
    wire N__16677;
    wire N__16676;
    wire N__16673;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16665;
    wire N__16664;
    wire N__16663;
    wire N__16654;
    wire N__16651;
    wire N__16646;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16596;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16458;
    wire N__16457;
    wire N__16452;
    wire N__16449;
    wire N__16448;
    wire N__16447;
    wire N__16444;
    wire N__16443;
    wire N__16442;
    wire N__16441;
    wire N__16440;
    wire N__16437;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16419;
    wire N__16414;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16319;
    wire N__16314;
    wire N__16313;
    wire N__16312;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16295;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16240;
    wire N__16239;
    wire N__16238;
    wire N__16235;
    wire N__16230;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16194;
    wire N__16193;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16149;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16128;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16065;
    wire N__16062;
    wire N__16061;
    wire N__16060;
    wire N__16057;
    wire N__16056;
    wire N__16055;
    wire N__16054;
    wire N__16047;
    wire N__16044;
    wire N__16043;
    wire N__16042;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16020;
    wire N__16015;
    wire N__16012;
    wire N__16007;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15991;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15981;
    wire N__15978;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15970;
    wire N__15969;
    wire N__15966;
    wire N__15965;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15950;
    wire N__15947;
    wire N__15942;
    wire N__15937;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15890;
    wire N__15883;
    wire N__15882;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15865;
    wire N__15864;
    wire N__15863;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15850;
    wire N__15849;
    wire N__15848;
    wire N__15847;
    wire N__15846;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15833;
    wire N__15830;
    wire N__15825;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15801;
    wire N__15798;
    wire N__15793;
    wire N__15772;
    wire N__15771;
    wire N__15770;
    wire N__15769;
    wire N__15766;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15758;
    wire N__15757;
    wire N__15754;
    wire N__15747;
    wire N__15746;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15709;
    wire N__15706;
    wire N__15701;
    wire N__15688;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15597;
    wire N__15596;
    wire N__15593;
    wire N__15588;
    wire N__15583;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15568;
    wire N__15567;
    wire N__15566;
    wire N__15563;
    wire N__15558;
    wire N__15553;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15483;
    wire N__15480;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15465;
    wire N__15462;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15436;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15424;
    wire N__15421;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15370;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15313;
    wire N__15310;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15288;
    wire N__15287;
    wire N__15284;
    wire N__15283;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15264;
    wire N__15261;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15253;
    wire N__15252;
    wire N__15249;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15234;
    wire N__15233;
    wire N__15230;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15175;
    wire N__15170;
    wire N__15169;
    wire N__15166;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15136;
    wire N__15133;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15108;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15091;
    wire N__15090;
    wire N__15089;
    wire N__15088;
    wire N__15087;
    wire N__15086;
    wire N__15085;
    wire N__15084;
    wire N__15083;
    wire N__15082;
    wire N__15079;
    wire N__15070;
    wire N__15067;
    wire N__15062;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15044;
    wire N__15041;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15025;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15008;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14993;
    wire N__14990;
    wire N__14985;
    wire N__14980;
    wire N__14977;
    wire N__14972;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14925;
    wire N__14920;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14910;
    wire N__14905;
    wire N__14904;
    wire N__14901;
    wire N__14896;
    wire N__14893;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14815;
    wire N__14814;
    wire N__14811;
    wire N__14810;
    wire N__14809;
    wire N__14808;
    wire N__14805;
    wire N__14800;
    wire N__14799;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14773;
    wire N__14770;
    wire N__14765;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14674;
    wire N__14671;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14652;
    wire N__14649;
    wire N__14646;
    wire N__14641;
    wire N__14638;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14580;
    wire N__14577;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14560;
    wire N__14559;
    wire N__14558;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14546;
    wire N__14543;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14466;
    wire N__14463;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14445;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14379;
    wire N__14378;
    wire N__14375;
    wire N__14370;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14187;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13995;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13963;
    wire N__13962;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13899;
    wire N__13898;
    wire N__13895;
    wire N__13890;
    wire N__13885;
    wire N__13882;
    wire N__13881;
    wire N__13880;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13866;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13823;
    wire N__13818;
    wire N__13815;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13803;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13707;
    wire N__13704;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13689;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13663;
    wire N__13660;
    wire N__13651;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13643;
    wire N__13640;
    wire N__13635;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13620;
    wire N__13619;
    wire N__13616;
    wire N__13611;
    wire N__13608;
    wire N__13603;
    wire N__13602;
    wire N__13599;
    wire N__13598;
    wire N__13597;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13572;
    wire N__13569;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13534;
    wire N__13533;
    wire N__13532;
    wire N__13527;
    wire N__13526;
    wire N__13525;
    wire N__13522;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13501;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13483;
    wire N__13482;
    wire N__13479;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13461;
    wire N__13460;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13430;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13420;
    wire N__13415;
    wire N__13410;
    wire N__13405;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13386;
    wire N__13385;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13375;
    wire N__13372;
    wire N__13367;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13335;
    wire N__13332;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13288;
    wire N__13285;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13273;
    wire N__13270;
    wire N__13269;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13257;
    wire N__13254;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13221;
    wire N__13220;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13174;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13134;
    wire N__13133;
    wire N__13130;
    wire N__13129;
    wire N__13128;
    wire N__13125;
    wire N__13124;
    wire N__13123;
    wire N__13118;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13104;
    wire N__13101;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13051;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13041;
    wire N__13040;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12975;
    wire N__12974;
    wire N__12973;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12867;
    wire N__12866;
    wire N__12865;
    wire N__12860;
    wire N__12855;
    wire N__12850;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12842;
    wire N__12839;
    wire N__12834;
    wire N__12829;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12821;
    wire N__12818;
    wire N__12813;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12790;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12778;
    wire N__12775;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12760;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12719;
    wire N__12714;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12289;
    wire N__12288;
    wire N__12287;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12198;
    wire N__12197;
    wire N__12196;
    wire N__12195;
    wire N__12188;
    wire N__12183;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12144;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12127;
    wire N__12124;
    wire N__12123;
    wire N__12120;
    wire N__12119;
    wire N__12116;
    wire N__12111;
    wire N__12106;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12073;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12034;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12019;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12001;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11971;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11959;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11947;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11935;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11920;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11908;
    wire N__11907;
    wire N__11906;
    wire N__11903;
    wire N__11898;
    wire N__11893;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11881;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11861;
    wire N__11856;
    wire N__11851;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11806;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11785;
    wire N__11782;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11767;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11604;
    wire N__11601;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11560;
    wire N__11557;
    wire N__11556;
    wire N__11555;
    wire N__11552;
    wire N__11547;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11511;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire VCCG0;
    wire GNDG0;
    wire \pid_alt.O_17 ;
    wire \pid_alt.O_6 ;
    wire \pid_alt.O_7 ;
    wire \pid_alt.O_10 ;
    wire \pid_alt.O_16 ;
    wire \pid_alt.O_12 ;
    wire \pid_alt.O_11 ;
    wire \pid_alt.O_13 ;
    wire \pid_alt.O_18 ;
    wire \pid_alt.O_14 ;
    wire \pid_alt.O_4 ;
    wire \pid_alt.O_5 ;
    wire \pid_alt.O_9 ;
    wire \pid_alt.O_15 ;
    wire \pid_alt.O_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_1_13_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire bfn_1_14_0_;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire bfn_1_15_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_1_16_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire drone_altitude_i_10;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire drone_altitude_i_11;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire drone_altitude_12;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire drone_altitude_13;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire drone_altitude_15;
    wire drone_altitude_i_7;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ;
    wire bfn_1_28_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire bfn_1_29_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_1_30_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire alt_kp_0;
    wire alt_kp_2;
    wire alt_kp_1;
    wire \pid_alt.source_p_enZ0 ;
    wire alt_kp_3;
    wire alt_kp_6;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4 ;
    wire \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lto13_1 ;
    wire \dron_frame_decoder_1.WDT10lt14_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.WDT10lt14_0_cascade_ ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire drone_altitude_0;
    wire \pid_alt.drone_altitude_i_0 ;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire drone_altitude_i_4;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire drone_altitude_i_5;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire drone_altitude_i_6;
    wire drone_altitude_1;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire \dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_ ;
    wire \dron_frame_decoder_1.source_Altitude8lt7_0_cascade_ ;
    wire drone_altitude_2;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire \dron_frame_decoder_1.source_Altitude8lt7_0 ;
    wire drone_altitude_3;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire alt_command_3;
    wire alt_command_1;
    wire \Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire alt_command_0;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire alt_command_2;
    wire \Commands_frame_decoder.source_CH1data8lt7_0 ;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire drone_altitude_i_8;
    wire drone_altitude_i_9;
    wire drone_altitude_14;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire bfn_2_19_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire throttle_command_3;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire throttle_command_6;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_2_20_0_;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire throttle_command_14;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire throttle_command_1;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_command_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire throttle_command_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire throttle_command_4;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire throttle_command_5;
    wire throttle_command_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_command_7;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_58_d_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_command_2;
    wire \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ;
    wire throttle_command_0;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.N_299 ;
    wire alt_kp_7;
    wire alt_kp_5;
    wire \dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_a3_0_3_1 ;
    wire \dron_frame_decoder_1.state_ns_0_a3_0_3_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \dron_frame_decoder_1.N_217_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \dron_frame_decoder_1.N_219 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_ ;
    wire \dron_frame_decoder_1.N_239 ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_2_0 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ;
    wire \dron_frame_decoder_1.N_243 ;
    wire alt_command_4;
    wire alt_command_5;
    wire alt_command_6;
    wire alt_command_7;
    wire \dron_frame_decoder_1.N_238_0 ;
    wire \dron_frame_decoder_1.N_237 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_0_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_ ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ;
    wire \dron_frame_decoder_1.N_230_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire uart_drone_data_rdy_debug_c;
    wire drone_frame_decoder_data_rdy_debug_c;
    wire \uart_pc.N_152_cascade_ ;
    wire \uart_pc.CO0_cascade_ ;
    wire \uart_pc.un1_state_7_0 ;
    wire throttle_command_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire throttle_command_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire throttle_command_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.N_303_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4 ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5 ;
    wire \ppm_encoder_1.throttle_RNIN3352Z0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire bfn_3_25_0_;
    wire \ppm_encoder_1.throttle_RNIALN65Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.throttle_RNI5V123Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.throttle_RNI82223Z0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.throttle_RNIJII96Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.throttle_RNIONI96Z0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire bfn_3_26_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.throttle_RNITSI96Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_3_27_0_;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.N_295 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_13_cascade_ ;
    wire \reset_module_System.reset6_3 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire bfn_4_12_0_;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_4_13_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_4_14_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_11 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_3_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.state_1_ns_0_a4_0_0_2 ;
    wire uart_drone_data_0;
    wire uart_drone_data_1;
    wire uart_drone_data_2;
    wire uart_drone_data_3;
    wire uart_drone_data_4;
    wire uart_drone_data_5;
    wire uart_drone_data_6;
    wire uart_drone_data_7;
    wire \uart_drone.state_1_sqmuxa_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_4_18_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire bfn_4_19_0_;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.WDT8lto13_1_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.N_300_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ;
    wire \ppm_encoder_1.N_139_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14 ;
    wire \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10 ;
    wire \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ;
    wire \ppm_encoder_1.N_318 ;
    wire \ppm_encoder_1.N_226 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire bfn_4_29_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_4_30_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.reset6_14 ;
    wire \Commands_frame_decoder.state_1_RNIVM1OZ0Z_6 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.state_1Z0Z_5 ;
    wire \Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0 ;
    wire \Commands_frame_decoder.state_1_ns_0_a4_0_3_2 ;
    wire \Commands_frame_decoder.N_323_cascade_ ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \Commands_frame_decoder.state_1Z0Z_2 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ;
    wire \Commands_frame_decoder.state_1Z0Z_3 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.state_1Z0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_drone.state_1_sqmuxa ;
    wire \Commands_frame_decoder.un1_state49_iZ0 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire \uart_drone.N_143_cascade_ ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire bfn_5_19_0_;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.N_302_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.N_296_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ;
    wire \ppm_encoder_1.N_237 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.N_237_cascade_ ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \uart_pc_sync.aux_2__0__0_0 ;
    wire \uart_pc_sync.aux_3__0__0_0 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire uart_commands_input_debug_c;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_144_1_cascade_ ;
    wire \uart_pc.state_1_sqmuxa ;
    wire \uart_pc.N_145 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.un1_state_2_0 ;
    wire bfn_7_19_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_7_20_0_;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.N_305_cascade_ ;
    wire \ppm_encoder_1.N_298 ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.N_304_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.N_319_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.N_590_i ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_7_28_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_7_29_0_;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_7_30_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_168_g ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0_Z0Z_0 ;
    wire \uart_drone_sync.aux_1__0_Z0Z_0 ;
    wire \uart_drone_sync.aux_2__0_Z0Z_0 ;
    wire \uart_drone_sync.aux_3__0_Z0Z_0 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire frame_decoder_CH2data_7;
    wire bfn_8_13_0_;
    wire frame_decoder_CH2data_1;
    wire \scaler_2.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH2data_2;
    wire \scaler_2.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH2data_3;
    wire frame_decoder_OFF2data_3;
    wire \scaler_2.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH2data_4;
    wire \scaler_2.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH2data_5;
    wire frame_decoder_OFF2data_5;
    wire \scaler_2.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH2data_6;
    wire frame_decoder_OFF2data_6;
    wire \scaler_2.un3_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_axb_7 ;
    wire \scaler_2.un3_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_7 ;
    wire \scaler_2.N_521_i_l_ofxZ0 ;
    wire bfn_8_14_0_;
    wire \scaler_2.un3_source_data_0_cry_8 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.un1_state_2_0 ;
    wire uart_drone_input_debug_c;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_145 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.N_144_1 ;
    wire \Commands_frame_decoder.state_1_RNO_4Z0Z_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire bfn_8_18_0_;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.stateZ0Z_4 ;
    wire bfn_8_19_0_;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire bfn_8_20_0_;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.N_301 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ;
    wire \ppm_encoder_1.N_144_17 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \ppm_encoder_1.N_144_17_cascade_ ;
    wire \ppm_encoder_1.N_144 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.N_590_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_158_d ;
    wire \ppm_encoder_1.PPM_STATE_58_d ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0__0_0 ;
    wire \uart_pc_sync.aux_1__0__0_0 ;
    wire frame_decoder_OFF2data_7;
    wire frame_decoder_OFF2data_1;
    wire frame_decoder_OFF2data_4;
    wire frame_decoder_OFF2data_2;
    wire bfn_9_13_0_;
    wire scaler_2_data_6;
    wire \scaler_2.un2_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_1_c_RNI14IK ;
    wire scaler_2_data_7;
    wire \scaler_2.un2_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_2_c_RNI48JK ;
    wire scaler_2_data_8;
    wire \scaler_2.un2_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ;
    wire scaler_2_data_9;
    wire \scaler_2.un2_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ;
    wire scaler_2_data_10;
    wire \scaler_2.un2_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ;
    wire scaler_2_data_11;
    wire \scaler_2.un2_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ;
    wire scaler_2_data_12;
    wire \scaler_2.un2_source_data_0_cry_7 ;
    wire \scaler_2.un2_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ;
    wire \scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ;
    wire scaler_2_data_13;
    wire bfn_9_14_0_;
    wire \scaler_2.un2_source_data_0_cry_9 ;
    wire scaler_2_data_14;
    wire scaler_2_data_5;
    wire scaler_3_data_5;
    wire scaler_4_data_5;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire scaler_2_data_4;
    wire scaler_3_data_4;
    wire scaler_4_data_4;
    wire \Commands_frame_decoder.N_282_0_cascade_ ;
    wire \Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1 ;
    wire \Commands_frame_decoder.source_CH1data8lto7Z0Z_1 ;
    wire \Commands_frame_decoder.N_319_cascade_ ;
    wire \Commands_frame_decoder.N_318 ;
    wire \Commands_frame_decoder.N_282_0 ;
    wire \Commands_frame_decoder.state_1_RNO_1Z0Z_0 ;
    wire \Commands_frame_decoder.state_1_ns_i_0_0_cascade_ ;
    wire \Commands_frame_decoder.state_1Z0Z_0 ;
    wire \Commands_frame_decoder.N_323 ;
    wire \Commands_frame_decoder.state_1_ns_0_a4_0_2_1 ;
    wire \Commands_frame_decoder.state_1Z0Z_1 ;
    wire bfn_9_19_0_;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire bfn_9_20_0_;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire pid_altitude_dv;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire frame_decoder_CH4data_7;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ;
    wire \scaler_2.un2_source_data_0 ;
    wire frame_decoder_OFF2data_0;
    wire frame_decoder_CH2data_0;
    wire \scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire frame_decoder_OFF4data_7;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNO_1 ;
    wire bfn_10_15_0_;
    wire scaler_4_data_6;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire scaler_4_data_7;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire scaler_4_data_8;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire scaler_4_data_9;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire scaler_4_data_10;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire scaler_4_data_11;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire scaler_4_data_12;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire scaler_4_data_13;
    wire bfn_10_16_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire \Commands_frame_decoder.state_1Z0Z_6 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.N_152 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \Commands_frame_decoder.state_1Z0Z_7 ;
    wire frame_decoder_OFF4data_0;
    wire bfn_11_14_0_;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un2_source_data_0 ;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire \scaler_4.N_545_i_l_ofxZ0 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire bfn_11_15_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire bfn_11_16_0_;
    wire scaler_3_data_6;
    wire \scaler_3.un2_source_data_0_cry_1 ;
    wire scaler_3_data_7;
    wire \scaler_3.un2_source_data_0_cry_2 ;
    wire scaler_3_data_8;
    wire \scaler_3.un2_source_data_0_cry_3 ;
    wire scaler_3_data_9;
    wire \scaler_3.un2_source_data_0_cry_4 ;
    wire scaler_3_data_10;
    wire \scaler_3.un2_source_data_0_cry_5 ;
    wire scaler_3_data_11;
    wire \scaler_3.un2_source_data_0_cry_6 ;
    wire scaler_3_data_12;
    wire \scaler_3.un2_source_data_0_cry_7 ;
    wire \scaler_3.un2_source_data_0_cry_8 ;
    wire scaler_3_data_13;
    wire bfn_11_17_0_;
    wire \scaler_3.un2_source_data_0_cry_9 ;
    wire scaler_3_data_14;
    wire pc_frame_decoder_dv_0_g;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \Commands_frame_decoder.state_1Z0Z_10 ;
    wire \Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_ ;
    wire \Commands_frame_decoder.N_292 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.CO0 ;
    wire bfn_11_19_0_;
    wire \Commands_frame_decoder.count8_axb_1 ;
    wire \Commands_frame_decoder.count8_cry_0 ;
    wire \Commands_frame_decoder.count_i_2 ;
    wire \Commands_frame_decoder.count8_cry_1 ;
    wire \Commands_frame_decoder.count8 ;
    wire \Commands_frame_decoder.count8_THRU_CO ;
    wire reset_system;
    wire \Commands_frame_decoder.count8_THRU_CO_cascade_ ;
    wire \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_ ;
    wire \Commands_frame_decoder.countZ0Z_2 ;
    wire \Commands_frame_decoder.CO0 ;
    wire \Commands_frame_decoder.CO0_cascade_ ;
    wire \Commands_frame_decoder.countZ0Z_1 ;
    wire pc_frame_decoder_dv_0;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_CH4data_0;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire bfn_12_15_0_;
    wire \scaler_3.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH3data_2;
    wire \scaler_3.un3_source_data_0_cry_1_c_RNI44VK ;
    wire \scaler_3.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH3data_3;
    wire \scaler_3.un3_source_data_0_cry_2_c_RNI780L ;
    wire \scaler_3.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH3data_4;
    wire \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ;
    wire \scaler_3.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH3data_5;
    wire \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ;
    wire \scaler_3.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH3data_6;
    wire \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ;
    wire \scaler_3.un3_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_6_c_RNILUAN ;
    wire \scaler_3.un3_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_7 ;
    wire \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ;
    wire bfn_12_16_0_;
    wire \scaler_3.un3_source_data_0_cry_8 ;
    wire \scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ;
    wire \scaler_3.N_533_i_l_ofxZ0 ;
    wire \scaler_3.un2_source_data_0 ;
    wire frame_decoder_CH3data_0;
    wire \scaler_3.un2_source_data_0_cry_1_c_RNO_0 ;
    wire \scaler_3.un3_source_data_0_axb_7 ;
    wire frame_decoder_CH3data_1;
    wire frame_decoder_CH3data_7;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire pc_frame_decoder_dv;
    wire CONSTANT_ONE_NET;
    wire \Commands_frame_decoder.count8_0_i ;
    wire \Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0 ;
    wire \Commands_frame_decoder.state_1_ns_i_a4_2_0_0 ;
    wire \Commands_frame_decoder.count8_0 ;
    wire frame_decoder_OFF4data_3;
    wire frame_decoder_OFF4data_6;
    wire uart_pc_data_2;
    wire frame_decoder_OFF3data_2;
    wire uart_pc_data_6;
    wire frame_decoder_OFF3data_6;
    wire uart_pc_data_3;
    wire frame_decoder_OFF3data_3;
    wire uart_pc_data_4;
    wire frame_decoder_OFF3data_4;
    wire uart_pc_data_5;
    wire frame_decoder_OFF3data_5;
    wire uart_pc_data_1;
    wire frame_decoder_OFF3data_1;
    wire uart_pc_data_7;
    wire frame_decoder_OFF3data_7;
    wire uart_pc_data_0;
    wire frame_decoder_OFF3data_0;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa ;
    wire \Commands_frame_decoder.state_1Z0Z_8 ;
    wire \Commands_frame_decoder.N_316 ;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa ;
    wire \Commands_frame_decoder.state_1Z0Z_9 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire reset_system_g;

    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__27295),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__27264),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__11359,N__11377,N__11392,N__11407,N__11422,N__11437,N__11227,N__11242,N__11257,N__11272,N__11284,N__11299,N__11314,N__11329,N__11188,N__12091}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__13195,N__12018,N__13174,N__16630,N__12037,N__11806,N__11785,N__11824}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,\pid_alt.O_18 ,\pid_alt.O_17 ,\pid_alt.O_16 ,\pid_alt.O_15 ,\pid_alt.O_14 ,\pid_alt.O_13 ,\pid_alt.O_12 ,\pid_alt.O_11 ,\pid_alt.O_10 ,\pid_alt.O_9 ,\pid_alt.O_8 ,\pid_alt.O_7 ,\pid_alt.O_6 ,\pid_alt.O_5 ,\pid_alt.O_4 ,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56}));
    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__29942),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__29944),
            .DIN(N__29943),
            .DOUT(N__29942),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__29944),
            .PADOUT(N__29943),
            .PADIN(N__29942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__29933),
            .DIN(N__29932),
            .DOUT(N__29931),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__29933),
            .PADOUT(N__29932),
            .PADIN(N__29931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__29924),
            .DIN(N__29923),
            .DOUT(N__29922),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__29924),
            .PADOUT(N__29923),
            .PADIN(N__29922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__29915),
            .DIN(N__29914),
            .DOUT(N__29913),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__29915),
            .PADOUT(N__29914),
            .PADIN(N__29913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15523),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_drone_data_rdy_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_drone_data_rdy_debug_obuf_iopad (
            .OE(N__29906),
            .DIN(N__29905),
            .DOUT(N__29904),
            .PACKAGEPIN(uart_drone_data_rdy_debug));
    defparam uart_drone_data_rdy_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_drone_data_rdy_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_drone_data_rdy_debug_obuf_preio (
            .PADOEN(N__29906),
            .PADOUT(N__29905),
            .PADIN(N__29904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_commands_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_commands_input_debug_obuf_iopad (
            .OE(N__29897),
            .DIN(N__29896),
            .DOUT(N__29895),
            .PACKAGEPIN(uart_commands_input_debug));
    defparam uart_commands_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_commands_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_commands_input_debug_obuf_preio (
            .PADOEN(N__29897),
            .PADOUT(N__29896),
            .PADIN(N__29895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam drone_frame_decoder_data_rdy_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD drone_frame_decoder_data_rdy_debug_obuf_iopad (
            .OE(N__29888),
            .DIN(N__29887),
            .DOUT(N__29886),
            .PACKAGEPIN(drone_frame_decoder_data_rdy_debug));
    defparam drone_frame_decoder_data_rdy_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam drone_frame_decoder_data_rdy_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO drone_frame_decoder_data_rdy_debug_obuf_preio (
            .PADOEN(N__29888),
            .PADOUT(N__29887),
            .PADIN(N__29886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13846),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_drone_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_drone_input_debug_obuf_iopad (
            .OE(N__29879),
            .DIN(N__29878),
            .DOUT(N__29877),
            .PACKAGEPIN(uart_drone_input_debug));
    defparam uart_drone_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_drone_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_drone_input_debug_obuf_preio (
            .PADOEN(N__29879),
            .PADOUT(N__29878),
            .PADIN(N__29877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21749),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__7203 (
            .O(N__29860),
            .I(N__29857));
    LocalMux I__7202 (
            .O(N__29857),
            .I(N__29853));
    InMux I__7201 (
            .O(N__29856),
            .I(N__29850));
    Span4Mux_h I__7200 (
            .O(N__29853),
            .I(N__29840));
    LocalMux I__7199 (
            .O(N__29850),
            .I(N__29840));
    InMux I__7198 (
            .O(N__29849),
            .I(N__29835));
    InMux I__7197 (
            .O(N__29848),
            .I(N__29832));
    InMux I__7196 (
            .O(N__29847),
            .I(N__29828));
    InMux I__7195 (
            .O(N__29846),
            .I(N__29823));
    InMux I__7194 (
            .O(N__29845),
            .I(N__29820));
    Span4Mux_v I__7193 (
            .O(N__29840),
            .I(N__29817));
    InMux I__7192 (
            .O(N__29839),
            .I(N__29814));
    InMux I__7191 (
            .O(N__29838),
            .I(N__29811));
    LocalMux I__7190 (
            .O(N__29835),
            .I(N__29808));
    LocalMux I__7189 (
            .O(N__29832),
            .I(N__29805));
    InMux I__7188 (
            .O(N__29831),
            .I(N__29802));
    LocalMux I__7187 (
            .O(N__29828),
            .I(N__29799));
    InMux I__7186 (
            .O(N__29827),
            .I(N__29796));
    CascadeMux I__7185 (
            .O(N__29826),
            .I(N__29793));
    LocalMux I__7184 (
            .O(N__29823),
            .I(N__29790));
    LocalMux I__7183 (
            .O(N__29820),
            .I(N__29787));
    Sp12to4 I__7182 (
            .O(N__29817),
            .I(N__29782));
    LocalMux I__7181 (
            .O(N__29814),
            .I(N__29782));
    LocalMux I__7180 (
            .O(N__29811),
            .I(N__29779));
    Span4Mux_v I__7179 (
            .O(N__29808),
            .I(N__29774));
    Span4Mux_h I__7178 (
            .O(N__29805),
            .I(N__29774));
    LocalMux I__7177 (
            .O(N__29802),
            .I(N__29771));
    Span4Mux_h I__7176 (
            .O(N__29799),
            .I(N__29766));
    LocalMux I__7175 (
            .O(N__29796),
            .I(N__29766));
    InMux I__7174 (
            .O(N__29793),
            .I(N__29763));
    Span4Mux_h I__7173 (
            .O(N__29790),
            .I(N__29760));
    Span4Mux_h I__7172 (
            .O(N__29787),
            .I(N__29757));
    Span12Mux_h I__7171 (
            .O(N__29782),
            .I(N__29754));
    Span4Mux_v I__7170 (
            .O(N__29779),
            .I(N__29745));
    Span4Mux_h I__7169 (
            .O(N__29774),
            .I(N__29745));
    Span4Mux_v I__7168 (
            .O(N__29771),
            .I(N__29745));
    Span4Mux_v I__7167 (
            .O(N__29766),
            .I(N__29745));
    LocalMux I__7166 (
            .O(N__29763),
            .I(uart_pc_data_0));
    Odrv4 I__7165 (
            .O(N__29760),
            .I(uart_pc_data_0));
    Odrv4 I__7164 (
            .O(N__29757),
            .I(uart_pc_data_0));
    Odrv12 I__7163 (
            .O(N__29754),
            .I(uart_pc_data_0));
    Odrv4 I__7162 (
            .O(N__29745),
            .I(uart_pc_data_0));
    InMux I__7161 (
            .O(N__29734),
            .I(N__29731));
    LocalMux I__7160 (
            .O(N__29731),
            .I(N__29726));
    InMux I__7159 (
            .O(N__29730),
            .I(N__29723));
    CascadeMux I__7158 (
            .O(N__29729),
            .I(N__29719));
    Span4Mux_h I__7157 (
            .O(N__29726),
            .I(N__29716));
    LocalMux I__7156 (
            .O(N__29723),
            .I(N__29713));
    InMux I__7155 (
            .O(N__29722),
            .I(N__29710));
    InMux I__7154 (
            .O(N__29719),
            .I(N__29707));
    Odrv4 I__7153 (
            .O(N__29716),
            .I(frame_decoder_OFF3data_0));
    Odrv12 I__7152 (
            .O(N__29713),
            .I(frame_decoder_OFF3data_0));
    LocalMux I__7151 (
            .O(N__29710),
            .I(frame_decoder_OFF3data_0));
    LocalMux I__7150 (
            .O(N__29707),
            .I(frame_decoder_OFF3data_0));
    InMux I__7149 (
            .O(N__29698),
            .I(N__29695));
    LocalMux I__7148 (
            .O(N__29695),
            .I(N__29692));
    Span4Mux_h I__7147 (
            .O(N__29692),
            .I(N__29689));
    Odrv4 I__7146 (
            .O(N__29689),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    CascadeMux I__7145 (
            .O(N__29686),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ));
    CEMux I__7144 (
            .O(N__29683),
            .I(N__29679));
    CEMux I__7143 (
            .O(N__29682),
            .I(N__29676));
    LocalMux I__7142 (
            .O(N__29679),
            .I(N__29673));
    LocalMux I__7141 (
            .O(N__29676),
            .I(N__29670));
    Span4Mux_v I__7140 (
            .O(N__29673),
            .I(N__29667));
    Span4Mux_v I__7139 (
            .O(N__29670),
            .I(N__29664));
    Odrv4 I__7138 (
            .O(N__29667),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    Odrv4 I__7137 (
            .O(N__29664),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__7136 (
            .O(N__29659),
            .I(N__29653));
    InMux I__7135 (
            .O(N__29658),
            .I(N__29650));
    InMux I__7134 (
            .O(N__29657),
            .I(N__29644));
    InMux I__7133 (
            .O(N__29656),
            .I(N__29641));
    LocalMux I__7132 (
            .O(N__29653),
            .I(N__29637));
    LocalMux I__7131 (
            .O(N__29650),
            .I(N__29634));
    InMux I__7130 (
            .O(N__29649),
            .I(N__29631));
    InMux I__7129 (
            .O(N__29648),
            .I(N__29628));
    InMux I__7128 (
            .O(N__29647),
            .I(N__29625));
    LocalMux I__7127 (
            .O(N__29644),
            .I(N__29622));
    LocalMux I__7126 (
            .O(N__29641),
            .I(N__29619));
    InMux I__7125 (
            .O(N__29640),
            .I(N__29615));
    Span4Mux_v I__7124 (
            .O(N__29637),
            .I(N__29610));
    Span4Mux_h I__7123 (
            .O(N__29634),
            .I(N__29601));
    LocalMux I__7122 (
            .O(N__29631),
            .I(N__29601));
    LocalMux I__7121 (
            .O(N__29628),
            .I(N__29601));
    LocalMux I__7120 (
            .O(N__29625),
            .I(N__29601));
    Span4Mux_v I__7119 (
            .O(N__29622),
            .I(N__29595));
    Span4Mux_h I__7118 (
            .O(N__29619),
            .I(N__29595));
    InMux I__7117 (
            .O(N__29618),
            .I(N__29592));
    LocalMux I__7116 (
            .O(N__29615),
            .I(N__29584));
    InMux I__7115 (
            .O(N__29614),
            .I(N__29579));
    InMux I__7114 (
            .O(N__29613),
            .I(N__29579));
    Span4Mux_h I__7113 (
            .O(N__29610),
            .I(N__29574));
    Span4Mux_v I__7112 (
            .O(N__29601),
            .I(N__29574));
    InMux I__7111 (
            .O(N__29600),
            .I(N__29571));
    Span4Mux_h I__7110 (
            .O(N__29595),
            .I(N__29568));
    LocalMux I__7109 (
            .O(N__29592),
            .I(N__29565));
    InMux I__7108 (
            .O(N__29591),
            .I(N__29558));
    InMux I__7107 (
            .O(N__29590),
            .I(N__29558));
    InMux I__7106 (
            .O(N__29589),
            .I(N__29558));
    InMux I__7105 (
            .O(N__29588),
            .I(N__29553));
    InMux I__7104 (
            .O(N__29587),
            .I(N__29553));
    Span4Mux_v I__7103 (
            .O(N__29584),
            .I(N__29548));
    LocalMux I__7102 (
            .O(N__29579),
            .I(N__29548));
    Span4Mux_h I__7101 (
            .O(N__29574),
            .I(N__29545));
    LocalMux I__7100 (
            .O(N__29571),
            .I(uart_pc_data_rdy));
    Odrv4 I__7099 (
            .O(N__29568),
            .I(uart_pc_data_rdy));
    Odrv4 I__7098 (
            .O(N__29565),
            .I(uart_pc_data_rdy));
    LocalMux I__7097 (
            .O(N__29558),
            .I(uart_pc_data_rdy));
    LocalMux I__7096 (
            .O(N__29553),
            .I(uart_pc_data_rdy));
    Odrv4 I__7095 (
            .O(N__29548),
            .I(uart_pc_data_rdy));
    Odrv4 I__7094 (
            .O(N__29545),
            .I(uart_pc_data_rdy));
    CascadeMux I__7093 (
            .O(N__29530),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ));
    CEMux I__7092 (
            .O(N__29527),
            .I(N__29524));
    LocalMux I__7091 (
            .O(N__29524),
            .I(N__29520));
    CEMux I__7090 (
            .O(N__29523),
            .I(N__29517));
    Span4Mux_h I__7089 (
            .O(N__29520),
            .I(N__29514));
    LocalMux I__7088 (
            .O(N__29517),
            .I(N__29511));
    Odrv4 I__7087 (
            .O(N__29514),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    Odrv12 I__7086 (
            .O(N__29511),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    InMux I__7085 (
            .O(N__29506),
            .I(N__29502));
    InMux I__7084 (
            .O(N__29505),
            .I(N__29499));
    LocalMux I__7083 (
            .O(N__29502),
            .I(N__29496));
    LocalMux I__7082 (
            .O(N__29499),
            .I(N__29493));
    Span4Mux_h I__7081 (
            .O(N__29496),
            .I(N__29490));
    Span4Mux_v I__7080 (
            .O(N__29493),
            .I(N__29487));
    Odrv4 I__7079 (
            .O(N__29490),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa ));
    Odrv4 I__7078 (
            .O(N__29487),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa ));
    InMux I__7077 (
            .O(N__29482),
            .I(N__29478));
    InMux I__7076 (
            .O(N__29481),
            .I(N__29475));
    LocalMux I__7075 (
            .O(N__29478),
            .I(\Commands_frame_decoder.state_1Z0Z_8 ));
    LocalMux I__7074 (
            .O(N__29475),
            .I(\Commands_frame_decoder.state_1Z0Z_8 ));
    InMux I__7073 (
            .O(N__29470),
            .I(N__29464));
    InMux I__7072 (
            .O(N__29469),
            .I(N__29464));
    LocalMux I__7071 (
            .O(N__29464),
            .I(N__29452));
    InMux I__7070 (
            .O(N__29463),
            .I(N__29449));
    InMux I__7069 (
            .O(N__29462),
            .I(N__29442));
    InMux I__7068 (
            .O(N__29461),
            .I(N__29442));
    InMux I__7067 (
            .O(N__29460),
            .I(N__29442));
    InMux I__7066 (
            .O(N__29459),
            .I(N__29437));
    InMux I__7065 (
            .O(N__29458),
            .I(N__29437));
    InMux I__7064 (
            .O(N__29457),
            .I(N__29430));
    InMux I__7063 (
            .O(N__29456),
            .I(N__29430));
    InMux I__7062 (
            .O(N__29455),
            .I(N__29430));
    Span12Mux_h I__7061 (
            .O(N__29452),
            .I(N__29423));
    LocalMux I__7060 (
            .O(N__29449),
            .I(N__29423));
    LocalMux I__7059 (
            .O(N__29442),
            .I(N__29423));
    LocalMux I__7058 (
            .O(N__29437),
            .I(N__29420));
    LocalMux I__7057 (
            .O(N__29430),
            .I(N__29417));
    Odrv12 I__7056 (
            .O(N__29423),
            .I(\Commands_frame_decoder.N_316 ));
    Odrv4 I__7055 (
            .O(N__29420),
            .I(\Commands_frame_decoder.N_316 ));
    Odrv4 I__7054 (
            .O(N__29417),
            .I(\Commands_frame_decoder.N_316 ));
    InMux I__7053 (
            .O(N__29410),
            .I(N__29407));
    LocalMux I__7052 (
            .O(N__29407),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa ));
    InMux I__7051 (
            .O(N__29404),
            .I(N__29400));
    InMux I__7050 (
            .O(N__29403),
            .I(N__29397));
    LocalMux I__7049 (
            .O(N__29400),
            .I(\Commands_frame_decoder.state_1Z0Z_9 ));
    LocalMux I__7048 (
            .O(N__29397),
            .I(\Commands_frame_decoder.state_1Z0Z_9 ));
    ClkMux I__7047 (
            .O(N__29392),
            .I(N__28987));
    ClkMux I__7046 (
            .O(N__29391),
            .I(N__28987));
    ClkMux I__7045 (
            .O(N__29390),
            .I(N__28987));
    ClkMux I__7044 (
            .O(N__29389),
            .I(N__28987));
    ClkMux I__7043 (
            .O(N__29388),
            .I(N__28987));
    ClkMux I__7042 (
            .O(N__29387),
            .I(N__28987));
    ClkMux I__7041 (
            .O(N__29386),
            .I(N__28987));
    ClkMux I__7040 (
            .O(N__29385),
            .I(N__28987));
    ClkMux I__7039 (
            .O(N__29384),
            .I(N__28987));
    ClkMux I__7038 (
            .O(N__29383),
            .I(N__28987));
    ClkMux I__7037 (
            .O(N__29382),
            .I(N__28987));
    ClkMux I__7036 (
            .O(N__29381),
            .I(N__28987));
    ClkMux I__7035 (
            .O(N__29380),
            .I(N__28987));
    ClkMux I__7034 (
            .O(N__29379),
            .I(N__28987));
    ClkMux I__7033 (
            .O(N__29378),
            .I(N__28987));
    ClkMux I__7032 (
            .O(N__29377),
            .I(N__28987));
    ClkMux I__7031 (
            .O(N__29376),
            .I(N__28987));
    ClkMux I__7030 (
            .O(N__29375),
            .I(N__28987));
    ClkMux I__7029 (
            .O(N__29374),
            .I(N__28987));
    ClkMux I__7028 (
            .O(N__29373),
            .I(N__28987));
    ClkMux I__7027 (
            .O(N__29372),
            .I(N__28987));
    ClkMux I__7026 (
            .O(N__29371),
            .I(N__28987));
    ClkMux I__7025 (
            .O(N__29370),
            .I(N__28987));
    ClkMux I__7024 (
            .O(N__29369),
            .I(N__28987));
    ClkMux I__7023 (
            .O(N__29368),
            .I(N__28987));
    ClkMux I__7022 (
            .O(N__29367),
            .I(N__28987));
    ClkMux I__7021 (
            .O(N__29366),
            .I(N__28987));
    ClkMux I__7020 (
            .O(N__29365),
            .I(N__28987));
    ClkMux I__7019 (
            .O(N__29364),
            .I(N__28987));
    ClkMux I__7018 (
            .O(N__29363),
            .I(N__28987));
    ClkMux I__7017 (
            .O(N__29362),
            .I(N__28987));
    ClkMux I__7016 (
            .O(N__29361),
            .I(N__28987));
    ClkMux I__7015 (
            .O(N__29360),
            .I(N__28987));
    ClkMux I__7014 (
            .O(N__29359),
            .I(N__28987));
    ClkMux I__7013 (
            .O(N__29358),
            .I(N__28987));
    ClkMux I__7012 (
            .O(N__29357),
            .I(N__28987));
    ClkMux I__7011 (
            .O(N__29356),
            .I(N__28987));
    ClkMux I__7010 (
            .O(N__29355),
            .I(N__28987));
    ClkMux I__7009 (
            .O(N__29354),
            .I(N__28987));
    ClkMux I__7008 (
            .O(N__29353),
            .I(N__28987));
    ClkMux I__7007 (
            .O(N__29352),
            .I(N__28987));
    ClkMux I__7006 (
            .O(N__29351),
            .I(N__28987));
    ClkMux I__7005 (
            .O(N__29350),
            .I(N__28987));
    ClkMux I__7004 (
            .O(N__29349),
            .I(N__28987));
    ClkMux I__7003 (
            .O(N__29348),
            .I(N__28987));
    ClkMux I__7002 (
            .O(N__29347),
            .I(N__28987));
    ClkMux I__7001 (
            .O(N__29346),
            .I(N__28987));
    ClkMux I__7000 (
            .O(N__29345),
            .I(N__28987));
    ClkMux I__6999 (
            .O(N__29344),
            .I(N__28987));
    ClkMux I__6998 (
            .O(N__29343),
            .I(N__28987));
    ClkMux I__6997 (
            .O(N__29342),
            .I(N__28987));
    ClkMux I__6996 (
            .O(N__29341),
            .I(N__28987));
    ClkMux I__6995 (
            .O(N__29340),
            .I(N__28987));
    ClkMux I__6994 (
            .O(N__29339),
            .I(N__28987));
    ClkMux I__6993 (
            .O(N__29338),
            .I(N__28987));
    ClkMux I__6992 (
            .O(N__29337),
            .I(N__28987));
    ClkMux I__6991 (
            .O(N__29336),
            .I(N__28987));
    ClkMux I__6990 (
            .O(N__29335),
            .I(N__28987));
    ClkMux I__6989 (
            .O(N__29334),
            .I(N__28987));
    ClkMux I__6988 (
            .O(N__29333),
            .I(N__28987));
    ClkMux I__6987 (
            .O(N__29332),
            .I(N__28987));
    ClkMux I__6986 (
            .O(N__29331),
            .I(N__28987));
    ClkMux I__6985 (
            .O(N__29330),
            .I(N__28987));
    ClkMux I__6984 (
            .O(N__29329),
            .I(N__28987));
    ClkMux I__6983 (
            .O(N__29328),
            .I(N__28987));
    ClkMux I__6982 (
            .O(N__29327),
            .I(N__28987));
    ClkMux I__6981 (
            .O(N__29326),
            .I(N__28987));
    ClkMux I__6980 (
            .O(N__29325),
            .I(N__28987));
    ClkMux I__6979 (
            .O(N__29324),
            .I(N__28987));
    ClkMux I__6978 (
            .O(N__29323),
            .I(N__28987));
    ClkMux I__6977 (
            .O(N__29322),
            .I(N__28987));
    ClkMux I__6976 (
            .O(N__29321),
            .I(N__28987));
    ClkMux I__6975 (
            .O(N__29320),
            .I(N__28987));
    ClkMux I__6974 (
            .O(N__29319),
            .I(N__28987));
    ClkMux I__6973 (
            .O(N__29318),
            .I(N__28987));
    ClkMux I__6972 (
            .O(N__29317),
            .I(N__28987));
    ClkMux I__6971 (
            .O(N__29316),
            .I(N__28987));
    ClkMux I__6970 (
            .O(N__29315),
            .I(N__28987));
    ClkMux I__6969 (
            .O(N__29314),
            .I(N__28987));
    ClkMux I__6968 (
            .O(N__29313),
            .I(N__28987));
    ClkMux I__6967 (
            .O(N__29312),
            .I(N__28987));
    ClkMux I__6966 (
            .O(N__29311),
            .I(N__28987));
    ClkMux I__6965 (
            .O(N__29310),
            .I(N__28987));
    ClkMux I__6964 (
            .O(N__29309),
            .I(N__28987));
    ClkMux I__6963 (
            .O(N__29308),
            .I(N__28987));
    ClkMux I__6962 (
            .O(N__29307),
            .I(N__28987));
    ClkMux I__6961 (
            .O(N__29306),
            .I(N__28987));
    ClkMux I__6960 (
            .O(N__29305),
            .I(N__28987));
    ClkMux I__6959 (
            .O(N__29304),
            .I(N__28987));
    ClkMux I__6958 (
            .O(N__29303),
            .I(N__28987));
    ClkMux I__6957 (
            .O(N__29302),
            .I(N__28987));
    ClkMux I__6956 (
            .O(N__29301),
            .I(N__28987));
    ClkMux I__6955 (
            .O(N__29300),
            .I(N__28987));
    ClkMux I__6954 (
            .O(N__29299),
            .I(N__28987));
    ClkMux I__6953 (
            .O(N__29298),
            .I(N__28987));
    ClkMux I__6952 (
            .O(N__29297),
            .I(N__28987));
    ClkMux I__6951 (
            .O(N__29296),
            .I(N__28987));
    ClkMux I__6950 (
            .O(N__29295),
            .I(N__28987));
    ClkMux I__6949 (
            .O(N__29294),
            .I(N__28987));
    ClkMux I__6948 (
            .O(N__29293),
            .I(N__28987));
    ClkMux I__6947 (
            .O(N__29292),
            .I(N__28987));
    ClkMux I__6946 (
            .O(N__29291),
            .I(N__28987));
    ClkMux I__6945 (
            .O(N__29290),
            .I(N__28987));
    ClkMux I__6944 (
            .O(N__29289),
            .I(N__28987));
    ClkMux I__6943 (
            .O(N__29288),
            .I(N__28987));
    ClkMux I__6942 (
            .O(N__29287),
            .I(N__28987));
    ClkMux I__6941 (
            .O(N__29286),
            .I(N__28987));
    ClkMux I__6940 (
            .O(N__29285),
            .I(N__28987));
    ClkMux I__6939 (
            .O(N__29284),
            .I(N__28987));
    ClkMux I__6938 (
            .O(N__29283),
            .I(N__28987));
    ClkMux I__6937 (
            .O(N__29282),
            .I(N__28987));
    ClkMux I__6936 (
            .O(N__29281),
            .I(N__28987));
    ClkMux I__6935 (
            .O(N__29280),
            .I(N__28987));
    ClkMux I__6934 (
            .O(N__29279),
            .I(N__28987));
    ClkMux I__6933 (
            .O(N__29278),
            .I(N__28987));
    ClkMux I__6932 (
            .O(N__29277),
            .I(N__28987));
    ClkMux I__6931 (
            .O(N__29276),
            .I(N__28987));
    ClkMux I__6930 (
            .O(N__29275),
            .I(N__28987));
    ClkMux I__6929 (
            .O(N__29274),
            .I(N__28987));
    ClkMux I__6928 (
            .O(N__29273),
            .I(N__28987));
    ClkMux I__6927 (
            .O(N__29272),
            .I(N__28987));
    ClkMux I__6926 (
            .O(N__29271),
            .I(N__28987));
    ClkMux I__6925 (
            .O(N__29270),
            .I(N__28987));
    ClkMux I__6924 (
            .O(N__29269),
            .I(N__28987));
    ClkMux I__6923 (
            .O(N__29268),
            .I(N__28987));
    ClkMux I__6922 (
            .O(N__29267),
            .I(N__28987));
    ClkMux I__6921 (
            .O(N__29266),
            .I(N__28987));
    ClkMux I__6920 (
            .O(N__29265),
            .I(N__28987));
    ClkMux I__6919 (
            .O(N__29264),
            .I(N__28987));
    ClkMux I__6918 (
            .O(N__29263),
            .I(N__28987));
    ClkMux I__6917 (
            .O(N__29262),
            .I(N__28987));
    ClkMux I__6916 (
            .O(N__29261),
            .I(N__28987));
    ClkMux I__6915 (
            .O(N__29260),
            .I(N__28987));
    ClkMux I__6914 (
            .O(N__29259),
            .I(N__28987));
    ClkMux I__6913 (
            .O(N__29258),
            .I(N__28987));
    GlobalMux I__6912 (
            .O(N__28987),
            .I(N__28984));
    gio2CtrlBuf I__6911 (
            .O(N__28984),
            .I(clk_system_c_g));
    CascadeMux I__6910 (
            .O(N__28981),
            .I(N__28973));
    CascadeMux I__6909 (
            .O(N__28980),
            .I(N__28969));
    CascadeMux I__6908 (
            .O(N__28979),
            .I(N__28965));
    InMux I__6907 (
            .O(N__28978),
            .I(N__28921));
    InMux I__6906 (
            .O(N__28977),
            .I(N__28916));
    InMux I__6905 (
            .O(N__28976),
            .I(N__28916));
    InMux I__6904 (
            .O(N__28973),
            .I(N__28913));
    InMux I__6903 (
            .O(N__28972),
            .I(N__28908));
    InMux I__6902 (
            .O(N__28969),
            .I(N__28908));
    InMux I__6901 (
            .O(N__28968),
            .I(N__28905));
    InMux I__6900 (
            .O(N__28965),
            .I(N__28900));
    InMux I__6899 (
            .O(N__28964),
            .I(N__28900));
    InMux I__6898 (
            .O(N__28963),
            .I(N__28897));
    InMux I__6897 (
            .O(N__28962),
            .I(N__28892));
    InMux I__6896 (
            .O(N__28961),
            .I(N__28892));
    InMux I__6895 (
            .O(N__28960),
            .I(N__28889));
    InMux I__6894 (
            .O(N__28959),
            .I(N__28878));
    InMux I__6893 (
            .O(N__28958),
            .I(N__28878));
    InMux I__6892 (
            .O(N__28957),
            .I(N__28878));
    InMux I__6891 (
            .O(N__28956),
            .I(N__28878));
    InMux I__6890 (
            .O(N__28955),
            .I(N__28878));
    InMux I__6889 (
            .O(N__28954),
            .I(N__28867));
    InMux I__6888 (
            .O(N__28953),
            .I(N__28867));
    InMux I__6887 (
            .O(N__28952),
            .I(N__28867));
    InMux I__6886 (
            .O(N__28951),
            .I(N__28867));
    InMux I__6885 (
            .O(N__28950),
            .I(N__28867));
    InMux I__6884 (
            .O(N__28949),
            .I(N__28862));
    InMux I__6883 (
            .O(N__28948),
            .I(N__28862));
    InMux I__6882 (
            .O(N__28947),
            .I(N__28855));
    InMux I__6881 (
            .O(N__28946),
            .I(N__28855));
    InMux I__6880 (
            .O(N__28945),
            .I(N__28855));
    InMux I__6879 (
            .O(N__28944),
            .I(N__28844));
    InMux I__6878 (
            .O(N__28943),
            .I(N__28844));
    InMux I__6877 (
            .O(N__28942),
            .I(N__28844));
    InMux I__6876 (
            .O(N__28941),
            .I(N__28844));
    InMux I__6875 (
            .O(N__28940),
            .I(N__28844));
    InMux I__6874 (
            .O(N__28939),
            .I(N__28841));
    InMux I__6873 (
            .O(N__28938),
            .I(N__28838));
    InMux I__6872 (
            .O(N__28937),
            .I(N__28835));
    InMux I__6871 (
            .O(N__28936),
            .I(N__28830));
    InMux I__6870 (
            .O(N__28935),
            .I(N__28830));
    InMux I__6869 (
            .O(N__28934),
            .I(N__28827));
    InMux I__6868 (
            .O(N__28933),
            .I(N__28824));
    InMux I__6867 (
            .O(N__28932),
            .I(N__28821));
    InMux I__6866 (
            .O(N__28931),
            .I(N__28818));
    InMux I__6865 (
            .O(N__28930),
            .I(N__28815));
    InMux I__6864 (
            .O(N__28929),
            .I(N__28812));
    InMux I__6863 (
            .O(N__28928),
            .I(N__28809));
    InMux I__6862 (
            .O(N__28927),
            .I(N__28806));
    InMux I__6861 (
            .O(N__28926),
            .I(N__28803));
    InMux I__6860 (
            .O(N__28925),
            .I(N__28800));
    InMux I__6859 (
            .O(N__28924),
            .I(N__28797));
    LocalMux I__6858 (
            .O(N__28921),
            .I(N__28708));
    LocalMux I__6857 (
            .O(N__28916),
            .I(N__28705));
    LocalMux I__6856 (
            .O(N__28913),
            .I(N__28702));
    LocalMux I__6855 (
            .O(N__28908),
            .I(N__28699));
    LocalMux I__6854 (
            .O(N__28905),
            .I(N__28696));
    LocalMux I__6853 (
            .O(N__28900),
            .I(N__28693));
    LocalMux I__6852 (
            .O(N__28897),
            .I(N__28690));
    LocalMux I__6851 (
            .O(N__28892),
            .I(N__28687));
    LocalMux I__6850 (
            .O(N__28889),
            .I(N__28684));
    LocalMux I__6849 (
            .O(N__28878),
            .I(N__28681));
    LocalMux I__6848 (
            .O(N__28867),
            .I(N__28678));
    LocalMux I__6847 (
            .O(N__28862),
            .I(N__28675));
    LocalMux I__6846 (
            .O(N__28855),
            .I(N__28672));
    LocalMux I__6845 (
            .O(N__28844),
            .I(N__28669));
    LocalMux I__6844 (
            .O(N__28841),
            .I(N__28666));
    LocalMux I__6843 (
            .O(N__28838),
            .I(N__28663));
    LocalMux I__6842 (
            .O(N__28835),
            .I(N__28660));
    LocalMux I__6841 (
            .O(N__28830),
            .I(N__28657));
    LocalMux I__6840 (
            .O(N__28827),
            .I(N__28654));
    LocalMux I__6839 (
            .O(N__28824),
            .I(N__28651));
    LocalMux I__6838 (
            .O(N__28821),
            .I(N__28648));
    LocalMux I__6837 (
            .O(N__28818),
            .I(N__28645));
    LocalMux I__6836 (
            .O(N__28815),
            .I(N__28642));
    LocalMux I__6835 (
            .O(N__28812),
            .I(N__28639));
    LocalMux I__6834 (
            .O(N__28809),
            .I(N__28636));
    LocalMux I__6833 (
            .O(N__28806),
            .I(N__28633));
    LocalMux I__6832 (
            .O(N__28803),
            .I(N__28630));
    LocalMux I__6831 (
            .O(N__28800),
            .I(N__28627));
    LocalMux I__6830 (
            .O(N__28797),
            .I(N__28624));
    SRMux I__6829 (
            .O(N__28796),
            .I(N__28393));
    SRMux I__6828 (
            .O(N__28795),
            .I(N__28393));
    SRMux I__6827 (
            .O(N__28794),
            .I(N__28393));
    SRMux I__6826 (
            .O(N__28793),
            .I(N__28393));
    SRMux I__6825 (
            .O(N__28792),
            .I(N__28393));
    SRMux I__6824 (
            .O(N__28791),
            .I(N__28393));
    SRMux I__6823 (
            .O(N__28790),
            .I(N__28393));
    SRMux I__6822 (
            .O(N__28789),
            .I(N__28393));
    SRMux I__6821 (
            .O(N__28788),
            .I(N__28393));
    SRMux I__6820 (
            .O(N__28787),
            .I(N__28393));
    SRMux I__6819 (
            .O(N__28786),
            .I(N__28393));
    SRMux I__6818 (
            .O(N__28785),
            .I(N__28393));
    SRMux I__6817 (
            .O(N__28784),
            .I(N__28393));
    SRMux I__6816 (
            .O(N__28783),
            .I(N__28393));
    SRMux I__6815 (
            .O(N__28782),
            .I(N__28393));
    SRMux I__6814 (
            .O(N__28781),
            .I(N__28393));
    SRMux I__6813 (
            .O(N__28780),
            .I(N__28393));
    SRMux I__6812 (
            .O(N__28779),
            .I(N__28393));
    SRMux I__6811 (
            .O(N__28778),
            .I(N__28393));
    SRMux I__6810 (
            .O(N__28777),
            .I(N__28393));
    SRMux I__6809 (
            .O(N__28776),
            .I(N__28393));
    SRMux I__6808 (
            .O(N__28775),
            .I(N__28393));
    SRMux I__6807 (
            .O(N__28774),
            .I(N__28393));
    SRMux I__6806 (
            .O(N__28773),
            .I(N__28393));
    SRMux I__6805 (
            .O(N__28772),
            .I(N__28393));
    SRMux I__6804 (
            .O(N__28771),
            .I(N__28393));
    SRMux I__6803 (
            .O(N__28770),
            .I(N__28393));
    SRMux I__6802 (
            .O(N__28769),
            .I(N__28393));
    SRMux I__6801 (
            .O(N__28768),
            .I(N__28393));
    SRMux I__6800 (
            .O(N__28767),
            .I(N__28393));
    SRMux I__6799 (
            .O(N__28766),
            .I(N__28393));
    SRMux I__6798 (
            .O(N__28765),
            .I(N__28393));
    SRMux I__6797 (
            .O(N__28764),
            .I(N__28393));
    SRMux I__6796 (
            .O(N__28763),
            .I(N__28393));
    SRMux I__6795 (
            .O(N__28762),
            .I(N__28393));
    SRMux I__6794 (
            .O(N__28761),
            .I(N__28393));
    SRMux I__6793 (
            .O(N__28760),
            .I(N__28393));
    SRMux I__6792 (
            .O(N__28759),
            .I(N__28393));
    SRMux I__6791 (
            .O(N__28758),
            .I(N__28393));
    SRMux I__6790 (
            .O(N__28757),
            .I(N__28393));
    SRMux I__6789 (
            .O(N__28756),
            .I(N__28393));
    SRMux I__6788 (
            .O(N__28755),
            .I(N__28393));
    SRMux I__6787 (
            .O(N__28754),
            .I(N__28393));
    SRMux I__6786 (
            .O(N__28753),
            .I(N__28393));
    SRMux I__6785 (
            .O(N__28752),
            .I(N__28393));
    SRMux I__6784 (
            .O(N__28751),
            .I(N__28393));
    SRMux I__6783 (
            .O(N__28750),
            .I(N__28393));
    SRMux I__6782 (
            .O(N__28749),
            .I(N__28393));
    SRMux I__6781 (
            .O(N__28748),
            .I(N__28393));
    SRMux I__6780 (
            .O(N__28747),
            .I(N__28393));
    SRMux I__6779 (
            .O(N__28746),
            .I(N__28393));
    SRMux I__6778 (
            .O(N__28745),
            .I(N__28393));
    SRMux I__6777 (
            .O(N__28744),
            .I(N__28393));
    SRMux I__6776 (
            .O(N__28743),
            .I(N__28393));
    SRMux I__6775 (
            .O(N__28742),
            .I(N__28393));
    SRMux I__6774 (
            .O(N__28741),
            .I(N__28393));
    SRMux I__6773 (
            .O(N__28740),
            .I(N__28393));
    SRMux I__6772 (
            .O(N__28739),
            .I(N__28393));
    SRMux I__6771 (
            .O(N__28738),
            .I(N__28393));
    SRMux I__6770 (
            .O(N__28737),
            .I(N__28393));
    SRMux I__6769 (
            .O(N__28736),
            .I(N__28393));
    SRMux I__6768 (
            .O(N__28735),
            .I(N__28393));
    SRMux I__6767 (
            .O(N__28734),
            .I(N__28393));
    SRMux I__6766 (
            .O(N__28733),
            .I(N__28393));
    SRMux I__6765 (
            .O(N__28732),
            .I(N__28393));
    SRMux I__6764 (
            .O(N__28731),
            .I(N__28393));
    SRMux I__6763 (
            .O(N__28730),
            .I(N__28393));
    SRMux I__6762 (
            .O(N__28729),
            .I(N__28393));
    SRMux I__6761 (
            .O(N__28728),
            .I(N__28393));
    SRMux I__6760 (
            .O(N__28727),
            .I(N__28393));
    SRMux I__6759 (
            .O(N__28726),
            .I(N__28393));
    SRMux I__6758 (
            .O(N__28725),
            .I(N__28393));
    SRMux I__6757 (
            .O(N__28724),
            .I(N__28393));
    SRMux I__6756 (
            .O(N__28723),
            .I(N__28393));
    SRMux I__6755 (
            .O(N__28722),
            .I(N__28393));
    SRMux I__6754 (
            .O(N__28721),
            .I(N__28393));
    SRMux I__6753 (
            .O(N__28720),
            .I(N__28393));
    SRMux I__6752 (
            .O(N__28719),
            .I(N__28393));
    SRMux I__6751 (
            .O(N__28718),
            .I(N__28393));
    SRMux I__6750 (
            .O(N__28717),
            .I(N__28393));
    SRMux I__6749 (
            .O(N__28716),
            .I(N__28393));
    SRMux I__6748 (
            .O(N__28715),
            .I(N__28393));
    SRMux I__6747 (
            .O(N__28714),
            .I(N__28393));
    SRMux I__6746 (
            .O(N__28713),
            .I(N__28393));
    SRMux I__6745 (
            .O(N__28712),
            .I(N__28393));
    SRMux I__6744 (
            .O(N__28711),
            .I(N__28393));
    Glb2LocalMux I__6743 (
            .O(N__28708),
            .I(N__28393));
    Glb2LocalMux I__6742 (
            .O(N__28705),
            .I(N__28393));
    Glb2LocalMux I__6741 (
            .O(N__28702),
            .I(N__28393));
    Glb2LocalMux I__6740 (
            .O(N__28699),
            .I(N__28393));
    Glb2LocalMux I__6739 (
            .O(N__28696),
            .I(N__28393));
    Glb2LocalMux I__6738 (
            .O(N__28693),
            .I(N__28393));
    Glb2LocalMux I__6737 (
            .O(N__28690),
            .I(N__28393));
    Glb2LocalMux I__6736 (
            .O(N__28687),
            .I(N__28393));
    Glb2LocalMux I__6735 (
            .O(N__28684),
            .I(N__28393));
    Glb2LocalMux I__6734 (
            .O(N__28681),
            .I(N__28393));
    Glb2LocalMux I__6733 (
            .O(N__28678),
            .I(N__28393));
    Glb2LocalMux I__6732 (
            .O(N__28675),
            .I(N__28393));
    Glb2LocalMux I__6731 (
            .O(N__28672),
            .I(N__28393));
    Glb2LocalMux I__6730 (
            .O(N__28669),
            .I(N__28393));
    Glb2LocalMux I__6729 (
            .O(N__28666),
            .I(N__28393));
    Glb2LocalMux I__6728 (
            .O(N__28663),
            .I(N__28393));
    Glb2LocalMux I__6727 (
            .O(N__28660),
            .I(N__28393));
    Glb2LocalMux I__6726 (
            .O(N__28657),
            .I(N__28393));
    Glb2LocalMux I__6725 (
            .O(N__28654),
            .I(N__28393));
    Glb2LocalMux I__6724 (
            .O(N__28651),
            .I(N__28393));
    Glb2LocalMux I__6723 (
            .O(N__28648),
            .I(N__28393));
    Glb2LocalMux I__6722 (
            .O(N__28645),
            .I(N__28393));
    Glb2LocalMux I__6721 (
            .O(N__28642),
            .I(N__28393));
    Glb2LocalMux I__6720 (
            .O(N__28639),
            .I(N__28393));
    Glb2LocalMux I__6719 (
            .O(N__28636),
            .I(N__28393));
    Glb2LocalMux I__6718 (
            .O(N__28633),
            .I(N__28393));
    Glb2LocalMux I__6717 (
            .O(N__28630),
            .I(N__28393));
    Glb2LocalMux I__6716 (
            .O(N__28627),
            .I(N__28393));
    Glb2LocalMux I__6715 (
            .O(N__28624),
            .I(N__28393));
    GlobalMux I__6714 (
            .O(N__28393),
            .I(N__28390));
    gio2CtrlBuf I__6713 (
            .O(N__28390),
            .I(reset_system_g));
    CascadeMux I__6712 (
            .O(N__28387),
            .I(N__28384));
    InMux I__6711 (
            .O(N__28384),
            .I(N__28381));
    LocalMux I__6710 (
            .O(N__28381),
            .I(N__28378));
    Odrv12 I__6709 (
            .O(N__28378),
            .I(frame_decoder_OFF4data_3));
    CascadeMux I__6708 (
            .O(N__28375),
            .I(N__28372));
    InMux I__6707 (
            .O(N__28372),
            .I(N__28369));
    LocalMux I__6706 (
            .O(N__28369),
            .I(N__28366));
    Odrv4 I__6705 (
            .O(N__28366),
            .I(frame_decoder_OFF4data_6));
    InMux I__6704 (
            .O(N__28363),
            .I(N__28357));
    CascadeMux I__6703 (
            .O(N__28362),
            .I(N__28350));
    InMux I__6702 (
            .O(N__28361),
            .I(N__28347));
    InMux I__6701 (
            .O(N__28360),
            .I(N__28344));
    LocalMux I__6700 (
            .O(N__28357),
            .I(N__28341));
    InMux I__6699 (
            .O(N__28356),
            .I(N__28338));
    InMux I__6698 (
            .O(N__28355),
            .I(N__28335));
    InMux I__6697 (
            .O(N__28354),
            .I(N__28332));
    InMux I__6696 (
            .O(N__28353),
            .I(N__28329));
    InMux I__6695 (
            .O(N__28350),
            .I(N__28326));
    LocalMux I__6694 (
            .O(N__28347),
            .I(N__28323));
    LocalMux I__6693 (
            .O(N__28344),
            .I(N__28316));
    Span4Mux_v I__6692 (
            .O(N__28341),
            .I(N__28316));
    LocalMux I__6691 (
            .O(N__28338),
            .I(N__28316));
    LocalMux I__6690 (
            .O(N__28335),
            .I(N__28313));
    LocalMux I__6689 (
            .O(N__28332),
            .I(N__28302));
    LocalMux I__6688 (
            .O(N__28329),
            .I(N__28302));
    LocalMux I__6687 (
            .O(N__28326),
            .I(N__28299));
    Span4Mux_v I__6686 (
            .O(N__28323),
            .I(N__28294));
    Span4Mux_h I__6685 (
            .O(N__28316),
            .I(N__28294));
    Span4Mux_h I__6684 (
            .O(N__28313),
            .I(N__28291));
    InMux I__6683 (
            .O(N__28312),
            .I(N__28288));
    InMux I__6682 (
            .O(N__28311),
            .I(N__28285));
    InMux I__6681 (
            .O(N__28310),
            .I(N__28282));
    InMux I__6680 (
            .O(N__28309),
            .I(N__28279));
    InMux I__6679 (
            .O(N__28308),
            .I(N__28276));
    InMux I__6678 (
            .O(N__28307),
            .I(N__28273));
    Span12Mux_h I__6677 (
            .O(N__28302),
            .I(N__28270));
    Span4Mux_v I__6676 (
            .O(N__28299),
            .I(N__28267));
    Span4Mux_h I__6675 (
            .O(N__28294),
            .I(N__28260));
    Span4Mux_v I__6674 (
            .O(N__28291),
            .I(N__28260));
    LocalMux I__6673 (
            .O(N__28288),
            .I(N__28260));
    LocalMux I__6672 (
            .O(N__28285),
            .I(N__28251));
    LocalMux I__6671 (
            .O(N__28282),
            .I(N__28251));
    LocalMux I__6670 (
            .O(N__28279),
            .I(N__28251));
    LocalMux I__6669 (
            .O(N__28276),
            .I(N__28251));
    LocalMux I__6668 (
            .O(N__28273),
            .I(uart_pc_data_2));
    Odrv12 I__6667 (
            .O(N__28270),
            .I(uart_pc_data_2));
    Odrv4 I__6666 (
            .O(N__28267),
            .I(uart_pc_data_2));
    Odrv4 I__6665 (
            .O(N__28260),
            .I(uart_pc_data_2));
    Odrv12 I__6664 (
            .O(N__28251),
            .I(uart_pc_data_2));
    CascadeMux I__6663 (
            .O(N__28240),
            .I(N__28237));
    InMux I__6662 (
            .O(N__28237),
            .I(N__28234));
    LocalMux I__6661 (
            .O(N__28234),
            .I(frame_decoder_OFF3data_2));
    InMux I__6660 (
            .O(N__28231),
            .I(N__28225));
    InMux I__6659 (
            .O(N__28230),
            .I(N__28222));
    InMux I__6658 (
            .O(N__28229),
            .I(N__28217));
    InMux I__6657 (
            .O(N__28228),
            .I(N__28214));
    LocalMux I__6656 (
            .O(N__28225),
            .I(N__28210));
    LocalMux I__6655 (
            .O(N__28222),
            .I(N__28207));
    InMux I__6654 (
            .O(N__28221),
            .I(N__28204));
    InMux I__6653 (
            .O(N__28220),
            .I(N__28200));
    LocalMux I__6652 (
            .O(N__28217),
            .I(N__28195));
    LocalMux I__6651 (
            .O(N__28214),
            .I(N__28195));
    InMux I__6650 (
            .O(N__28213),
            .I(N__28191));
    Span4Mux_v I__6649 (
            .O(N__28210),
            .I(N__28188));
    Span4Mux_s3_h I__6648 (
            .O(N__28207),
            .I(N__28185));
    LocalMux I__6647 (
            .O(N__28204),
            .I(N__28182));
    InMux I__6646 (
            .O(N__28203),
            .I(N__28179));
    LocalMux I__6645 (
            .O(N__28200),
            .I(N__28176));
    Span4Mux_v I__6644 (
            .O(N__28195),
            .I(N__28172));
    InMux I__6643 (
            .O(N__28194),
            .I(N__28169));
    LocalMux I__6642 (
            .O(N__28191),
            .I(N__28165));
    Span4Mux_h I__6641 (
            .O(N__28188),
            .I(N__28154));
    Span4Mux_v I__6640 (
            .O(N__28185),
            .I(N__28154));
    Span4Mux_v I__6639 (
            .O(N__28182),
            .I(N__28154));
    LocalMux I__6638 (
            .O(N__28179),
            .I(N__28154));
    Span4Mux_v I__6637 (
            .O(N__28176),
            .I(N__28154));
    CascadeMux I__6636 (
            .O(N__28175),
            .I(N__28151));
    Sp12to4 I__6635 (
            .O(N__28172),
            .I(N__28146));
    LocalMux I__6634 (
            .O(N__28169),
            .I(N__28146));
    InMux I__6633 (
            .O(N__28168),
            .I(N__28143));
    Span12Mux_v I__6632 (
            .O(N__28165),
            .I(N__28138));
    Sp12to4 I__6631 (
            .O(N__28154),
            .I(N__28138));
    InMux I__6630 (
            .O(N__28151),
            .I(N__28135));
    Odrv12 I__6629 (
            .O(N__28146),
            .I(uart_pc_data_6));
    LocalMux I__6628 (
            .O(N__28143),
            .I(uart_pc_data_6));
    Odrv12 I__6627 (
            .O(N__28138),
            .I(uart_pc_data_6));
    LocalMux I__6626 (
            .O(N__28135),
            .I(uart_pc_data_6));
    CascadeMux I__6625 (
            .O(N__28126),
            .I(N__28123));
    InMux I__6624 (
            .O(N__28123),
            .I(N__28120));
    LocalMux I__6623 (
            .O(N__28120),
            .I(frame_decoder_OFF3data_6));
    InMux I__6622 (
            .O(N__28117),
            .I(N__28110));
    InMux I__6621 (
            .O(N__28116),
            .I(N__28107));
    InMux I__6620 (
            .O(N__28115),
            .I(N__28102));
    InMux I__6619 (
            .O(N__28114),
            .I(N__28099));
    InMux I__6618 (
            .O(N__28113),
            .I(N__28095));
    LocalMux I__6617 (
            .O(N__28110),
            .I(N__28092));
    LocalMux I__6616 (
            .O(N__28107),
            .I(N__28089));
    InMux I__6615 (
            .O(N__28106),
            .I(N__28086));
    InMux I__6614 (
            .O(N__28105),
            .I(N__28083));
    LocalMux I__6613 (
            .O(N__28102),
            .I(N__28080));
    LocalMux I__6612 (
            .O(N__28099),
            .I(N__28077));
    InMux I__6611 (
            .O(N__28098),
            .I(N__28073));
    LocalMux I__6610 (
            .O(N__28095),
            .I(N__28070));
    Span4Mux_v I__6609 (
            .O(N__28092),
            .I(N__28065));
    Span4Mux_v I__6608 (
            .O(N__28089),
            .I(N__28065));
    LocalMux I__6607 (
            .O(N__28086),
            .I(N__28060));
    LocalMux I__6606 (
            .O(N__28083),
            .I(N__28053));
    Span4Mux_h I__6605 (
            .O(N__28080),
            .I(N__28053));
    Span4Mux_v I__6604 (
            .O(N__28077),
            .I(N__28053));
    InMux I__6603 (
            .O(N__28076),
            .I(N__28050));
    LocalMux I__6602 (
            .O(N__28073),
            .I(N__28045));
    Span4Mux_v I__6601 (
            .O(N__28070),
            .I(N__28045));
    Span4Mux_h I__6600 (
            .O(N__28065),
            .I(N__28042));
    InMux I__6599 (
            .O(N__28064),
            .I(N__28039));
    InMux I__6598 (
            .O(N__28063),
            .I(N__28036));
    Span12Mux_v I__6597 (
            .O(N__28060),
            .I(N__28033));
    Span4Mux_h I__6596 (
            .O(N__28053),
            .I(N__28028));
    LocalMux I__6595 (
            .O(N__28050),
            .I(N__28028));
    Span4Mux_v I__6594 (
            .O(N__28045),
            .I(N__28021));
    Span4Mux_h I__6593 (
            .O(N__28042),
            .I(N__28021));
    LocalMux I__6592 (
            .O(N__28039),
            .I(N__28021));
    LocalMux I__6591 (
            .O(N__28036),
            .I(uart_pc_data_3));
    Odrv12 I__6590 (
            .O(N__28033),
            .I(uart_pc_data_3));
    Odrv4 I__6589 (
            .O(N__28028),
            .I(uart_pc_data_3));
    Odrv4 I__6588 (
            .O(N__28021),
            .I(uart_pc_data_3));
    CascadeMux I__6587 (
            .O(N__28012),
            .I(N__28009));
    InMux I__6586 (
            .O(N__28009),
            .I(N__28006));
    LocalMux I__6585 (
            .O(N__28006),
            .I(frame_decoder_OFF3data_3));
    InMux I__6584 (
            .O(N__28003),
            .I(N__27997));
    InMux I__6583 (
            .O(N__28002),
            .I(N__27994));
    InMux I__6582 (
            .O(N__28001),
            .I(N__27990));
    InMux I__6581 (
            .O(N__28000),
            .I(N__27986));
    LocalMux I__6580 (
            .O(N__27997),
            .I(N__27981));
    LocalMux I__6579 (
            .O(N__27994),
            .I(N__27981));
    InMux I__6578 (
            .O(N__27993),
            .I(N__27978));
    LocalMux I__6577 (
            .O(N__27990),
            .I(N__27973));
    InMux I__6576 (
            .O(N__27989),
            .I(N__27969));
    LocalMux I__6575 (
            .O(N__27986),
            .I(N__27964));
    Span4Mux_v I__6574 (
            .O(N__27981),
            .I(N__27964));
    LocalMux I__6573 (
            .O(N__27978),
            .I(N__27961));
    InMux I__6572 (
            .O(N__27977),
            .I(N__27958));
    CascadeMux I__6571 (
            .O(N__27976),
            .I(N__27953));
    Span4Mux_v I__6570 (
            .O(N__27973),
            .I(N__27950));
    InMux I__6569 (
            .O(N__27972),
            .I(N__27947));
    LocalMux I__6568 (
            .O(N__27969),
            .I(N__27940));
    Span4Mux_h I__6567 (
            .O(N__27964),
            .I(N__27940));
    Span4Mux_v I__6566 (
            .O(N__27961),
            .I(N__27940));
    LocalMux I__6565 (
            .O(N__27958),
            .I(N__27937));
    InMux I__6564 (
            .O(N__27957),
            .I(N__27934));
    InMux I__6563 (
            .O(N__27956),
            .I(N__27931));
    InMux I__6562 (
            .O(N__27953),
            .I(N__27928));
    Span4Mux_h I__6561 (
            .O(N__27950),
            .I(N__27925));
    LocalMux I__6560 (
            .O(N__27947),
            .I(N__27920));
    Span4Mux_h I__6559 (
            .O(N__27940),
            .I(N__27920));
    Span4Mux_h I__6558 (
            .O(N__27937),
            .I(N__27917));
    LocalMux I__6557 (
            .O(N__27934),
            .I(N__27914));
    LocalMux I__6556 (
            .O(N__27931),
            .I(uart_pc_data_4));
    LocalMux I__6555 (
            .O(N__27928),
            .I(uart_pc_data_4));
    Odrv4 I__6554 (
            .O(N__27925),
            .I(uart_pc_data_4));
    Odrv4 I__6553 (
            .O(N__27920),
            .I(uart_pc_data_4));
    Odrv4 I__6552 (
            .O(N__27917),
            .I(uart_pc_data_4));
    Odrv4 I__6551 (
            .O(N__27914),
            .I(uart_pc_data_4));
    CascadeMux I__6550 (
            .O(N__27901),
            .I(N__27898));
    InMux I__6549 (
            .O(N__27898),
            .I(N__27895));
    LocalMux I__6548 (
            .O(N__27895),
            .I(frame_decoder_OFF3data_4));
    InMux I__6547 (
            .O(N__27892),
            .I(N__27887));
    InMux I__6546 (
            .O(N__27891),
            .I(N__27884));
    InMux I__6545 (
            .O(N__27890),
            .I(N__27880));
    LocalMux I__6544 (
            .O(N__27887),
            .I(N__27875));
    LocalMux I__6543 (
            .O(N__27884),
            .I(N__27875));
    InMux I__6542 (
            .O(N__27883),
            .I(N__27872));
    LocalMux I__6541 (
            .O(N__27880),
            .I(N__27864));
    Span4Mux_v I__6540 (
            .O(N__27875),
            .I(N__27864));
    LocalMux I__6539 (
            .O(N__27872),
            .I(N__27861));
    InMux I__6538 (
            .O(N__27871),
            .I(N__27858));
    InMux I__6537 (
            .O(N__27870),
            .I(N__27854));
    InMux I__6536 (
            .O(N__27869),
            .I(N__27849));
    Span4Mux_h I__6535 (
            .O(N__27864),
            .I(N__27842));
    Span4Mux_v I__6534 (
            .O(N__27861),
            .I(N__27842));
    LocalMux I__6533 (
            .O(N__27858),
            .I(N__27842));
    InMux I__6532 (
            .O(N__27857),
            .I(N__27839));
    LocalMux I__6531 (
            .O(N__27854),
            .I(N__27836));
    InMux I__6530 (
            .O(N__27853),
            .I(N__27833));
    InMux I__6529 (
            .O(N__27852),
            .I(N__27830));
    LocalMux I__6528 (
            .O(N__27849),
            .I(N__27827));
    Span4Mux_h I__6527 (
            .O(N__27842),
            .I(N__27820));
    LocalMux I__6526 (
            .O(N__27839),
            .I(N__27820));
    Span4Mux_v I__6525 (
            .O(N__27836),
            .I(N__27813));
    LocalMux I__6524 (
            .O(N__27833),
            .I(N__27813));
    LocalMux I__6523 (
            .O(N__27830),
            .I(N__27813));
    Span4Mux_v I__6522 (
            .O(N__27827),
            .I(N__27809));
    InMux I__6521 (
            .O(N__27826),
            .I(N__27806));
    InMux I__6520 (
            .O(N__27825),
            .I(N__27803));
    Span4Mux_v I__6519 (
            .O(N__27820),
            .I(N__27800));
    Span4Mux_h I__6518 (
            .O(N__27813),
            .I(N__27797));
    InMux I__6517 (
            .O(N__27812),
            .I(N__27794));
    Odrv4 I__6516 (
            .O(N__27809),
            .I(uart_pc_data_5));
    LocalMux I__6515 (
            .O(N__27806),
            .I(uart_pc_data_5));
    LocalMux I__6514 (
            .O(N__27803),
            .I(uart_pc_data_5));
    Odrv4 I__6513 (
            .O(N__27800),
            .I(uart_pc_data_5));
    Odrv4 I__6512 (
            .O(N__27797),
            .I(uart_pc_data_5));
    LocalMux I__6511 (
            .O(N__27794),
            .I(uart_pc_data_5));
    InMux I__6510 (
            .O(N__27781),
            .I(N__27778));
    LocalMux I__6509 (
            .O(N__27778),
            .I(frame_decoder_OFF3data_5));
    InMux I__6508 (
            .O(N__27775),
            .I(N__27771));
    InMux I__6507 (
            .O(N__27774),
            .I(N__27764));
    LocalMux I__6506 (
            .O(N__27771),
            .I(N__27760));
    InMux I__6505 (
            .O(N__27770),
            .I(N__27757));
    CascadeMux I__6504 (
            .O(N__27769),
            .I(N__27754));
    InMux I__6503 (
            .O(N__27768),
            .I(N__27751));
    InMux I__6502 (
            .O(N__27767),
            .I(N__27748));
    LocalMux I__6501 (
            .O(N__27764),
            .I(N__27745));
    InMux I__6500 (
            .O(N__27763),
            .I(N__27742));
    Span4Mux_v I__6499 (
            .O(N__27760),
            .I(N__27737));
    LocalMux I__6498 (
            .O(N__27757),
            .I(N__27737));
    InMux I__6497 (
            .O(N__27754),
            .I(N__27733));
    LocalMux I__6496 (
            .O(N__27751),
            .I(N__27730));
    LocalMux I__6495 (
            .O(N__27748),
            .I(N__27727));
    Span4Mux_v I__6494 (
            .O(N__27745),
            .I(N__27724));
    LocalMux I__6493 (
            .O(N__27742),
            .I(N__27719));
    Span4Mux_v I__6492 (
            .O(N__27737),
            .I(N__27719));
    InMux I__6491 (
            .O(N__27736),
            .I(N__27715));
    LocalMux I__6490 (
            .O(N__27733),
            .I(N__27710));
    Span4Mux_h I__6489 (
            .O(N__27730),
            .I(N__27707));
    Span4Mux_h I__6488 (
            .O(N__27727),
            .I(N__27704));
    Span4Mux_v I__6487 (
            .O(N__27724),
            .I(N__27699));
    Span4Mux_h I__6486 (
            .O(N__27719),
            .I(N__27699));
    InMux I__6485 (
            .O(N__27718),
            .I(N__27696));
    LocalMux I__6484 (
            .O(N__27715),
            .I(N__27693));
    InMux I__6483 (
            .O(N__27714),
            .I(N__27690));
    InMux I__6482 (
            .O(N__27713),
            .I(N__27687));
    Span4Mux_h I__6481 (
            .O(N__27710),
            .I(N__27684));
    Span4Mux_h I__6480 (
            .O(N__27707),
            .I(N__27679));
    Span4Mux_v I__6479 (
            .O(N__27704),
            .I(N__27679));
    Span4Mux_h I__6478 (
            .O(N__27699),
            .I(N__27674));
    LocalMux I__6477 (
            .O(N__27696),
            .I(N__27674));
    Span4Mux_h I__6476 (
            .O(N__27693),
            .I(N__27669));
    LocalMux I__6475 (
            .O(N__27690),
            .I(N__27669));
    LocalMux I__6474 (
            .O(N__27687),
            .I(uart_pc_data_1));
    Odrv4 I__6473 (
            .O(N__27684),
            .I(uart_pc_data_1));
    Odrv4 I__6472 (
            .O(N__27679),
            .I(uart_pc_data_1));
    Odrv4 I__6471 (
            .O(N__27674),
            .I(uart_pc_data_1));
    Odrv4 I__6470 (
            .O(N__27669),
            .I(uart_pc_data_1));
    CascadeMux I__6469 (
            .O(N__27658),
            .I(N__27655));
    InMux I__6468 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__6467 (
            .O(N__27652),
            .I(frame_decoder_OFF3data_1));
    InMux I__6466 (
            .O(N__27649),
            .I(N__27643));
    InMux I__6465 (
            .O(N__27648),
            .I(N__27640));
    InMux I__6464 (
            .O(N__27647),
            .I(N__27636));
    InMux I__6463 (
            .O(N__27646),
            .I(N__27633));
    LocalMux I__6462 (
            .O(N__27643),
            .I(N__27627));
    LocalMux I__6461 (
            .O(N__27640),
            .I(N__27627));
    InMux I__6460 (
            .O(N__27639),
            .I(N__27624));
    LocalMux I__6459 (
            .O(N__27636),
            .I(N__27618));
    LocalMux I__6458 (
            .O(N__27633),
            .I(N__27614));
    InMux I__6457 (
            .O(N__27632),
            .I(N__27611));
    Span4Mux_v I__6456 (
            .O(N__27627),
            .I(N__27606));
    LocalMux I__6455 (
            .O(N__27624),
            .I(N__27606));
    InMux I__6454 (
            .O(N__27623),
            .I(N__27602));
    InMux I__6453 (
            .O(N__27622),
            .I(N__27599));
    InMux I__6452 (
            .O(N__27621),
            .I(N__27596));
    Span4Mux_v I__6451 (
            .O(N__27618),
            .I(N__27593));
    InMux I__6450 (
            .O(N__27617),
            .I(N__27590));
    Span4Mux_v I__6449 (
            .O(N__27614),
            .I(N__27587));
    LocalMux I__6448 (
            .O(N__27611),
            .I(N__27584));
    Span4Mux_v I__6447 (
            .O(N__27606),
            .I(N__27581));
    InMux I__6446 (
            .O(N__27605),
            .I(N__27578));
    LocalMux I__6445 (
            .O(N__27602),
            .I(N__27572));
    LocalMux I__6444 (
            .O(N__27599),
            .I(N__27572));
    LocalMux I__6443 (
            .O(N__27596),
            .I(N__27569));
    Span4Mux_v I__6442 (
            .O(N__27593),
            .I(N__27564));
    LocalMux I__6441 (
            .O(N__27590),
            .I(N__27564));
    Sp12to4 I__6440 (
            .O(N__27587),
            .I(N__27555));
    Span12Mux_v I__6439 (
            .O(N__27584),
            .I(N__27555));
    Sp12to4 I__6438 (
            .O(N__27581),
            .I(N__27555));
    LocalMux I__6437 (
            .O(N__27578),
            .I(N__27555));
    InMux I__6436 (
            .O(N__27577),
            .I(N__27552));
    Span4Mux_h I__6435 (
            .O(N__27572),
            .I(N__27549));
    Span4Mux_h I__6434 (
            .O(N__27569),
            .I(N__27544));
    Span4Mux_h I__6433 (
            .O(N__27564),
            .I(N__27544));
    Odrv12 I__6432 (
            .O(N__27555),
            .I(uart_pc_data_7));
    LocalMux I__6431 (
            .O(N__27552),
            .I(uart_pc_data_7));
    Odrv4 I__6430 (
            .O(N__27549),
            .I(uart_pc_data_7));
    Odrv4 I__6429 (
            .O(N__27544),
            .I(uart_pc_data_7));
    CascadeMux I__6428 (
            .O(N__27535),
            .I(N__27532));
    InMux I__6427 (
            .O(N__27532),
            .I(N__27526));
    InMux I__6426 (
            .O(N__27531),
            .I(N__27526));
    LocalMux I__6425 (
            .O(N__27526),
            .I(frame_decoder_OFF3data_7));
    InMux I__6424 (
            .O(N__27523),
            .I(N__27520));
    LocalMux I__6423 (
            .O(N__27520),
            .I(\scaler_3.N_533_i_l_ofxZ0 ));
    InMux I__6422 (
            .O(N__27517),
            .I(N__27512));
    CascadeMux I__6421 (
            .O(N__27516),
            .I(N__27509));
    InMux I__6420 (
            .O(N__27515),
            .I(N__27505));
    LocalMux I__6419 (
            .O(N__27512),
            .I(N__27502));
    InMux I__6418 (
            .O(N__27509),
            .I(N__27497));
    InMux I__6417 (
            .O(N__27508),
            .I(N__27497));
    LocalMux I__6416 (
            .O(N__27505),
            .I(\scaler_3.un2_source_data_0 ));
    Odrv12 I__6415 (
            .O(N__27502),
            .I(\scaler_3.un2_source_data_0 ));
    LocalMux I__6414 (
            .O(N__27497),
            .I(\scaler_3.un2_source_data_0 ));
    InMux I__6413 (
            .O(N__27490),
            .I(N__27484));
    InMux I__6412 (
            .O(N__27489),
            .I(N__27481));
    InMux I__6411 (
            .O(N__27488),
            .I(N__27478));
    InMux I__6410 (
            .O(N__27487),
            .I(N__27475));
    LocalMux I__6409 (
            .O(N__27484),
            .I(N__27470));
    LocalMux I__6408 (
            .O(N__27481),
            .I(N__27470));
    LocalMux I__6407 (
            .O(N__27478),
            .I(N__27465));
    LocalMux I__6406 (
            .O(N__27475),
            .I(N__27465));
    Span4Mux_v I__6405 (
            .O(N__27470),
            .I(N__27462));
    Span4Mux_v I__6404 (
            .O(N__27465),
            .I(N__27459));
    Odrv4 I__6403 (
            .O(N__27462),
            .I(frame_decoder_CH3data_0));
    Odrv4 I__6402 (
            .O(N__27459),
            .I(frame_decoder_CH3data_0));
    CascadeMux I__6401 (
            .O(N__27454),
            .I(N__27451));
    InMux I__6400 (
            .O(N__27451),
            .I(N__27448));
    LocalMux I__6399 (
            .O(N__27448),
            .I(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ));
    InMux I__6398 (
            .O(N__27445),
            .I(N__27442));
    LocalMux I__6397 (
            .O(N__27442),
            .I(\scaler_3.un3_source_data_0_axb_7 ));
    InMux I__6396 (
            .O(N__27439),
            .I(N__27436));
    LocalMux I__6395 (
            .O(N__27436),
            .I(N__27433));
    Odrv4 I__6394 (
            .O(N__27433),
            .I(frame_decoder_CH3data_1));
    InMux I__6393 (
            .O(N__27430),
            .I(N__27424));
    InMux I__6392 (
            .O(N__27429),
            .I(N__27424));
    LocalMux I__6391 (
            .O(N__27424),
            .I(frame_decoder_CH3data_7));
    CEMux I__6390 (
            .O(N__27421),
            .I(N__27418));
    LocalMux I__6389 (
            .O(N__27418),
            .I(N__27414));
    CEMux I__6388 (
            .O(N__27417),
            .I(N__27411));
    Span4Mux_v I__6387 (
            .O(N__27414),
            .I(N__27408));
    LocalMux I__6386 (
            .O(N__27411),
            .I(N__27405));
    Span4Mux_v I__6385 (
            .O(N__27408),
            .I(N__27401));
    Span4Mux_h I__6384 (
            .O(N__27405),
            .I(N__27398));
    CEMux I__6383 (
            .O(N__27404),
            .I(N__27395));
    Odrv4 I__6382 (
            .O(N__27401),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    Odrv4 I__6381 (
            .O(N__27398),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    LocalMux I__6380 (
            .O(N__27395),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    CascadeMux I__6379 (
            .O(N__27388),
            .I(N__27384));
    InMux I__6378 (
            .O(N__27387),
            .I(N__27381));
    InMux I__6377 (
            .O(N__27384),
            .I(N__27378));
    LocalMux I__6376 (
            .O(N__27381),
            .I(N__27375));
    LocalMux I__6375 (
            .O(N__27378),
            .I(N__27371));
    Span4Mux_v I__6374 (
            .O(N__27375),
            .I(N__27368));
    InMux I__6373 (
            .O(N__27374),
            .I(N__27365));
    Span4Mux_h I__6372 (
            .O(N__27371),
            .I(N__27362));
    Odrv4 I__6371 (
            .O(N__27368),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__6370 (
            .O(N__27365),
            .I(\Commands_frame_decoder.preinitZ0 ));
    Odrv4 I__6369 (
            .O(N__27362),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__6368 (
            .O(N__27355),
            .I(N__27352));
    LocalMux I__6367 (
            .O(N__27352),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    InMux I__6366 (
            .O(N__27349),
            .I(N__27343));
    InMux I__6365 (
            .O(N__27348),
            .I(N__27338));
    InMux I__6364 (
            .O(N__27347),
            .I(N__27338));
    InMux I__6363 (
            .O(N__27346),
            .I(N__27334));
    LocalMux I__6362 (
            .O(N__27343),
            .I(N__27329));
    LocalMux I__6361 (
            .O(N__27338),
            .I(N__27329));
    CascadeMux I__6360 (
            .O(N__27337),
            .I(N__27326));
    LocalMux I__6359 (
            .O(N__27334),
            .I(N__27323));
    Span4Mux_h I__6358 (
            .O(N__27329),
            .I(N__27320));
    InMux I__6357 (
            .O(N__27326),
            .I(N__27317));
    Span12Mux_v I__6356 (
            .O(N__27323),
            .I(N__27314));
    Odrv4 I__6355 (
            .O(N__27320),
            .I(pc_frame_decoder_dv));
    LocalMux I__6354 (
            .O(N__27317),
            .I(pc_frame_decoder_dv));
    Odrv12 I__6353 (
            .O(N__27314),
            .I(pc_frame_decoder_dv));
    CascadeMux I__6352 (
            .O(N__27307),
            .I(N__27303));
    CascadeMux I__6351 (
            .O(N__27306),
            .I(N__27300));
    InMux I__6350 (
            .O(N__27303),
            .I(N__27292));
    InMux I__6349 (
            .O(N__27300),
            .I(N__27289));
    CascadeMux I__6348 (
            .O(N__27299),
            .I(N__27286));
    InMux I__6347 (
            .O(N__27298),
            .I(N__27283));
    CascadeMux I__6346 (
            .O(N__27297),
            .I(N__27280));
    CascadeMux I__6345 (
            .O(N__27296),
            .I(N__27277));
    InMux I__6344 (
            .O(N__27295),
            .I(N__27261));
    LocalMux I__6343 (
            .O(N__27292),
            .I(N__27258));
    LocalMux I__6342 (
            .O(N__27289),
            .I(N__27255));
    InMux I__6341 (
            .O(N__27286),
            .I(N__27252));
    LocalMux I__6340 (
            .O(N__27283),
            .I(N__27249));
    InMux I__6339 (
            .O(N__27280),
            .I(N__27246));
    InMux I__6338 (
            .O(N__27277),
            .I(N__27243));
    CascadeMux I__6337 (
            .O(N__27276),
            .I(N__27240));
    CascadeMux I__6336 (
            .O(N__27275),
            .I(N__27237));
    CascadeMux I__6335 (
            .O(N__27274),
            .I(N__27234));
    InMux I__6334 (
            .O(N__27273),
            .I(N__27231));
    CascadeMux I__6333 (
            .O(N__27272),
            .I(N__27228));
    CascadeMux I__6332 (
            .O(N__27271),
            .I(N__27225));
    CascadeMux I__6331 (
            .O(N__27270),
            .I(N__27222));
    CascadeMux I__6330 (
            .O(N__27269),
            .I(N__27219));
    CascadeMux I__6329 (
            .O(N__27268),
            .I(N__27216));
    CascadeMux I__6328 (
            .O(N__27267),
            .I(N__27213));
    CascadeMux I__6327 (
            .O(N__27266),
            .I(N__27210));
    CascadeMux I__6326 (
            .O(N__27265),
            .I(N__27203));
    InMux I__6325 (
            .O(N__27264),
            .I(N__27200));
    LocalMux I__6324 (
            .O(N__27261),
            .I(N__27197));
    Span4Mux_h I__6323 (
            .O(N__27258),
            .I(N__27194));
    Span4Mux_v I__6322 (
            .O(N__27255),
            .I(N__27189));
    LocalMux I__6321 (
            .O(N__27252),
            .I(N__27189));
    Span4Mux_h I__6320 (
            .O(N__27249),
            .I(N__27182));
    LocalMux I__6319 (
            .O(N__27246),
            .I(N__27182));
    LocalMux I__6318 (
            .O(N__27243),
            .I(N__27182));
    InMux I__6317 (
            .O(N__27240),
            .I(N__27179));
    InMux I__6316 (
            .O(N__27237),
            .I(N__27176));
    InMux I__6315 (
            .O(N__27234),
            .I(N__27173));
    LocalMux I__6314 (
            .O(N__27231),
            .I(N__27170));
    InMux I__6313 (
            .O(N__27228),
            .I(N__27161));
    InMux I__6312 (
            .O(N__27225),
            .I(N__27161));
    InMux I__6311 (
            .O(N__27222),
            .I(N__27161));
    InMux I__6310 (
            .O(N__27219),
            .I(N__27161));
    InMux I__6309 (
            .O(N__27216),
            .I(N__27154));
    InMux I__6308 (
            .O(N__27213),
            .I(N__27154));
    InMux I__6307 (
            .O(N__27210),
            .I(N__27154));
    CascadeMux I__6306 (
            .O(N__27209),
            .I(N__27151));
    CascadeMux I__6305 (
            .O(N__27208),
            .I(N__27148));
    CascadeMux I__6304 (
            .O(N__27207),
            .I(N__27145));
    CascadeMux I__6303 (
            .O(N__27206),
            .I(N__27142));
    InMux I__6302 (
            .O(N__27203),
            .I(N__27139));
    LocalMux I__6301 (
            .O(N__27200),
            .I(N__27136));
    Span4Mux_v I__6300 (
            .O(N__27197),
            .I(N__27133));
    Span4Mux_v I__6299 (
            .O(N__27194),
            .I(N__27124));
    Span4Mux_h I__6298 (
            .O(N__27189),
            .I(N__27124));
    Span4Mux_h I__6297 (
            .O(N__27182),
            .I(N__27124));
    LocalMux I__6296 (
            .O(N__27179),
            .I(N__27124));
    LocalMux I__6295 (
            .O(N__27176),
            .I(N__27119));
    LocalMux I__6294 (
            .O(N__27173),
            .I(N__27119));
    Span4Mux_v I__6293 (
            .O(N__27170),
            .I(N__27116));
    LocalMux I__6292 (
            .O(N__27161),
            .I(N__27111));
    LocalMux I__6291 (
            .O(N__27154),
            .I(N__27111));
    InMux I__6290 (
            .O(N__27151),
            .I(N__27108));
    InMux I__6289 (
            .O(N__27148),
            .I(N__27103));
    InMux I__6288 (
            .O(N__27145),
            .I(N__27103));
    InMux I__6287 (
            .O(N__27142),
            .I(N__27100));
    LocalMux I__6286 (
            .O(N__27139),
            .I(N__27097));
    Span4Mux_v I__6285 (
            .O(N__27136),
            .I(N__27094));
    Span4Mux_v I__6284 (
            .O(N__27133),
            .I(N__27091));
    Span4Mux_h I__6283 (
            .O(N__27124),
            .I(N__27088));
    Span4Mux_s3_v I__6282 (
            .O(N__27119),
            .I(N__27085));
    Span4Mux_v I__6281 (
            .O(N__27116),
            .I(N__27082));
    Span4Mux_h I__6280 (
            .O(N__27111),
            .I(N__27079));
    LocalMux I__6279 (
            .O(N__27108),
            .I(N__27072));
    LocalMux I__6278 (
            .O(N__27103),
            .I(N__27072));
    LocalMux I__6277 (
            .O(N__27100),
            .I(N__27072));
    Span12Mux_v I__6276 (
            .O(N__27097),
            .I(N__27069));
    Sp12to4 I__6275 (
            .O(N__27094),
            .I(N__27066));
    Span4Mux_v I__6274 (
            .O(N__27091),
            .I(N__27059));
    Span4Mux_v I__6273 (
            .O(N__27088),
            .I(N__27059));
    Span4Mux_v I__6272 (
            .O(N__27085),
            .I(N__27059));
    Span4Mux_h I__6271 (
            .O(N__27082),
            .I(N__27052));
    Span4Mux_v I__6270 (
            .O(N__27079),
            .I(N__27052));
    Span4Mux_v I__6269 (
            .O(N__27072),
            .I(N__27052));
    Odrv12 I__6268 (
            .O(N__27069),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6267 (
            .O(N__27066),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6266 (
            .O(N__27059),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6265 (
            .O(N__27052),
            .I(CONSTANT_ONE_NET));
    InMux I__6264 (
            .O(N__27043),
            .I(N__27039));
    InMux I__6263 (
            .O(N__27042),
            .I(N__27036));
    LocalMux I__6262 (
            .O(N__27039),
            .I(\Commands_frame_decoder.count8_0_i ));
    LocalMux I__6261 (
            .O(N__27036),
            .I(\Commands_frame_decoder.count8_0_i ));
    InMux I__6260 (
            .O(N__27031),
            .I(N__27027));
    InMux I__6259 (
            .O(N__27030),
            .I(N__27024));
    LocalMux I__6258 (
            .O(N__27027),
            .I(\Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0 ));
    LocalMux I__6257 (
            .O(N__27024),
            .I(\Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0 ));
    InMux I__6256 (
            .O(N__27019),
            .I(N__27014));
    InMux I__6255 (
            .O(N__27018),
            .I(N__27009));
    InMux I__6254 (
            .O(N__27017),
            .I(N__27009));
    LocalMux I__6253 (
            .O(N__27014),
            .I(\Commands_frame_decoder.state_1_ns_i_a4_2_0_0 ));
    LocalMux I__6252 (
            .O(N__27009),
            .I(\Commands_frame_decoder.state_1_ns_i_a4_2_0_0 ));
    InMux I__6251 (
            .O(N__27004),
            .I(N__26998));
    InMux I__6250 (
            .O(N__27003),
            .I(N__26995));
    InMux I__6249 (
            .O(N__27002),
            .I(N__26990));
    InMux I__6248 (
            .O(N__27001),
            .I(N__26990));
    LocalMux I__6247 (
            .O(N__26998),
            .I(\Commands_frame_decoder.count8_0 ));
    LocalMux I__6246 (
            .O(N__26995),
            .I(\Commands_frame_decoder.count8_0 ));
    LocalMux I__6245 (
            .O(N__26990),
            .I(\Commands_frame_decoder.count8_0 ));
    InMux I__6244 (
            .O(N__26983),
            .I(N__26980));
    LocalMux I__6243 (
            .O(N__26980),
            .I(frame_decoder_CH3data_2));
    CascadeMux I__6242 (
            .O(N__26977),
            .I(N__26974));
    InMux I__6241 (
            .O(N__26974),
            .I(N__26968));
    InMux I__6240 (
            .O(N__26973),
            .I(N__26968));
    LocalMux I__6239 (
            .O(N__26968),
            .I(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ));
    InMux I__6238 (
            .O(N__26965),
            .I(\scaler_3.un3_source_data_0_cry_1 ));
    InMux I__6237 (
            .O(N__26962),
            .I(N__26959));
    LocalMux I__6236 (
            .O(N__26959),
            .I(frame_decoder_CH3data_3));
    CascadeMux I__6235 (
            .O(N__26956),
            .I(N__26953));
    InMux I__6234 (
            .O(N__26953),
            .I(N__26947));
    InMux I__6233 (
            .O(N__26952),
            .I(N__26947));
    LocalMux I__6232 (
            .O(N__26947),
            .I(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ));
    InMux I__6231 (
            .O(N__26944),
            .I(\scaler_3.un3_source_data_0_cry_2 ));
    InMux I__6230 (
            .O(N__26941),
            .I(N__26938));
    LocalMux I__6229 (
            .O(N__26938),
            .I(frame_decoder_CH3data_4));
    CascadeMux I__6228 (
            .O(N__26935),
            .I(N__26932));
    InMux I__6227 (
            .O(N__26932),
            .I(N__26926));
    InMux I__6226 (
            .O(N__26931),
            .I(N__26926));
    LocalMux I__6225 (
            .O(N__26926),
            .I(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ));
    InMux I__6224 (
            .O(N__26923),
            .I(\scaler_3.un3_source_data_0_cry_3 ));
    CascadeMux I__6223 (
            .O(N__26920),
            .I(N__26917));
    InMux I__6222 (
            .O(N__26917),
            .I(N__26914));
    LocalMux I__6221 (
            .O(N__26914),
            .I(frame_decoder_CH3data_5));
    CascadeMux I__6220 (
            .O(N__26911),
            .I(N__26908));
    InMux I__6219 (
            .O(N__26908),
            .I(N__26902));
    InMux I__6218 (
            .O(N__26907),
            .I(N__26902));
    LocalMux I__6217 (
            .O(N__26902),
            .I(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ));
    InMux I__6216 (
            .O(N__26899),
            .I(\scaler_3.un3_source_data_0_cry_4 ));
    InMux I__6215 (
            .O(N__26896),
            .I(N__26893));
    LocalMux I__6214 (
            .O(N__26893),
            .I(frame_decoder_CH3data_6));
    CascadeMux I__6213 (
            .O(N__26890),
            .I(N__26887));
    InMux I__6212 (
            .O(N__26887),
            .I(N__26881));
    InMux I__6211 (
            .O(N__26886),
            .I(N__26881));
    LocalMux I__6210 (
            .O(N__26881),
            .I(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ));
    InMux I__6209 (
            .O(N__26878),
            .I(\scaler_3.un3_source_data_0_cry_5 ));
    CascadeMux I__6208 (
            .O(N__26875),
            .I(N__26872));
    InMux I__6207 (
            .O(N__26872),
            .I(N__26866));
    InMux I__6206 (
            .O(N__26871),
            .I(N__26866));
    LocalMux I__6205 (
            .O(N__26866),
            .I(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ));
    InMux I__6204 (
            .O(N__26863),
            .I(\scaler_3.un3_source_data_0_cry_6 ));
    InMux I__6203 (
            .O(N__26860),
            .I(N__26856));
    InMux I__6202 (
            .O(N__26859),
            .I(N__26853));
    LocalMux I__6201 (
            .O(N__26856),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    LocalMux I__6200 (
            .O(N__26853),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    InMux I__6199 (
            .O(N__26848),
            .I(bfn_12_16_0_));
    InMux I__6198 (
            .O(N__26845),
            .I(\scaler_3.un3_source_data_0_cry_8 ));
    CascadeMux I__6197 (
            .O(N__26842),
            .I(N__26839));
    InMux I__6196 (
            .O(N__26839),
            .I(N__26836));
    LocalMux I__6195 (
            .O(N__26836),
            .I(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ));
    IoInMux I__6194 (
            .O(N__26833),
            .I(N__26830));
    LocalMux I__6193 (
            .O(N__26830),
            .I(N__26827));
    Odrv4 I__6192 (
            .O(N__26827),
            .I(pc_frame_decoder_dv_0));
    CascadeMux I__6191 (
            .O(N__26824),
            .I(N__26821));
    InMux I__6190 (
            .O(N__26821),
            .I(N__26818));
    LocalMux I__6189 (
            .O(N__26818),
            .I(N__26815));
    Odrv4 I__6188 (
            .O(N__26815),
            .I(frame_decoder_CH4data_1));
    InMux I__6187 (
            .O(N__26812),
            .I(N__26807));
    InMux I__6186 (
            .O(N__26811),
            .I(N__26804));
    InMux I__6185 (
            .O(N__26810),
            .I(N__26801));
    LocalMux I__6184 (
            .O(N__26807),
            .I(N__26794));
    LocalMux I__6183 (
            .O(N__26804),
            .I(N__26794));
    LocalMux I__6182 (
            .O(N__26801),
            .I(N__26794));
    Span4Mux_v I__6181 (
            .O(N__26794),
            .I(N__26790));
    InMux I__6180 (
            .O(N__26793),
            .I(N__26787));
    Odrv4 I__6179 (
            .O(N__26790),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6178 (
            .O(N__26787),
            .I(frame_decoder_CH4data_0));
    CEMux I__6177 (
            .O(N__26782),
            .I(N__26778));
    CEMux I__6176 (
            .O(N__26781),
            .I(N__26775));
    LocalMux I__6175 (
            .O(N__26778),
            .I(N__26770));
    LocalMux I__6174 (
            .O(N__26775),
            .I(N__26767));
    CEMux I__6173 (
            .O(N__26774),
            .I(N__26764));
    CEMux I__6172 (
            .O(N__26773),
            .I(N__26761));
    Span4Mux_v I__6171 (
            .O(N__26770),
            .I(N__26754));
    Span4Mux_h I__6170 (
            .O(N__26767),
            .I(N__26754));
    LocalMux I__6169 (
            .O(N__26764),
            .I(N__26754));
    LocalMux I__6168 (
            .O(N__26761),
            .I(N__26751));
    Span4Mux_h I__6167 (
            .O(N__26754),
            .I(N__26748));
    Span4Mux_v I__6166 (
            .O(N__26751),
            .I(N__26745));
    Odrv4 I__6165 (
            .O(N__26748),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    Odrv4 I__6164 (
            .O(N__26745),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__6163 (
            .O(N__26740),
            .I(\scaler_3.un3_source_data_0_cry_0 ));
    InMux I__6162 (
            .O(N__26737),
            .I(N__26734));
    LocalMux I__6161 (
            .O(N__26734),
            .I(N__26731));
    Odrv4 I__6160 (
            .O(N__26731),
            .I(\uart_drone.CO0 ));
    InMux I__6159 (
            .O(N__26728),
            .I(N__26725));
    LocalMux I__6158 (
            .O(N__26725),
            .I(\Commands_frame_decoder.count8_axb_1 ));
    InMux I__6157 (
            .O(N__26722),
            .I(N__26719));
    LocalMux I__6156 (
            .O(N__26719),
            .I(\Commands_frame_decoder.count_i_2 ));
    InMux I__6155 (
            .O(N__26716),
            .I(\Commands_frame_decoder.count8 ));
    InMux I__6154 (
            .O(N__26713),
            .I(N__26710));
    LocalMux I__6153 (
            .O(N__26710),
            .I(\Commands_frame_decoder.count8_THRU_CO ));
    InMux I__6152 (
            .O(N__26707),
            .I(N__26704));
    LocalMux I__6151 (
            .O(N__26704),
            .I(N__26701));
    Span4Mux_v I__6150 (
            .O(N__26701),
            .I(N__26698));
    Span4Mux_v I__6149 (
            .O(N__26698),
            .I(N__26688));
    InMux I__6148 (
            .O(N__26697),
            .I(N__26680));
    InMux I__6147 (
            .O(N__26696),
            .I(N__26676));
    InMux I__6146 (
            .O(N__26695),
            .I(N__26671));
    InMux I__6145 (
            .O(N__26694),
            .I(N__26671));
    InMux I__6144 (
            .O(N__26693),
            .I(N__26664));
    InMux I__6143 (
            .O(N__26692),
            .I(N__26664));
    InMux I__6142 (
            .O(N__26691),
            .I(N__26664));
    Span4Mux_v I__6141 (
            .O(N__26688),
            .I(N__26661));
    InMux I__6140 (
            .O(N__26687),
            .I(N__26658));
    InMux I__6139 (
            .O(N__26686),
            .I(N__26648));
    InMux I__6138 (
            .O(N__26685),
            .I(N__26648));
    InMux I__6137 (
            .O(N__26684),
            .I(N__26648));
    InMux I__6136 (
            .O(N__26683),
            .I(N__26648));
    LocalMux I__6135 (
            .O(N__26680),
            .I(N__26643));
    IoInMux I__6134 (
            .O(N__26679),
            .I(N__26639));
    LocalMux I__6133 (
            .O(N__26676),
            .I(N__26632));
    LocalMux I__6132 (
            .O(N__26671),
            .I(N__26632));
    LocalMux I__6131 (
            .O(N__26664),
            .I(N__26632));
    Span4Mux_h I__6130 (
            .O(N__26661),
            .I(N__26627));
    LocalMux I__6129 (
            .O(N__26658),
            .I(N__26627));
    InMux I__6128 (
            .O(N__26657),
            .I(N__26618));
    LocalMux I__6127 (
            .O(N__26648),
            .I(N__26615));
    InMux I__6126 (
            .O(N__26647),
            .I(N__26612));
    InMux I__6125 (
            .O(N__26646),
            .I(N__26609));
    Span4Mux_h I__6124 (
            .O(N__26643),
            .I(N__26605));
    InMux I__6123 (
            .O(N__26642),
            .I(N__26602));
    LocalMux I__6122 (
            .O(N__26639),
            .I(N__26599));
    Span4Mux_v I__6121 (
            .O(N__26632),
            .I(N__26596));
    Span4Mux_v I__6120 (
            .O(N__26627),
            .I(N__26593));
    InMux I__6119 (
            .O(N__26626),
            .I(N__26590));
    InMux I__6118 (
            .O(N__26625),
            .I(N__26585));
    InMux I__6117 (
            .O(N__26624),
            .I(N__26585));
    InMux I__6116 (
            .O(N__26623),
            .I(N__26578));
    InMux I__6115 (
            .O(N__26622),
            .I(N__26578));
    InMux I__6114 (
            .O(N__26621),
            .I(N__26578));
    LocalMux I__6113 (
            .O(N__26618),
            .I(N__26575));
    Span4Mux_h I__6112 (
            .O(N__26615),
            .I(N__26568));
    LocalMux I__6111 (
            .O(N__26612),
            .I(N__26568));
    LocalMux I__6110 (
            .O(N__26609),
            .I(N__26568));
    InMux I__6109 (
            .O(N__26608),
            .I(N__26565));
    Sp12to4 I__6108 (
            .O(N__26605),
            .I(N__26560));
    LocalMux I__6107 (
            .O(N__26602),
            .I(N__26560));
    Span4Mux_s1_v I__6106 (
            .O(N__26599),
            .I(N__26557));
    Span4Mux_v I__6105 (
            .O(N__26596),
            .I(N__26552));
    Span4Mux_v I__6104 (
            .O(N__26593),
            .I(N__26552));
    LocalMux I__6103 (
            .O(N__26590),
            .I(N__26537));
    LocalMux I__6102 (
            .O(N__26585),
            .I(N__26537));
    LocalMux I__6101 (
            .O(N__26578),
            .I(N__26537));
    Span12Mux_h I__6100 (
            .O(N__26575),
            .I(N__26537));
    Sp12to4 I__6099 (
            .O(N__26568),
            .I(N__26537));
    LocalMux I__6098 (
            .O(N__26565),
            .I(N__26537));
    Span12Mux_s11_v I__6097 (
            .O(N__26560),
            .I(N__26537));
    Span4Mux_v I__6096 (
            .O(N__26557),
            .I(N__26534));
    Odrv4 I__6095 (
            .O(N__26552),
            .I(reset_system));
    Odrv12 I__6094 (
            .O(N__26537),
            .I(reset_system));
    Odrv4 I__6093 (
            .O(N__26534),
            .I(reset_system));
    CascadeMux I__6092 (
            .O(N__26527),
            .I(\Commands_frame_decoder.count8_THRU_CO_cascade_ ));
    CascadeMux I__6091 (
            .O(N__26524),
            .I(\Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_ ));
    InMux I__6090 (
            .O(N__26521),
            .I(N__26516));
    InMux I__6089 (
            .O(N__26520),
            .I(N__26511));
    InMux I__6088 (
            .O(N__26519),
            .I(N__26511));
    LocalMux I__6087 (
            .O(N__26516),
            .I(\Commands_frame_decoder.countZ0Z_2 ));
    LocalMux I__6086 (
            .O(N__26511),
            .I(\Commands_frame_decoder.countZ0Z_2 ));
    InMux I__6085 (
            .O(N__26506),
            .I(N__26503));
    LocalMux I__6084 (
            .O(N__26503),
            .I(\Commands_frame_decoder.CO0 ));
    CascadeMux I__6083 (
            .O(N__26500),
            .I(\Commands_frame_decoder.CO0_cascade_ ));
    InMux I__6082 (
            .O(N__26497),
            .I(N__26491));
    InMux I__6081 (
            .O(N__26496),
            .I(N__26484));
    InMux I__6080 (
            .O(N__26495),
            .I(N__26484));
    InMux I__6079 (
            .O(N__26494),
            .I(N__26484));
    LocalMux I__6078 (
            .O(N__26491),
            .I(\Commands_frame_decoder.countZ0Z_1 ));
    LocalMux I__6077 (
            .O(N__26484),
            .I(\Commands_frame_decoder.countZ0Z_1 ));
    InMux I__6076 (
            .O(N__26479),
            .I(N__26475));
    InMux I__6075 (
            .O(N__26478),
            .I(N__26472));
    LocalMux I__6074 (
            .O(N__26475),
            .I(N__26469));
    LocalMux I__6073 (
            .O(N__26472),
            .I(N__26466));
    Span12Mux_v I__6072 (
            .O(N__26469),
            .I(N__26463));
    Span4Mux_h I__6071 (
            .O(N__26466),
            .I(N__26460));
    Odrv12 I__6070 (
            .O(N__26463),
            .I(scaler_3_data_11));
    Odrv4 I__6069 (
            .O(N__26460),
            .I(scaler_3_data_11));
    InMux I__6068 (
            .O(N__26455),
            .I(\scaler_3.un2_source_data_0_cry_6 ));
    InMux I__6067 (
            .O(N__26452),
            .I(N__26448));
    InMux I__6066 (
            .O(N__26451),
            .I(N__26445));
    LocalMux I__6065 (
            .O(N__26448),
            .I(N__26442));
    LocalMux I__6064 (
            .O(N__26445),
            .I(N__26439));
    Span12Mux_v I__6063 (
            .O(N__26442),
            .I(N__26436));
    Span4Mux_h I__6062 (
            .O(N__26439),
            .I(N__26433));
    Odrv12 I__6061 (
            .O(N__26436),
            .I(scaler_3_data_12));
    Odrv4 I__6060 (
            .O(N__26433),
            .I(scaler_3_data_12));
    InMux I__6059 (
            .O(N__26428),
            .I(\scaler_3.un2_source_data_0_cry_7 ));
    InMux I__6058 (
            .O(N__26425),
            .I(N__26422));
    LocalMux I__6057 (
            .O(N__26422),
            .I(N__26418));
    InMux I__6056 (
            .O(N__26421),
            .I(N__26415));
    Span4Mux_h I__6055 (
            .O(N__26418),
            .I(N__26412));
    LocalMux I__6054 (
            .O(N__26415),
            .I(N__26409));
    Span4Mux_v I__6053 (
            .O(N__26412),
            .I(N__26406));
    Span4Mux_h I__6052 (
            .O(N__26409),
            .I(N__26403));
    Odrv4 I__6051 (
            .O(N__26406),
            .I(scaler_3_data_13));
    Odrv4 I__6050 (
            .O(N__26403),
            .I(scaler_3_data_13));
    InMux I__6049 (
            .O(N__26398),
            .I(bfn_11_17_0_));
    InMux I__6048 (
            .O(N__26395),
            .I(\scaler_3.un2_source_data_0_cry_9 ));
    InMux I__6047 (
            .O(N__26392),
            .I(N__26389));
    LocalMux I__6046 (
            .O(N__26389),
            .I(N__26386));
    Span4Mux_v I__6045 (
            .O(N__26386),
            .I(N__26383));
    Odrv4 I__6044 (
            .O(N__26383),
            .I(scaler_3_data_14));
    CEMux I__6043 (
            .O(N__26380),
            .I(N__26359));
    CEMux I__6042 (
            .O(N__26379),
            .I(N__26359));
    CEMux I__6041 (
            .O(N__26378),
            .I(N__26359));
    CEMux I__6040 (
            .O(N__26377),
            .I(N__26359));
    CEMux I__6039 (
            .O(N__26376),
            .I(N__26359));
    CEMux I__6038 (
            .O(N__26375),
            .I(N__26359));
    CEMux I__6037 (
            .O(N__26374),
            .I(N__26359));
    GlobalMux I__6036 (
            .O(N__26359),
            .I(N__26356));
    gio2CtrlBuf I__6035 (
            .O(N__26356),
            .I(pc_frame_decoder_dv_0_g));
    InMux I__6034 (
            .O(N__26353),
            .I(N__26350));
    LocalMux I__6033 (
            .O(N__26350),
            .I(N__26345));
    InMux I__6032 (
            .O(N__26349),
            .I(N__26342));
    InMux I__6031 (
            .O(N__26348),
            .I(N__26337));
    Span4Mux_v I__6030 (
            .O(N__26345),
            .I(N__26329));
    LocalMux I__6029 (
            .O(N__26342),
            .I(N__26329));
    InMux I__6028 (
            .O(N__26341),
            .I(N__26326));
    InMux I__6027 (
            .O(N__26340),
            .I(N__26323));
    LocalMux I__6026 (
            .O(N__26337),
            .I(N__26320));
    CascadeMux I__6025 (
            .O(N__26336),
            .I(N__26317));
    InMux I__6024 (
            .O(N__26335),
            .I(N__26314));
    InMux I__6023 (
            .O(N__26334),
            .I(N__26310));
    Span4Mux_h I__6022 (
            .O(N__26329),
            .I(N__26301));
    LocalMux I__6021 (
            .O(N__26326),
            .I(N__26301));
    LocalMux I__6020 (
            .O(N__26323),
            .I(N__26301));
    Span4Mux_h I__6019 (
            .O(N__26320),
            .I(N__26301));
    InMux I__6018 (
            .O(N__26317),
            .I(N__26298));
    LocalMux I__6017 (
            .O(N__26314),
            .I(N__26295));
    InMux I__6016 (
            .O(N__26313),
            .I(N__26292));
    LocalMux I__6015 (
            .O(N__26310),
            .I(N__26287));
    Span4Mux_v I__6014 (
            .O(N__26301),
            .I(N__26287));
    LocalMux I__6013 (
            .O(N__26298),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv12 I__6012 (
            .O(N__26295),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__6011 (
            .O(N__26292),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__6010 (
            .O(N__26287),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__6009 (
            .O(N__26278),
            .I(N__26275));
    LocalMux I__6008 (
            .O(N__26275),
            .I(N__26268));
    InMux I__6007 (
            .O(N__26274),
            .I(N__26265));
    InMux I__6006 (
            .O(N__26273),
            .I(N__26260));
    InMux I__6005 (
            .O(N__26272),
            .I(N__26257));
    InMux I__6004 (
            .O(N__26271),
            .I(N__26254));
    Span4Mux_h I__6003 (
            .O(N__26268),
            .I(N__26247));
    LocalMux I__6002 (
            .O(N__26265),
            .I(N__26247));
    InMux I__6001 (
            .O(N__26264),
            .I(N__26244));
    InMux I__6000 (
            .O(N__26263),
            .I(N__26240));
    LocalMux I__5999 (
            .O(N__26260),
            .I(N__26233));
    LocalMux I__5998 (
            .O(N__26257),
            .I(N__26233));
    LocalMux I__5997 (
            .O(N__26254),
            .I(N__26233));
    InMux I__5996 (
            .O(N__26253),
            .I(N__26228));
    InMux I__5995 (
            .O(N__26252),
            .I(N__26228));
    Sp12to4 I__5994 (
            .O(N__26247),
            .I(N__26223));
    LocalMux I__5993 (
            .O(N__26244),
            .I(N__26223));
    InMux I__5992 (
            .O(N__26243),
            .I(N__26220));
    LocalMux I__5991 (
            .O(N__26240),
            .I(N__26215));
    Span12Mux_v I__5990 (
            .O(N__26233),
            .I(N__26215));
    LocalMux I__5989 (
            .O(N__26228),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__5988 (
            .O(N__26223),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__5987 (
            .O(N__26220),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__5986 (
            .O(N__26215),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__5985 (
            .O(N__26206),
            .I(N__26203));
    LocalMux I__5984 (
            .O(N__26203),
            .I(N__26200));
    Span4Mux_h I__5983 (
            .O(N__26200),
            .I(N__26197));
    Odrv4 I__5982 (
            .O(N__26197),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__5981 (
            .O(N__26194),
            .I(N__26188));
    InMux I__5980 (
            .O(N__26193),
            .I(N__26188));
    LocalMux I__5979 (
            .O(N__26188),
            .I(N__26185));
    Span4Mux_h I__5978 (
            .O(N__26185),
            .I(N__26180));
    InMux I__5977 (
            .O(N__26184),
            .I(N__26175));
    InMux I__5976 (
            .O(N__26183),
            .I(N__26175));
    Odrv4 I__5975 (
            .O(N__26180),
            .I(\Commands_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__5974 (
            .O(N__26175),
            .I(\Commands_frame_decoder.state_1Z0Z_10 ));
    CascadeMux I__5973 (
            .O(N__26170),
            .I(\Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_ ));
    CascadeMux I__5972 (
            .O(N__26167),
            .I(N__26164));
    InMux I__5971 (
            .O(N__26164),
            .I(N__26158));
    InMux I__5970 (
            .O(N__26163),
            .I(N__26158));
    LocalMux I__5969 (
            .O(N__26158),
            .I(N__26155));
    Span4Mux_h I__5968 (
            .O(N__26155),
            .I(N__26152));
    Odrv4 I__5967 (
            .O(N__26152),
            .I(\Commands_frame_decoder.N_292 ));
    CascadeMux I__5966 (
            .O(N__26149),
            .I(N__26144));
    InMux I__5965 (
            .O(N__26148),
            .I(N__26141));
    InMux I__5964 (
            .O(N__26147),
            .I(N__26138));
    InMux I__5963 (
            .O(N__26144),
            .I(N__26134));
    LocalMux I__5962 (
            .O(N__26141),
            .I(N__26131));
    LocalMux I__5961 (
            .O(N__26138),
            .I(N__26128));
    InMux I__5960 (
            .O(N__26137),
            .I(N__26125));
    LocalMux I__5959 (
            .O(N__26134),
            .I(N__26116));
    Span4Mux_v I__5958 (
            .O(N__26131),
            .I(N__26116));
    Span4Mux_h I__5957 (
            .O(N__26128),
            .I(N__26116));
    LocalMux I__5956 (
            .O(N__26125),
            .I(N__26116));
    Odrv4 I__5955 (
            .O(N__26116),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__5954 (
            .O(N__26113),
            .I(N__26105));
    InMux I__5953 (
            .O(N__26112),
            .I(N__26102));
    InMux I__5952 (
            .O(N__26111),
            .I(N__26099));
    InMux I__5951 (
            .O(N__26110),
            .I(N__26096));
    InMux I__5950 (
            .O(N__26109),
            .I(N__26091));
    InMux I__5949 (
            .O(N__26108),
            .I(N__26087));
    LocalMux I__5948 (
            .O(N__26105),
            .I(N__26082));
    LocalMux I__5947 (
            .O(N__26102),
            .I(N__26082));
    LocalMux I__5946 (
            .O(N__26099),
            .I(N__26077));
    LocalMux I__5945 (
            .O(N__26096),
            .I(N__26077));
    InMux I__5944 (
            .O(N__26095),
            .I(N__26074));
    InMux I__5943 (
            .O(N__26094),
            .I(N__26069));
    LocalMux I__5942 (
            .O(N__26091),
            .I(N__26066));
    InMux I__5941 (
            .O(N__26090),
            .I(N__26063));
    LocalMux I__5940 (
            .O(N__26087),
            .I(N__26058));
    Span4Mux_v I__5939 (
            .O(N__26082),
            .I(N__26058));
    Span4Mux_v I__5938 (
            .O(N__26077),
            .I(N__26053));
    LocalMux I__5937 (
            .O(N__26074),
            .I(N__26053));
    InMux I__5936 (
            .O(N__26073),
            .I(N__26048));
    InMux I__5935 (
            .O(N__26072),
            .I(N__26048));
    LocalMux I__5934 (
            .O(N__26069),
            .I(N__26043));
    Span4Mux_h I__5933 (
            .O(N__26066),
            .I(N__26043));
    LocalMux I__5932 (
            .O(N__26063),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__5931 (
            .O(N__26058),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__5930 (
            .O(N__26053),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__5929 (
            .O(N__26048),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__5928 (
            .O(N__26043),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__5927 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__5926 (
            .O(N__26029),
            .I(N__26026));
    Odrv4 I__5925 (
            .O(N__26026),
            .I(\scaler_4.N_545_i_l_ofxZ0 ));
    InMux I__5924 (
            .O(N__26023),
            .I(N__26019));
    InMux I__5923 (
            .O(N__26022),
            .I(N__26016));
    LocalMux I__5922 (
            .O(N__26019),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__5921 (
            .O(N__26016),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    InMux I__5920 (
            .O(N__26011),
            .I(bfn_11_15_0_));
    InMux I__5919 (
            .O(N__26008),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CascadeMux I__5918 (
            .O(N__26005),
            .I(N__26002));
    InMux I__5917 (
            .O(N__26002),
            .I(N__25999));
    LocalMux I__5916 (
            .O(N__25999),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__5915 (
            .O(N__25996),
            .I(N__25993));
    LocalMux I__5914 (
            .O(N__25993),
            .I(N__25990));
    Span4Mux_v I__5913 (
            .O(N__25990),
            .I(N__25987));
    Span4Mux_h I__5912 (
            .O(N__25987),
            .I(N__25983));
    InMux I__5911 (
            .O(N__25986),
            .I(N__25980));
    Span4Mux_h I__5910 (
            .O(N__25983),
            .I(N__25975));
    LocalMux I__5909 (
            .O(N__25980),
            .I(N__25975));
    Span4Mux_v I__5908 (
            .O(N__25975),
            .I(N__25972));
    Odrv4 I__5907 (
            .O(N__25972),
            .I(scaler_3_data_6));
    InMux I__5906 (
            .O(N__25969),
            .I(\scaler_3.un2_source_data_0_cry_1 ));
    InMux I__5905 (
            .O(N__25966),
            .I(N__25963));
    LocalMux I__5904 (
            .O(N__25963),
            .I(N__25960));
    Span4Mux_v I__5903 (
            .O(N__25960),
            .I(N__25956));
    InMux I__5902 (
            .O(N__25959),
            .I(N__25953));
    Span4Mux_h I__5901 (
            .O(N__25956),
            .I(N__25948));
    LocalMux I__5900 (
            .O(N__25953),
            .I(N__25948));
    Span4Mux_h I__5899 (
            .O(N__25948),
            .I(N__25945));
    Odrv4 I__5898 (
            .O(N__25945),
            .I(scaler_3_data_7));
    InMux I__5897 (
            .O(N__25942),
            .I(\scaler_3.un2_source_data_0_cry_2 ));
    InMux I__5896 (
            .O(N__25939),
            .I(N__25936));
    LocalMux I__5895 (
            .O(N__25936),
            .I(N__25932));
    InMux I__5894 (
            .O(N__25935),
            .I(N__25929));
    Span4Mux_v I__5893 (
            .O(N__25932),
            .I(N__25924));
    LocalMux I__5892 (
            .O(N__25929),
            .I(N__25924));
    Span4Mux_h I__5891 (
            .O(N__25924),
            .I(N__25921));
    Odrv4 I__5890 (
            .O(N__25921),
            .I(scaler_3_data_8));
    InMux I__5889 (
            .O(N__25918),
            .I(\scaler_3.un2_source_data_0_cry_3 ));
    InMux I__5888 (
            .O(N__25915),
            .I(N__25912));
    LocalMux I__5887 (
            .O(N__25912),
            .I(N__25908));
    InMux I__5886 (
            .O(N__25911),
            .I(N__25905));
    Span4Mux_v I__5885 (
            .O(N__25908),
            .I(N__25902));
    LocalMux I__5884 (
            .O(N__25905),
            .I(N__25899));
    Span4Mux_h I__5883 (
            .O(N__25902),
            .I(N__25894));
    Span4Mux_h I__5882 (
            .O(N__25899),
            .I(N__25894));
    Odrv4 I__5881 (
            .O(N__25894),
            .I(scaler_3_data_9));
    InMux I__5880 (
            .O(N__25891),
            .I(\scaler_3.un2_source_data_0_cry_4 ));
    InMux I__5879 (
            .O(N__25888),
            .I(N__25884));
    InMux I__5878 (
            .O(N__25887),
            .I(N__25881));
    LocalMux I__5877 (
            .O(N__25884),
            .I(N__25878));
    LocalMux I__5876 (
            .O(N__25881),
            .I(N__25875));
    Span12Mux_s11_h I__5875 (
            .O(N__25878),
            .I(N__25872));
    Span4Mux_h I__5874 (
            .O(N__25875),
            .I(N__25869));
    Odrv12 I__5873 (
            .O(N__25872),
            .I(scaler_3_data_10));
    Odrv4 I__5872 (
            .O(N__25869),
            .I(scaler_3_data_10));
    InMux I__5871 (
            .O(N__25864),
            .I(\scaler_3.un2_source_data_0_cry_5 ));
    InMux I__5870 (
            .O(N__25861),
            .I(N__25857));
    InMux I__5869 (
            .O(N__25860),
            .I(N__25853));
    LocalMux I__5868 (
            .O(N__25857),
            .I(N__25849));
    CascadeMux I__5867 (
            .O(N__25856),
            .I(N__25846));
    LocalMux I__5866 (
            .O(N__25853),
            .I(N__25843));
    InMux I__5865 (
            .O(N__25852),
            .I(N__25840));
    Span4Mux_v I__5864 (
            .O(N__25849),
            .I(N__25837));
    InMux I__5863 (
            .O(N__25846),
            .I(N__25834));
    Odrv4 I__5862 (
            .O(N__25843),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__5861 (
            .O(N__25840),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__5860 (
            .O(N__25837),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__5859 (
            .O(N__25834),
            .I(frame_decoder_OFF4data_0));
    InMux I__5858 (
            .O(N__25825),
            .I(N__25822));
    LocalMux I__5857 (
            .O(N__25822),
            .I(frame_decoder_OFF4data_1));
    InMux I__5856 (
            .O(N__25819),
            .I(N__25815));
    InMux I__5855 (
            .O(N__25818),
            .I(N__25812));
    LocalMux I__5854 (
            .O(N__25815),
            .I(N__25806));
    LocalMux I__5853 (
            .O(N__25812),
            .I(N__25806));
    CascadeMux I__5852 (
            .O(N__25811),
            .I(N__25803));
    Span4Mux_h I__5851 (
            .O(N__25806),
            .I(N__25799));
    InMux I__5850 (
            .O(N__25803),
            .I(N__25794));
    InMux I__5849 (
            .O(N__25802),
            .I(N__25794));
    Odrv4 I__5848 (
            .O(N__25799),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__5847 (
            .O(N__25794),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__5846 (
            .O(N__25789),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__5845 (
            .O(N__25786),
            .I(N__25783));
    LocalMux I__5844 (
            .O(N__25783),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__5843 (
            .O(N__25780),
            .I(N__25777));
    InMux I__5842 (
            .O(N__25777),
            .I(N__25774));
    LocalMux I__5841 (
            .O(N__25774),
            .I(frame_decoder_OFF4data_2));
    CascadeMux I__5840 (
            .O(N__25771),
            .I(N__25768));
    InMux I__5839 (
            .O(N__25768),
            .I(N__25762));
    InMux I__5838 (
            .O(N__25767),
            .I(N__25762));
    LocalMux I__5837 (
            .O(N__25762),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__5836 (
            .O(N__25759),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__5835 (
            .O(N__25756),
            .I(N__25753));
    LocalMux I__5834 (
            .O(N__25753),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__5833 (
            .O(N__25750),
            .I(N__25747));
    InMux I__5832 (
            .O(N__25747),
            .I(N__25741));
    InMux I__5831 (
            .O(N__25746),
            .I(N__25741));
    LocalMux I__5830 (
            .O(N__25741),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__5829 (
            .O(N__25738),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__5828 (
            .O(N__25735),
            .I(N__25732));
    LocalMux I__5827 (
            .O(N__25732),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__5826 (
            .O(N__25729),
            .I(N__25726));
    InMux I__5825 (
            .O(N__25726),
            .I(N__25723));
    LocalMux I__5824 (
            .O(N__25723),
            .I(N__25720));
    Odrv4 I__5823 (
            .O(N__25720),
            .I(frame_decoder_OFF4data_4));
    CascadeMux I__5822 (
            .O(N__25717),
            .I(N__25714));
    InMux I__5821 (
            .O(N__25714),
            .I(N__25708));
    InMux I__5820 (
            .O(N__25713),
            .I(N__25708));
    LocalMux I__5819 (
            .O(N__25708),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__5818 (
            .O(N__25705),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__5817 (
            .O(N__25702),
            .I(N__25699));
    LocalMux I__5816 (
            .O(N__25699),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__5815 (
            .O(N__25696),
            .I(N__25693));
    InMux I__5814 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__5813 (
            .O(N__25690),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__5812 (
            .O(N__25687),
            .I(N__25684));
    InMux I__5811 (
            .O(N__25684),
            .I(N__25678));
    InMux I__5810 (
            .O(N__25683),
            .I(N__25678));
    LocalMux I__5809 (
            .O(N__25678),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__5808 (
            .O(N__25675),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__5807 (
            .O(N__25672),
            .I(N__25669));
    LocalMux I__5806 (
            .O(N__25669),
            .I(N__25666));
    Odrv4 I__5805 (
            .O(N__25666),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__5804 (
            .O(N__25663),
            .I(N__25660));
    InMux I__5803 (
            .O(N__25660),
            .I(N__25654));
    InMux I__5802 (
            .O(N__25659),
            .I(N__25654));
    LocalMux I__5801 (
            .O(N__25654),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__5800 (
            .O(N__25651),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__5799 (
            .O(N__25648),
            .I(N__25645));
    LocalMux I__5798 (
            .O(N__25645),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    CascadeMux I__5797 (
            .O(N__25642),
            .I(N__25639));
    InMux I__5796 (
            .O(N__25639),
            .I(N__25633));
    InMux I__5795 (
            .O(N__25638),
            .I(N__25633));
    LocalMux I__5794 (
            .O(N__25633),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__5793 (
            .O(N__25630),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    CascadeMux I__5792 (
            .O(N__25627),
            .I(N__25624));
    InMux I__5791 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__5790 (
            .O(N__25621),
            .I(N__25618));
    Span4Mux_v I__5789 (
            .O(N__25618),
            .I(N__25613));
    CascadeMux I__5788 (
            .O(N__25617),
            .I(N__25609));
    InMux I__5787 (
            .O(N__25616),
            .I(N__25606));
    Span4Mux_h I__5786 (
            .O(N__25613),
            .I(N__25603));
    InMux I__5785 (
            .O(N__25612),
            .I(N__25598));
    InMux I__5784 (
            .O(N__25609),
            .I(N__25598));
    LocalMux I__5783 (
            .O(N__25606),
            .I(N__25595));
    Odrv4 I__5782 (
            .O(N__25603),
            .I(\Commands_frame_decoder.state_1Z0Z_6 ));
    LocalMux I__5781 (
            .O(N__25598),
            .I(\Commands_frame_decoder.state_1Z0Z_6 ));
    Odrv4 I__5780 (
            .O(N__25595),
            .I(\Commands_frame_decoder.state_1Z0Z_6 ));
    CascadeMux I__5779 (
            .O(N__25588),
            .I(N__25584));
    InMux I__5778 (
            .O(N__25587),
            .I(N__25579));
    InMux I__5777 (
            .O(N__25584),
            .I(N__25575));
    CascadeMux I__5776 (
            .O(N__25583),
            .I(N__25572));
    InMux I__5775 (
            .O(N__25582),
            .I(N__25568));
    LocalMux I__5774 (
            .O(N__25579),
            .I(N__25563));
    CascadeMux I__5773 (
            .O(N__25578),
            .I(N__25560));
    LocalMux I__5772 (
            .O(N__25575),
            .I(N__25557));
    InMux I__5771 (
            .O(N__25572),
            .I(N__25552));
    InMux I__5770 (
            .O(N__25571),
            .I(N__25552));
    LocalMux I__5769 (
            .O(N__25568),
            .I(N__25549));
    InMux I__5768 (
            .O(N__25567),
            .I(N__25544));
    InMux I__5767 (
            .O(N__25566),
            .I(N__25544));
    Span4Mux_h I__5766 (
            .O(N__25563),
            .I(N__25541));
    InMux I__5765 (
            .O(N__25560),
            .I(N__25538));
    Odrv12 I__5764 (
            .O(N__25557),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__5763 (
            .O(N__25552),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__5762 (
            .O(N__25549),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__5761 (
            .O(N__25544),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__5760 (
            .O(N__25541),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__5759 (
            .O(N__25538),
            .I(\uart_drone.stateZ0Z_3 ));
    InMux I__5758 (
            .O(N__25525),
            .I(N__25519));
    InMux I__5757 (
            .O(N__25524),
            .I(N__25516));
    InMux I__5756 (
            .O(N__25523),
            .I(N__25513));
    InMux I__5755 (
            .O(N__25522),
            .I(N__25510));
    LocalMux I__5754 (
            .O(N__25519),
            .I(N__25507));
    LocalMux I__5753 (
            .O(N__25516),
            .I(N__25502));
    LocalMux I__5752 (
            .O(N__25513),
            .I(N__25502));
    LocalMux I__5751 (
            .O(N__25510),
            .I(N__25499));
    Span4Mux_v I__5750 (
            .O(N__25507),
            .I(N__25494));
    Span4Mux_v I__5749 (
            .O(N__25502),
            .I(N__25494));
    Odrv4 I__5748 (
            .O(N__25499),
            .I(\uart_drone.N_152 ));
    Odrv4 I__5747 (
            .O(N__25494),
            .I(\uart_drone.N_152 ));
    InMux I__5746 (
            .O(N__25489),
            .I(N__25483));
    InMux I__5745 (
            .O(N__25488),
            .I(N__25483));
    LocalMux I__5744 (
            .O(N__25483),
            .I(\uart_drone.un1_state_7_0 ));
    InMux I__5743 (
            .O(N__25480),
            .I(N__25476));
    InMux I__5742 (
            .O(N__25479),
            .I(N__25473));
    LocalMux I__5741 (
            .O(N__25476),
            .I(\Commands_frame_decoder.state_1Z0Z_7 ));
    LocalMux I__5740 (
            .O(N__25473),
            .I(\Commands_frame_decoder.state_1Z0Z_7 ));
    InMux I__5739 (
            .O(N__25468),
            .I(N__25465));
    LocalMux I__5738 (
            .O(N__25465),
            .I(N__25462));
    Span4Mux_h I__5737 (
            .O(N__25462),
            .I(N__25458));
    InMux I__5736 (
            .O(N__25461),
            .I(N__25455));
    Span4Mux_v I__5735 (
            .O(N__25458),
            .I(N__25450));
    LocalMux I__5734 (
            .O(N__25455),
            .I(N__25450));
    Span4Mux_v I__5733 (
            .O(N__25450),
            .I(N__25447));
    Odrv4 I__5732 (
            .O(N__25447),
            .I(scaler_4_data_7));
    InMux I__5731 (
            .O(N__25444),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    InMux I__5730 (
            .O(N__25441),
            .I(N__25438));
    LocalMux I__5729 (
            .O(N__25438),
            .I(N__25434));
    InMux I__5728 (
            .O(N__25437),
            .I(N__25431));
    Span4Mux_v I__5727 (
            .O(N__25434),
            .I(N__25426));
    LocalMux I__5726 (
            .O(N__25431),
            .I(N__25426));
    Span4Mux_v I__5725 (
            .O(N__25426),
            .I(N__25423));
    Odrv4 I__5724 (
            .O(N__25423),
            .I(scaler_4_data_8));
    InMux I__5723 (
            .O(N__25420),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    InMux I__5722 (
            .O(N__25417),
            .I(N__25414));
    LocalMux I__5721 (
            .O(N__25414),
            .I(N__25410));
    InMux I__5720 (
            .O(N__25413),
            .I(N__25407));
    Span4Mux_v I__5719 (
            .O(N__25410),
            .I(N__25402));
    LocalMux I__5718 (
            .O(N__25407),
            .I(N__25402));
    Span4Mux_v I__5717 (
            .O(N__25402),
            .I(N__25399));
    Odrv4 I__5716 (
            .O(N__25399),
            .I(scaler_4_data_9));
    InMux I__5715 (
            .O(N__25396),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    InMux I__5714 (
            .O(N__25393),
            .I(N__25390));
    LocalMux I__5713 (
            .O(N__25390),
            .I(N__25386));
    InMux I__5712 (
            .O(N__25389),
            .I(N__25383));
    Span4Mux_v I__5711 (
            .O(N__25386),
            .I(N__25378));
    LocalMux I__5710 (
            .O(N__25383),
            .I(N__25378));
    Span4Mux_v I__5709 (
            .O(N__25378),
            .I(N__25375));
    Odrv4 I__5708 (
            .O(N__25375),
            .I(scaler_4_data_10));
    InMux I__5707 (
            .O(N__25372),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    InMux I__5706 (
            .O(N__25369),
            .I(N__25366));
    LocalMux I__5705 (
            .O(N__25366),
            .I(N__25362));
    InMux I__5704 (
            .O(N__25365),
            .I(N__25359));
    Span4Mux_v I__5703 (
            .O(N__25362),
            .I(N__25354));
    LocalMux I__5702 (
            .O(N__25359),
            .I(N__25354));
    Span4Mux_v I__5701 (
            .O(N__25354),
            .I(N__25351));
    Odrv4 I__5700 (
            .O(N__25351),
            .I(scaler_4_data_11));
    InMux I__5699 (
            .O(N__25348),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    InMux I__5698 (
            .O(N__25345),
            .I(N__25342));
    LocalMux I__5697 (
            .O(N__25342),
            .I(N__25338));
    InMux I__5696 (
            .O(N__25341),
            .I(N__25335));
    Span4Mux_v I__5695 (
            .O(N__25338),
            .I(N__25330));
    LocalMux I__5694 (
            .O(N__25335),
            .I(N__25330));
    Span4Mux_v I__5693 (
            .O(N__25330),
            .I(N__25327));
    Odrv4 I__5692 (
            .O(N__25327),
            .I(scaler_4_data_12));
    InMux I__5691 (
            .O(N__25324),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__5690 (
            .O(N__25321),
            .I(N__25318));
    LocalMux I__5689 (
            .O(N__25318),
            .I(N__25315));
    Span4Mux_v I__5688 (
            .O(N__25315),
            .I(N__25311));
    InMux I__5687 (
            .O(N__25314),
            .I(N__25308));
    Span4Mux_h I__5686 (
            .O(N__25311),
            .I(N__25303));
    LocalMux I__5685 (
            .O(N__25308),
            .I(N__25303));
    Span4Mux_v I__5684 (
            .O(N__25303),
            .I(N__25300));
    Odrv4 I__5683 (
            .O(N__25300),
            .I(scaler_4_data_13));
    InMux I__5682 (
            .O(N__25297),
            .I(bfn_10_16_0_));
    InMux I__5681 (
            .O(N__25294),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__5680 (
            .O(N__25291),
            .I(N__25288));
    LocalMux I__5679 (
            .O(N__25288),
            .I(N__25285));
    Span4Mux_h I__5678 (
            .O(N__25285),
            .I(N__25282));
    Span4Mux_v I__5677 (
            .O(N__25282),
            .I(N__25279));
    Odrv4 I__5676 (
            .O(N__25279),
            .I(scaler_4_data_14));
    InMux I__5675 (
            .O(N__25276),
            .I(N__25272));
    InMux I__5674 (
            .O(N__25275),
            .I(N__25268));
    LocalMux I__5673 (
            .O(N__25272),
            .I(N__25265));
    CascadeMux I__5672 (
            .O(N__25271),
            .I(N__25262));
    LocalMux I__5671 (
            .O(N__25268),
            .I(N__25258));
    Span4Mux_h I__5670 (
            .O(N__25265),
            .I(N__25255));
    InMux I__5669 (
            .O(N__25262),
            .I(N__25250));
    InMux I__5668 (
            .O(N__25261),
            .I(N__25250));
    Odrv4 I__5667 (
            .O(N__25258),
            .I(\scaler_2.un2_source_data_0 ));
    Odrv4 I__5666 (
            .O(N__25255),
            .I(\scaler_2.un2_source_data_0 ));
    LocalMux I__5665 (
            .O(N__25250),
            .I(\scaler_2.un2_source_data_0 ));
    InMux I__5664 (
            .O(N__25243),
            .I(N__25238));
    InMux I__5663 (
            .O(N__25242),
            .I(N__25235));
    CascadeMux I__5662 (
            .O(N__25241),
            .I(N__25231));
    LocalMux I__5661 (
            .O(N__25238),
            .I(N__25228));
    LocalMux I__5660 (
            .O(N__25235),
            .I(N__25225));
    InMux I__5659 (
            .O(N__25234),
            .I(N__25222));
    InMux I__5658 (
            .O(N__25231),
            .I(N__25219));
    Odrv12 I__5657 (
            .O(N__25228),
            .I(frame_decoder_OFF2data_0));
    Odrv4 I__5656 (
            .O(N__25225),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__5655 (
            .O(N__25222),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__5654 (
            .O(N__25219),
            .I(frame_decoder_OFF2data_0));
    InMux I__5653 (
            .O(N__25210),
            .I(N__25205));
    InMux I__5652 (
            .O(N__25209),
            .I(N__25202));
    InMux I__5651 (
            .O(N__25208),
            .I(N__25199));
    LocalMux I__5650 (
            .O(N__25205),
            .I(N__25195));
    LocalMux I__5649 (
            .O(N__25202),
            .I(N__25192));
    LocalMux I__5648 (
            .O(N__25199),
            .I(N__25189));
    InMux I__5647 (
            .O(N__25198),
            .I(N__25186));
    Span4Mux_v I__5646 (
            .O(N__25195),
            .I(N__25183));
    Span12Mux_h I__5645 (
            .O(N__25192),
            .I(N__25180));
    Span4Mux_h I__5644 (
            .O(N__25189),
            .I(N__25177));
    LocalMux I__5643 (
            .O(N__25186),
            .I(N__25174));
    Odrv4 I__5642 (
            .O(N__25183),
            .I(frame_decoder_CH2data_0));
    Odrv12 I__5641 (
            .O(N__25180),
            .I(frame_decoder_CH2data_0));
    Odrv4 I__5640 (
            .O(N__25177),
            .I(frame_decoder_CH2data_0));
    Odrv4 I__5639 (
            .O(N__25174),
            .I(frame_decoder_CH2data_0));
    CascadeMux I__5638 (
            .O(N__25165),
            .I(N__25162));
    InMux I__5637 (
            .O(N__25162),
            .I(N__25159));
    LocalMux I__5636 (
            .O(N__25159),
            .I(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__5635 (
            .O(N__25156),
            .I(N__25150));
    InMux I__5634 (
            .O(N__25155),
            .I(N__25150));
    LocalMux I__5633 (
            .O(N__25150),
            .I(frame_decoder_OFF4data_7));
    CascadeMux I__5632 (
            .O(N__25147),
            .I(N__25144));
    InMux I__5631 (
            .O(N__25144),
            .I(N__25141));
    LocalMux I__5630 (
            .O(N__25141),
            .I(N__25138));
    Span4Mux_h I__5629 (
            .O(N__25138),
            .I(N__25135));
    Odrv4 I__5628 (
            .O(N__25135),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ));
    InMux I__5627 (
            .O(N__25132),
            .I(N__25128));
    InMux I__5626 (
            .O(N__25131),
            .I(N__25125));
    LocalMux I__5625 (
            .O(N__25128),
            .I(N__25122));
    LocalMux I__5624 (
            .O(N__25125),
            .I(N__25119));
    Span12Mux_v I__5623 (
            .O(N__25122),
            .I(N__25116));
    Span4Mux_v I__5622 (
            .O(N__25119),
            .I(N__25113));
    Odrv12 I__5621 (
            .O(N__25116),
            .I(scaler_4_data_6));
    Odrv4 I__5620 (
            .O(N__25113),
            .I(scaler_4_data_6));
    InMux I__5619 (
            .O(N__25108),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    InMux I__5618 (
            .O(N__25105),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__5617 (
            .O(N__25102),
            .I(bfn_9_20_0_));
    InMux I__5616 (
            .O(N__25099),
            .I(N__25095));
    InMux I__5615 (
            .O(N__25098),
            .I(N__25092));
    LocalMux I__5614 (
            .O(N__25095),
            .I(N__25089));
    LocalMux I__5613 (
            .O(N__25092),
            .I(N__25084));
    Span4Mux_h I__5612 (
            .O(N__25089),
            .I(N__25084));
    Span4Mux_v I__5611 (
            .O(N__25084),
            .I(N__25081));
    Odrv4 I__5610 (
            .O(N__25081),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    CEMux I__5609 (
            .O(N__25078),
            .I(N__25073));
    CEMux I__5608 (
            .O(N__25077),
            .I(N__25070));
    CEMux I__5607 (
            .O(N__25076),
            .I(N__25067));
    LocalMux I__5606 (
            .O(N__25073),
            .I(N__25062));
    LocalMux I__5605 (
            .O(N__25070),
            .I(N__25057));
    LocalMux I__5604 (
            .O(N__25067),
            .I(N__25057));
    CEMux I__5603 (
            .O(N__25066),
            .I(N__25054));
    CEMux I__5602 (
            .O(N__25065),
            .I(N__25051));
    Span4Mux_h I__5601 (
            .O(N__25062),
            .I(N__25043));
    Span4Mux_h I__5600 (
            .O(N__25057),
            .I(N__25043));
    LocalMux I__5599 (
            .O(N__25054),
            .I(N__25043));
    LocalMux I__5598 (
            .O(N__25051),
            .I(N__25039));
    CEMux I__5597 (
            .O(N__25050),
            .I(N__25036));
    Sp12to4 I__5596 (
            .O(N__25043),
            .I(N__25033));
    CEMux I__5595 (
            .O(N__25042),
            .I(N__25030));
    Span4Mux_h I__5594 (
            .O(N__25039),
            .I(N__25025));
    LocalMux I__5593 (
            .O(N__25036),
            .I(N__25025));
    Span12Mux_s4_h I__5592 (
            .O(N__25033),
            .I(N__25020));
    LocalMux I__5591 (
            .O(N__25030),
            .I(N__25020));
    Odrv4 I__5590 (
            .O(N__25025),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv12 I__5589 (
            .O(N__25020),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    InMux I__5588 (
            .O(N__25015),
            .I(N__25012));
    LocalMux I__5587 (
            .O(N__25012),
            .I(N__25009));
    Odrv4 I__5586 (
            .O(N__25009),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__5585 (
            .O(N__25006),
            .I(N__25002));
    InMux I__5584 (
            .O(N__25005),
            .I(N__24998));
    LocalMux I__5583 (
            .O(N__25002),
            .I(N__24995));
    CascadeMux I__5582 (
            .O(N__25001),
            .I(N__24992));
    LocalMux I__5581 (
            .O(N__24998),
            .I(N__24987));
    Span4Mux_h I__5580 (
            .O(N__24995),
            .I(N__24987));
    InMux I__5579 (
            .O(N__24992),
            .I(N__24984));
    Span4Mux_h I__5578 (
            .O(N__24987),
            .I(N__24981));
    LocalMux I__5577 (
            .O(N__24984),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    Odrv4 I__5576 (
            .O(N__24981),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__5575 (
            .O(N__24976),
            .I(N__24973));
    LocalMux I__5574 (
            .O(N__24973),
            .I(N__24970));
    Odrv12 I__5573 (
            .O(N__24970),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    CascadeMux I__5572 (
            .O(N__24967),
            .I(N__24956));
    CascadeMux I__5571 (
            .O(N__24966),
            .I(N__24951));
    CascadeMux I__5570 (
            .O(N__24965),
            .I(N__24944));
    CascadeMux I__5569 (
            .O(N__24964),
            .I(N__24941));
    CascadeMux I__5568 (
            .O(N__24963),
            .I(N__24935));
    CascadeMux I__5567 (
            .O(N__24962),
            .I(N__24932));
    CascadeMux I__5566 (
            .O(N__24961),
            .I(N__24929));
    CascadeMux I__5565 (
            .O(N__24960),
            .I(N__24926));
    CascadeMux I__5564 (
            .O(N__24959),
            .I(N__24923));
    InMux I__5563 (
            .O(N__24956),
            .I(N__24920));
    InMux I__5562 (
            .O(N__24955),
            .I(N__24917));
    InMux I__5561 (
            .O(N__24954),
            .I(N__24914));
    InMux I__5560 (
            .O(N__24951),
            .I(N__24904));
    InMux I__5559 (
            .O(N__24950),
            .I(N__24891));
    InMux I__5558 (
            .O(N__24949),
            .I(N__24891));
    InMux I__5557 (
            .O(N__24948),
            .I(N__24891));
    InMux I__5556 (
            .O(N__24947),
            .I(N__24891));
    InMux I__5555 (
            .O(N__24944),
            .I(N__24891));
    InMux I__5554 (
            .O(N__24941),
            .I(N__24891));
    InMux I__5553 (
            .O(N__24940),
            .I(N__24880));
    InMux I__5552 (
            .O(N__24939),
            .I(N__24880));
    InMux I__5551 (
            .O(N__24938),
            .I(N__24880));
    InMux I__5550 (
            .O(N__24935),
            .I(N__24880));
    InMux I__5549 (
            .O(N__24932),
            .I(N__24880));
    InMux I__5548 (
            .O(N__24929),
            .I(N__24877));
    InMux I__5547 (
            .O(N__24926),
            .I(N__24874));
    InMux I__5546 (
            .O(N__24923),
            .I(N__24871));
    LocalMux I__5545 (
            .O(N__24920),
            .I(N__24857));
    LocalMux I__5544 (
            .O(N__24917),
            .I(N__24857));
    LocalMux I__5543 (
            .O(N__24914),
            .I(N__24857));
    InMux I__5542 (
            .O(N__24913),
            .I(N__24854));
    CascadeMux I__5541 (
            .O(N__24912),
            .I(N__24850));
    CascadeMux I__5540 (
            .O(N__24911),
            .I(N__24847));
    CascadeMux I__5539 (
            .O(N__24910),
            .I(N__24844));
    CascadeMux I__5538 (
            .O(N__24909),
            .I(N__24837));
    CascadeMux I__5537 (
            .O(N__24908),
            .I(N__24834));
    InMux I__5536 (
            .O(N__24907),
            .I(N__24831));
    LocalMux I__5535 (
            .O(N__24904),
            .I(N__24828));
    LocalMux I__5534 (
            .O(N__24891),
            .I(N__24823));
    LocalMux I__5533 (
            .O(N__24880),
            .I(N__24823));
    LocalMux I__5532 (
            .O(N__24877),
            .I(N__24820));
    LocalMux I__5531 (
            .O(N__24874),
            .I(N__24815));
    LocalMux I__5530 (
            .O(N__24871),
            .I(N__24815));
    CascadeMux I__5529 (
            .O(N__24870),
            .I(N__24812));
    CascadeMux I__5528 (
            .O(N__24869),
            .I(N__24809));
    CascadeMux I__5527 (
            .O(N__24868),
            .I(N__24806));
    InMux I__5526 (
            .O(N__24867),
            .I(N__24799));
    InMux I__5525 (
            .O(N__24866),
            .I(N__24799));
    InMux I__5524 (
            .O(N__24865),
            .I(N__24799));
    InMux I__5523 (
            .O(N__24864),
            .I(N__24794));
    Span4Mux_v I__5522 (
            .O(N__24857),
            .I(N__24791));
    LocalMux I__5521 (
            .O(N__24854),
            .I(N__24788));
    InMux I__5520 (
            .O(N__24853),
            .I(N__24779));
    InMux I__5519 (
            .O(N__24850),
            .I(N__24779));
    InMux I__5518 (
            .O(N__24847),
            .I(N__24779));
    InMux I__5517 (
            .O(N__24844),
            .I(N__24779));
    InMux I__5516 (
            .O(N__24843),
            .I(N__24770));
    InMux I__5515 (
            .O(N__24842),
            .I(N__24770));
    InMux I__5514 (
            .O(N__24841),
            .I(N__24770));
    InMux I__5513 (
            .O(N__24840),
            .I(N__24770));
    InMux I__5512 (
            .O(N__24837),
            .I(N__24767));
    InMux I__5511 (
            .O(N__24834),
            .I(N__24764));
    LocalMux I__5510 (
            .O(N__24831),
            .I(N__24761));
    Span4Mux_v I__5509 (
            .O(N__24828),
            .I(N__24754));
    Span4Mux_v I__5508 (
            .O(N__24823),
            .I(N__24754));
    Span4Mux_h I__5507 (
            .O(N__24820),
            .I(N__24754));
    Span4Mux_v I__5506 (
            .O(N__24815),
            .I(N__24751));
    InMux I__5505 (
            .O(N__24812),
            .I(N__24744));
    InMux I__5504 (
            .O(N__24809),
            .I(N__24744));
    InMux I__5503 (
            .O(N__24806),
            .I(N__24744));
    LocalMux I__5502 (
            .O(N__24799),
            .I(N__24741));
    CascadeMux I__5501 (
            .O(N__24798),
            .I(N__24738));
    InMux I__5500 (
            .O(N__24797),
            .I(N__24735));
    LocalMux I__5499 (
            .O(N__24794),
            .I(N__24732));
    Span4Mux_h I__5498 (
            .O(N__24791),
            .I(N__24727));
    Span4Mux_h I__5497 (
            .O(N__24788),
            .I(N__24727));
    LocalMux I__5496 (
            .O(N__24779),
            .I(N__24714));
    LocalMux I__5495 (
            .O(N__24770),
            .I(N__24714));
    LocalMux I__5494 (
            .O(N__24767),
            .I(N__24714));
    LocalMux I__5493 (
            .O(N__24764),
            .I(N__24714));
    Span4Mux_v I__5492 (
            .O(N__24761),
            .I(N__24714));
    Span4Mux_h I__5491 (
            .O(N__24754),
            .I(N__24714));
    Span4Mux_h I__5490 (
            .O(N__24751),
            .I(N__24707));
    LocalMux I__5489 (
            .O(N__24744),
            .I(N__24707));
    Span4Mux_h I__5488 (
            .O(N__24741),
            .I(N__24707));
    InMux I__5487 (
            .O(N__24738),
            .I(N__24704));
    LocalMux I__5486 (
            .O(N__24735),
            .I(N__24701));
    Span4Mux_v I__5485 (
            .O(N__24732),
            .I(N__24696));
    Span4Mux_v I__5484 (
            .O(N__24727),
            .I(N__24696));
    Span4Mux_v I__5483 (
            .O(N__24714),
            .I(N__24693));
    Span4Mux_v I__5482 (
            .O(N__24707),
            .I(N__24690));
    LocalMux I__5481 (
            .O(N__24704),
            .I(N__24685));
    Span4Mux_v I__5480 (
            .O(N__24701),
            .I(N__24685));
    Odrv4 I__5479 (
            .O(N__24696),
            .I(pid_altitude_dv));
    Odrv4 I__5478 (
            .O(N__24693),
            .I(pid_altitude_dv));
    Odrv4 I__5477 (
            .O(N__24690),
            .I(pid_altitude_dv));
    Odrv4 I__5476 (
            .O(N__24685),
            .I(pid_altitude_dv));
    InMux I__5475 (
            .O(N__24676),
            .I(N__24671));
    InMux I__5474 (
            .O(N__24675),
            .I(N__24668));
    InMux I__5473 (
            .O(N__24674),
            .I(N__24665));
    LocalMux I__5472 (
            .O(N__24671),
            .I(N__24660));
    LocalMux I__5471 (
            .O(N__24668),
            .I(N__24660));
    LocalMux I__5470 (
            .O(N__24665),
            .I(N__24655));
    Span4Mux_h I__5469 (
            .O(N__24660),
            .I(N__24655));
    Odrv4 I__5468 (
            .O(N__24655),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__5467 (
            .O(N__24652),
            .I(N__24648));
    InMux I__5466 (
            .O(N__24651),
            .I(N__24645));
    LocalMux I__5465 (
            .O(N__24648),
            .I(N__24642));
    LocalMux I__5464 (
            .O(N__24645),
            .I(N__24639));
    Odrv4 I__5463 (
            .O(N__24642),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    Odrv12 I__5462 (
            .O(N__24639),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__5461 (
            .O(N__24634),
            .I(N__24628));
    InMux I__5460 (
            .O(N__24633),
            .I(N__24628));
    LocalMux I__5459 (
            .O(N__24628),
            .I(frame_decoder_CH4data_7));
    CEMux I__5458 (
            .O(N__24625),
            .I(N__24621));
    CEMux I__5457 (
            .O(N__24624),
            .I(N__24618));
    LocalMux I__5456 (
            .O(N__24621),
            .I(N__24614));
    LocalMux I__5455 (
            .O(N__24618),
            .I(N__24611));
    CEMux I__5454 (
            .O(N__24617),
            .I(N__24608));
    Span4Mux_h I__5453 (
            .O(N__24614),
            .I(N__24605));
    Span4Mux_v I__5452 (
            .O(N__24611),
            .I(N__24600));
    LocalMux I__5451 (
            .O(N__24608),
            .I(N__24600));
    Span4Mux_h I__5450 (
            .O(N__24605),
            .I(N__24597));
    Sp12to4 I__5449 (
            .O(N__24600),
            .I(N__24594));
    Odrv4 I__5448 (
            .O(N__24597),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    Odrv12 I__5447 (
            .O(N__24594),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    InMux I__5446 (
            .O(N__24589),
            .I(N__24586));
    LocalMux I__5445 (
            .O(N__24586),
            .I(N__24583));
    Span4Mux_v I__5444 (
            .O(N__24583),
            .I(N__24580));
    Span4Mux_h I__5443 (
            .O(N__24580),
            .I(N__24577));
    Span4Mux_h I__5442 (
            .O(N__24577),
            .I(N__24574));
    Odrv4 I__5441 (
            .O(N__24574),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__5440 (
            .O(N__24571),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__5439 (
            .O(N__24568),
            .I(N__24565));
    LocalMux I__5438 (
            .O(N__24565),
            .I(N__24562));
    Span4Mux_v I__5437 (
            .O(N__24562),
            .I(N__24559));
    Odrv4 I__5436 (
            .O(N__24559),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__5435 (
            .O(N__24556),
            .I(\ppm_encoder_1.un1_elevator_cry_7 ));
    InMux I__5434 (
            .O(N__24553),
            .I(N__24550));
    LocalMux I__5433 (
            .O(N__24550),
            .I(N__24547));
    Span4Mux_v I__5432 (
            .O(N__24547),
            .I(N__24544));
    Span4Mux_h I__5431 (
            .O(N__24544),
            .I(N__24541));
    Odrv4 I__5430 (
            .O(N__24541),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__5429 (
            .O(N__24538),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__5428 (
            .O(N__24535),
            .I(N__24532));
    LocalMux I__5427 (
            .O(N__24532),
            .I(N__24529));
    Odrv4 I__5426 (
            .O(N__24529),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__5425 (
            .O(N__24526),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__5424 (
            .O(N__24523),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__5423 (
            .O(N__24520),
            .I(N__24517));
    LocalMux I__5422 (
            .O(N__24517),
            .I(N__24514));
    Odrv4 I__5421 (
            .O(N__24514),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__5420 (
            .O(N__24511),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__5419 (
            .O(N__24508),
            .I(N__24505));
    LocalMux I__5418 (
            .O(N__24505),
            .I(N__24502));
    Span4Mux_h I__5417 (
            .O(N__24502),
            .I(N__24499));
    Span4Mux_v I__5416 (
            .O(N__24499),
            .I(N__24495));
    CascadeMux I__5415 (
            .O(N__24498),
            .I(N__24492));
    Span4Mux_v I__5414 (
            .O(N__24495),
            .I(N__24489));
    InMux I__5413 (
            .O(N__24492),
            .I(N__24486));
    Odrv4 I__5412 (
            .O(N__24489),
            .I(scaler_3_data_4));
    LocalMux I__5411 (
            .O(N__24486),
            .I(scaler_3_data_4));
    InMux I__5410 (
            .O(N__24481),
            .I(N__24478));
    LocalMux I__5409 (
            .O(N__24478),
            .I(N__24475));
    Span4Mux_h I__5408 (
            .O(N__24475),
            .I(N__24472));
    Span4Mux_h I__5407 (
            .O(N__24472),
            .I(N__24469));
    Span4Mux_v I__5406 (
            .O(N__24469),
            .I(N__24465));
    CascadeMux I__5405 (
            .O(N__24468),
            .I(N__24462));
    Span4Mux_v I__5404 (
            .O(N__24465),
            .I(N__24459));
    InMux I__5403 (
            .O(N__24462),
            .I(N__24456));
    Odrv4 I__5402 (
            .O(N__24459),
            .I(scaler_4_data_4));
    LocalMux I__5401 (
            .O(N__24456),
            .I(scaler_4_data_4));
    CascadeMux I__5400 (
            .O(N__24451),
            .I(\Commands_frame_decoder.N_282_0_cascade_ ));
    InMux I__5399 (
            .O(N__24448),
            .I(N__24444));
    InMux I__5398 (
            .O(N__24447),
            .I(N__24441));
    LocalMux I__5397 (
            .O(N__24444),
            .I(N__24436));
    LocalMux I__5396 (
            .O(N__24441),
            .I(N__24436));
    Odrv4 I__5395 (
            .O(N__24436),
            .I(\Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1 ));
    InMux I__5394 (
            .O(N__24433),
            .I(N__24430));
    LocalMux I__5393 (
            .O(N__24430),
            .I(N__24427));
    Span4Mux_h I__5392 (
            .O(N__24427),
            .I(N__24424));
    Span4Mux_h I__5391 (
            .O(N__24424),
            .I(N__24421));
    Odrv4 I__5390 (
            .O(N__24421),
            .I(\Commands_frame_decoder.source_CH1data8lto7Z0Z_1 ));
    CascadeMux I__5389 (
            .O(N__24418),
            .I(\Commands_frame_decoder.N_319_cascade_ ));
    InMux I__5388 (
            .O(N__24415),
            .I(N__24412));
    LocalMux I__5387 (
            .O(N__24412),
            .I(\Commands_frame_decoder.N_318 ));
    InMux I__5386 (
            .O(N__24409),
            .I(N__24406));
    LocalMux I__5385 (
            .O(N__24406),
            .I(\Commands_frame_decoder.N_282_0 ));
    InMux I__5384 (
            .O(N__24403),
            .I(N__24400));
    LocalMux I__5383 (
            .O(N__24400),
            .I(\Commands_frame_decoder.state_1_RNO_1Z0Z_0 ));
    CascadeMux I__5382 (
            .O(N__24397),
            .I(\Commands_frame_decoder.state_1_ns_i_0_0_cascade_ ));
    CascadeMux I__5381 (
            .O(N__24394),
            .I(N__24390));
    InMux I__5380 (
            .O(N__24393),
            .I(N__24385));
    InMux I__5379 (
            .O(N__24390),
            .I(N__24385));
    LocalMux I__5378 (
            .O(N__24385),
            .I(\Commands_frame_decoder.state_1Z0Z_0 ));
    InMux I__5377 (
            .O(N__24382),
            .I(N__24376));
    InMux I__5376 (
            .O(N__24381),
            .I(N__24376));
    LocalMux I__5375 (
            .O(N__24376),
            .I(N__24373));
    Span4Mux_h I__5374 (
            .O(N__24373),
            .I(N__24370));
    Odrv4 I__5373 (
            .O(N__24370),
            .I(\Commands_frame_decoder.N_323 ));
    InMux I__5372 (
            .O(N__24367),
            .I(N__24364));
    LocalMux I__5371 (
            .O(N__24364),
            .I(\Commands_frame_decoder.state_1_ns_0_a4_0_2_1 ));
    InMux I__5370 (
            .O(N__24361),
            .I(N__24358));
    LocalMux I__5369 (
            .O(N__24358),
            .I(N__24355));
    Span4Mux_h I__5368 (
            .O(N__24355),
            .I(N__24350));
    CascadeMux I__5367 (
            .O(N__24354),
            .I(N__24347));
    CascadeMux I__5366 (
            .O(N__24353),
            .I(N__24344));
    Span4Mux_h I__5365 (
            .O(N__24350),
            .I(N__24340));
    InMux I__5364 (
            .O(N__24347),
            .I(N__24333));
    InMux I__5363 (
            .O(N__24344),
            .I(N__24333));
    InMux I__5362 (
            .O(N__24343),
            .I(N__24333));
    Odrv4 I__5361 (
            .O(N__24340),
            .I(\Commands_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__5360 (
            .O(N__24333),
            .I(\Commands_frame_decoder.state_1Z0Z_1 ));
    InMux I__5359 (
            .O(N__24328),
            .I(N__24324));
    InMux I__5358 (
            .O(N__24327),
            .I(N__24321));
    LocalMux I__5357 (
            .O(N__24324),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    LocalMux I__5356 (
            .O(N__24321),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    CascadeMux I__5355 (
            .O(N__24316),
            .I(N__24313));
    InMux I__5354 (
            .O(N__24313),
            .I(N__24310));
    LocalMux I__5353 (
            .O(N__24310),
            .I(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ));
    InMux I__5352 (
            .O(N__24307),
            .I(N__24303));
    InMux I__5351 (
            .O(N__24306),
            .I(N__24300));
    LocalMux I__5350 (
            .O(N__24303),
            .I(N__24297));
    LocalMux I__5349 (
            .O(N__24300),
            .I(N__24294));
    Span12Mux_s9_h I__5348 (
            .O(N__24297),
            .I(N__24291));
    Span4Mux_v I__5347 (
            .O(N__24294),
            .I(N__24288));
    Odrv12 I__5346 (
            .O(N__24291),
            .I(scaler_2_data_13));
    Odrv4 I__5345 (
            .O(N__24288),
            .I(scaler_2_data_13));
    InMux I__5344 (
            .O(N__24283),
            .I(bfn_9_14_0_));
    InMux I__5343 (
            .O(N__24280),
            .I(\scaler_2.un2_source_data_0_cry_9 ));
    InMux I__5342 (
            .O(N__24277),
            .I(N__24274));
    LocalMux I__5341 (
            .O(N__24274),
            .I(N__24271));
    Span4Mux_v I__5340 (
            .O(N__24271),
            .I(N__24268));
    Odrv4 I__5339 (
            .O(N__24268),
            .I(scaler_2_data_14));
    InMux I__5338 (
            .O(N__24265),
            .I(N__24262));
    LocalMux I__5337 (
            .O(N__24262),
            .I(N__24259));
    Sp12to4 I__5336 (
            .O(N__24259),
            .I(N__24256));
    Span12Mux_v I__5335 (
            .O(N__24256),
            .I(N__24253));
    Odrv12 I__5334 (
            .O(N__24253),
            .I(scaler_2_data_5));
    InMux I__5333 (
            .O(N__24250),
            .I(N__24247));
    LocalMux I__5332 (
            .O(N__24247),
            .I(N__24244));
    Span4Mux_h I__5331 (
            .O(N__24244),
            .I(N__24241));
    Span4Mux_v I__5330 (
            .O(N__24241),
            .I(N__24238));
    Span4Mux_v I__5329 (
            .O(N__24238),
            .I(N__24235));
    Odrv4 I__5328 (
            .O(N__24235),
            .I(scaler_3_data_5));
    InMux I__5327 (
            .O(N__24232),
            .I(N__24229));
    LocalMux I__5326 (
            .O(N__24229),
            .I(N__24226));
    Span4Mux_v I__5325 (
            .O(N__24226),
            .I(N__24223));
    Span4Mux_v I__5324 (
            .O(N__24223),
            .I(N__24220));
    Span4Mux_h I__5323 (
            .O(N__24220),
            .I(N__24217));
    Odrv4 I__5322 (
            .O(N__24217),
            .I(scaler_4_data_5));
    InMux I__5321 (
            .O(N__24214),
            .I(N__24211));
    LocalMux I__5320 (
            .O(N__24211),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__5319 (
            .O(N__24208),
            .I(N__24205));
    LocalMux I__5318 (
            .O(N__24205),
            .I(N__24202));
    Span4Mux_v I__5317 (
            .O(N__24202),
            .I(N__24199));
    Span4Mux_v I__5316 (
            .O(N__24199),
            .I(N__24195));
    CascadeMux I__5315 (
            .O(N__24198),
            .I(N__24192));
    Span4Mux_h I__5314 (
            .O(N__24195),
            .I(N__24189));
    InMux I__5313 (
            .O(N__24192),
            .I(N__24186));
    Odrv4 I__5312 (
            .O(N__24189),
            .I(scaler_2_data_4));
    LocalMux I__5311 (
            .O(N__24186),
            .I(scaler_2_data_4));
    CascadeMux I__5310 (
            .O(N__24181),
            .I(N__24178));
    InMux I__5309 (
            .O(N__24178),
            .I(N__24175));
    LocalMux I__5308 (
            .O(N__24175),
            .I(frame_decoder_OFF2data_2));
    InMux I__5307 (
            .O(N__24172),
            .I(N__24169));
    LocalMux I__5306 (
            .O(N__24169),
            .I(N__24166));
    Span4Mux_v I__5305 (
            .O(N__24166),
            .I(N__24163));
    Span4Mux_h I__5304 (
            .O(N__24163),
            .I(N__24159));
    InMux I__5303 (
            .O(N__24162),
            .I(N__24156));
    Span4Mux_h I__5302 (
            .O(N__24159),
            .I(N__24151));
    LocalMux I__5301 (
            .O(N__24156),
            .I(N__24151));
    Sp12to4 I__5300 (
            .O(N__24151),
            .I(N__24148));
    Odrv12 I__5299 (
            .O(N__24148),
            .I(scaler_2_data_6));
    InMux I__5298 (
            .O(N__24145),
            .I(\scaler_2.un2_source_data_0_cry_1 ));
    CascadeMux I__5297 (
            .O(N__24142),
            .I(N__24139));
    InMux I__5296 (
            .O(N__24139),
            .I(N__24133));
    InMux I__5295 (
            .O(N__24138),
            .I(N__24133));
    LocalMux I__5294 (
            .O(N__24133),
            .I(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ));
    InMux I__5293 (
            .O(N__24130),
            .I(N__24126));
    InMux I__5292 (
            .O(N__24129),
            .I(N__24123));
    LocalMux I__5291 (
            .O(N__24126),
            .I(N__24120));
    LocalMux I__5290 (
            .O(N__24123),
            .I(N__24117));
    Span12Mux_s9_h I__5289 (
            .O(N__24120),
            .I(N__24114));
    Span4Mux_v I__5288 (
            .O(N__24117),
            .I(N__24111));
    Odrv12 I__5287 (
            .O(N__24114),
            .I(scaler_2_data_7));
    Odrv4 I__5286 (
            .O(N__24111),
            .I(scaler_2_data_7));
    InMux I__5285 (
            .O(N__24106),
            .I(\scaler_2.un2_source_data_0_cry_2 ));
    CascadeMux I__5284 (
            .O(N__24103),
            .I(N__24100));
    InMux I__5283 (
            .O(N__24100),
            .I(N__24094));
    InMux I__5282 (
            .O(N__24099),
            .I(N__24094));
    LocalMux I__5281 (
            .O(N__24094),
            .I(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ));
    InMux I__5280 (
            .O(N__24091),
            .I(N__24088));
    LocalMux I__5279 (
            .O(N__24088),
            .I(N__24085));
    Span4Mux_v I__5278 (
            .O(N__24085),
            .I(N__24081));
    InMux I__5277 (
            .O(N__24084),
            .I(N__24078));
    Span4Mux_h I__5276 (
            .O(N__24081),
            .I(N__24073));
    LocalMux I__5275 (
            .O(N__24078),
            .I(N__24073));
    Span4Mux_v I__5274 (
            .O(N__24073),
            .I(N__24070));
    Odrv4 I__5273 (
            .O(N__24070),
            .I(scaler_2_data_8));
    InMux I__5272 (
            .O(N__24067),
            .I(\scaler_2.un2_source_data_0_cry_3 ));
    CascadeMux I__5271 (
            .O(N__24064),
            .I(N__24061));
    InMux I__5270 (
            .O(N__24061),
            .I(N__24055));
    InMux I__5269 (
            .O(N__24060),
            .I(N__24055));
    LocalMux I__5268 (
            .O(N__24055),
            .I(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ));
    InMux I__5267 (
            .O(N__24052),
            .I(N__24049));
    LocalMux I__5266 (
            .O(N__24049),
            .I(N__24045));
    InMux I__5265 (
            .O(N__24048),
            .I(N__24042));
    Span4Mux_v I__5264 (
            .O(N__24045),
            .I(N__24039));
    LocalMux I__5263 (
            .O(N__24042),
            .I(N__24036));
    Span4Mux_v I__5262 (
            .O(N__24039),
            .I(N__24033));
    Span4Mux_v I__5261 (
            .O(N__24036),
            .I(N__24030));
    Odrv4 I__5260 (
            .O(N__24033),
            .I(scaler_2_data_9));
    Odrv4 I__5259 (
            .O(N__24030),
            .I(scaler_2_data_9));
    InMux I__5258 (
            .O(N__24025),
            .I(\scaler_2.un2_source_data_0_cry_4 ));
    CascadeMux I__5257 (
            .O(N__24022),
            .I(N__24019));
    InMux I__5256 (
            .O(N__24019),
            .I(N__24013));
    InMux I__5255 (
            .O(N__24018),
            .I(N__24013));
    LocalMux I__5254 (
            .O(N__24013),
            .I(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ));
    InMux I__5253 (
            .O(N__24010),
            .I(N__24007));
    LocalMux I__5252 (
            .O(N__24007),
            .I(N__24004));
    Span4Mux_h I__5251 (
            .O(N__24004),
            .I(N__24000));
    InMux I__5250 (
            .O(N__24003),
            .I(N__23997));
    Span4Mux_v I__5249 (
            .O(N__24000),
            .I(N__23994));
    LocalMux I__5248 (
            .O(N__23997),
            .I(N__23991));
    Span4Mux_v I__5247 (
            .O(N__23994),
            .I(N__23988));
    Span4Mux_v I__5246 (
            .O(N__23991),
            .I(N__23985));
    Odrv4 I__5245 (
            .O(N__23988),
            .I(scaler_2_data_10));
    Odrv4 I__5244 (
            .O(N__23985),
            .I(scaler_2_data_10));
    InMux I__5243 (
            .O(N__23980),
            .I(\scaler_2.un2_source_data_0_cry_5 ));
    CascadeMux I__5242 (
            .O(N__23977),
            .I(N__23974));
    InMux I__5241 (
            .O(N__23974),
            .I(N__23968));
    InMux I__5240 (
            .O(N__23973),
            .I(N__23968));
    LocalMux I__5239 (
            .O(N__23968),
            .I(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ));
    InMux I__5238 (
            .O(N__23965),
            .I(N__23962));
    LocalMux I__5237 (
            .O(N__23962),
            .I(N__23959));
    Span4Mux_v I__5236 (
            .O(N__23959),
            .I(N__23955));
    InMux I__5235 (
            .O(N__23958),
            .I(N__23952));
    Sp12to4 I__5234 (
            .O(N__23955),
            .I(N__23947));
    LocalMux I__5233 (
            .O(N__23952),
            .I(N__23947));
    Span12Mux_s9_h I__5232 (
            .O(N__23947),
            .I(N__23944));
    Odrv12 I__5231 (
            .O(N__23944),
            .I(scaler_2_data_11));
    InMux I__5230 (
            .O(N__23941),
            .I(\scaler_2.un2_source_data_0_cry_6 ));
    CascadeMux I__5229 (
            .O(N__23938),
            .I(N__23935));
    InMux I__5228 (
            .O(N__23935),
            .I(N__23929));
    InMux I__5227 (
            .O(N__23934),
            .I(N__23929));
    LocalMux I__5226 (
            .O(N__23929),
            .I(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ));
    InMux I__5225 (
            .O(N__23926),
            .I(N__23923));
    LocalMux I__5224 (
            .O(N__23923),
            .I(N__23920));
    Span4Mux_v I__5223 (
            .O(N__23920),
            .I(N__23916));
    InMux I__5222 (
            .O(N__23919),
            .I(N__23913));
    Sp12to4 I__5221 (
            .O(N__23916),
            .I(N__23910));
    LocalMux I__5220 (
            .O(N__23913),
            .I(N__23907));
    Span12Mux_s9_h I__5219 (
            .O(N__23910),
            .I(N__23904));
    Span4Mux_v I__5218 (
            .O(N__23907),
            .I(N__23901));
    Odrv12 I__5217 (
            .O(N__23904),
            .I(scaler_2_data_12));
    Odrv4 I__5216 (
            .O(N__23901),
            .I(scaler_2_data_12));
    InMux I__5215 (
            .O(N__23896),
            .I(\scaler_2.un2_source_data_0_cry_7 ));
    InMux I__5214 (
            .O(N__23893),
            .I(N__23890));
    LocalMux I__5213 (
            .O(N__23890),
            .I(N__23887));
    Span4Mux_s3_v I__5212 (
            .O(N__23887),
            .I(N__23882));
    InMux I__5211 (
            .O(N__23886),
            .I(N__23877));
    InMux I__5210 (
            .O(N__23885),
            .I(N__23877));
    Odrv4 I__5209 (
            .O(N__23882),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__5208 (
            .O(N__23877),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    CascadeMux I__5207 (
            .O(N__23872),
            .I(N__23867));
    CascadeMux I__5206 (
            .O(N__23871),
            .I(N__23864));
    InMux I__5205 (
            .O(N__23870),
            .I(N__23857));
    InMux I__5204 (
            .O(N__23867),
            .I(N__23857));
    InMux I__5203 (
            .O(N__23864),
            .I(N__23857));
    LocalMux I__5202 (
            .O(N__23857),
            .I(N__23854));
    Span4Mux_s3_v I__5201 (
            .O(N__23854),
            .I(N__23851));
    Span4Mux_v I__5200 (
            .O(N__23851),
            .I(N__23846));
    InMux I__5199 (
            .O(N__23850),
            .I(N__23843));
    InMux I__5198 (
            .O(N__23849),
            .I(N__23840));
    Sp12to4 I__5197 (
            .O(N__23846),
            .I(N__23835));
    LocalMux I__5196 (
            .O(N__23843),
            .I(N__23835));
    LocalMux I__5195 (
            .O(N__23840),
            .I(N__23832));
    Odrv12 I__5194 (
            .O(N__23835),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_158_d ));
    Odrv12 I__5193 (
            .O(N__23832),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_158_d ));
    InMux I__5192 (
            .O(N__23827),
            .I(N__23814));
    InMux I__5191 (
            .O(N__23826),
            .I(N__23814));
    InMux I__5190 (
            .O(N__23825),
            .I(N__23814));
    CascadeMux I__5189 (
            .O(N__23824),
            .I(N__23804));
    CascadeMux I__5188 (
            .O(N__23823),
            .I(N__23801));
    InMux I__5187 (
            .O(N__23822),
            .I(N__23789));
    InMux I__5186 (
            .O(N__23821),
            .I(N__23789));
    LocalMux I__5185 (
            .O(N__23814),
            .I(N__23781));
    CascadeMux I__5184 (
            .O(N__23813),
            .I(N__23777));
    CascadeMux I__5183 (
            .O(N__23812),
            .I(N__23774));
    CascadeMux I__5182 (
            .O(N__23811),
            .I(N__23768));
    CascadeMux I__5181 (
            .O(N__23810),
            .I(N__23764));
    CascadeMux I__5180 (
            .O(N__23809),
            .I(N__23757));
    InMux I__5179 (
            .O(N__23808),
            .I(N__23750));
    CascadeMux I__5178 (
            .O(N__23807),
            .I(N__23745));
    InMux I__5177 (
            .O(N__23804),
            .I(N__23737));
    InMux I__5176 (
            .O(N__23801),
            .I(N__23737));
    InMux I__5175 (
            .O(N__23800),
            .I(N__23737));
    CascadeMux I__5174 (
            .O(N__23799),
            .I(N__23734));
    CascadeMux I__5173 (
            .O(N__23798),
            .I(N__23728));
    InMux I__5172 (
            .O(N__23797),
            .I(N__23725));
    InMux I__5171 (
            .O(N__23796),
            .I(N__23717));
    InMux I__5170 (
            .O(N__23795),
            .I(N__23717));
    InMux I__5169 (
            .O(N__23794),
            .I(N__23717));
    LocalMux I__5168 (
            .O(N__23789),
            .I(N__23714));
    InMux I__5167 (
            .O(N__23788),
            .I(N__23703));
    InMux I__5166 (
            .O(N__23787),
            .I(N__23703));
    InMux I__5165 (
            .O(N__23786),
            .I(N__23703));
    InMux I__5164 (
            .O(N__23785),
            .I(N__23703));
    InMux I__5163 (
            .O(N__23784),
            .I(N__23703));
    Span4Mux_h I__5162 (
            .O(N__23781),
            .I(N__23699));
    InMux I__5161 (
            .O(N__23780),
            .I(N__23696));
    InMux I__5160 (
            .O(N__23777),
            .I(N__23687));
    InMux I__5159 (
            .O(N__23774),
            .I(N__23687));
    InMux I__5158 (
            .O(N__23773),
            .I(N__23687));
    InMux I__5157 (
            .O(N__23772),
            .I(N__23687));
    InMux I__5156 (
            .O(N__23771),
            .I(N__23676));
    InMux I__5155 (
            .O(N__23768),
            .I(N__23676));
    InMux I__5154 (
            .O(N__23767),
            .I(N__23676));
    InMux I__5153 (
            .O(N__23764),
            .I(N__23676));
    InMux I__5152 (
            .O(N__23763),
            .I(N__23676));
    InMux I__5151 (
            .O(N__23762),
            .I(N__23669));
    InMux I__5150 (
            .O(N__23761),
            .I(N__23669));
    InMux I__5149 (
            .O(N__23760),
            .I(N__23669));
    InMux I__5148 (
            .O(N__23757),
            .I(N__23658));
    InMux I__5147 (
            .O(N__23756),
            .I(N__23658));
    InMux I__5146 (
            .O(N__23755),
            .I(N__23658));
    InMux I__5145 (
            .O(N__23754),
            .I(N__23658));
    InMux I__5144 (
            .O(N__23753),
            .I(N__23658));
    LocalMux I__5143 (
            .O(N__23750),
            .I(N__23647));
    InMux I__5142 (
            .O(N__23749),
            .I(N__23638));
    InMux I__5141 (
            .O(N__23748),
            .I(N__23638));
    InMux I__5140 (
            .O(N__23745),
            .I(N__23638));
    InMux I__5139 (
            .O(N__23744),
            .I(N__23638));
    LocalMux I__5138 (
            .O(N__23737),
            .I(N__23635));
    InMux I__5137 (
            .O(N__23734),
            .I(N__23630));
    InMux I__5136 (
            .O(N__23733),
            .I(N__23630));
    InMux I__5135 (
            .O(N__23732),
            .I(N__23624));
    InMux I__5134 (
            .O(N__23731),
            .I(N__23624));
    InMux I__5133 (
            .O(N__23728),
            .I(N__23621));
    LocalMux I__5132 (
            .O(N__23725),
            .I(N__23618));
    CascadeMux I__5131 (
            .O(N__23724),
            .I(N__23614));
    LocalMux I__5130 (
            .O(N__23717),
            .I(N__23605));
    Span4Mux_h I__5129 (
            .O(N__23714),
            .I(N__23605));
    LocalMux I__5128 (
            .O(N__23703),
            .I(N__23605));
    CascadeMux I__5127 (
            .O(N__23702),
            .I(N__23602));
    Span4Mux_h I__5126 (
            .O(N__23699),
            .I(N__23588));
    LocalMux I__5125 (
            .O(N__23696),
            .I(N__23588));
    LocalMux I__5124 (
            .O(N__23687),
            .I(N__23588));
    LocalMux I__5123 (
            .O(N__23676),
            .I(N__23588));
    LocalMux I__5122 (
            .O(N__23669),
            .I(N__23588));
    LocalMux I__5121 (
            .O(N__23658),
            .I(N__23588));
    InMux I__5120 (
            .O(N__23657),
            .I(N__23575));
    InMux I__5119 (
            .O(N__23656),
            .I(N__23575));
    InMux I__5118 (
            .O(N__23655),
            .I(N__23575));
    InMux I__5117 (
            .O(N__23654),
            .I(N__23575));
    InMux I__5116 (
            .O(N__23653),
            .I(N__23575));
    InMux I__5115 (
            .O(N__23652),
            .I(N__23575));
    InMux I__5114 (
            .O(N__23651),
            .I(N__23570));
    InMux I__5113 (
            .O(N__23650),
            .I(N__23570));
    Span4Mux_v I__5112 (
            .O(N__23647),
            .I(N__23561));
    LocalMux I__5111 (
            .O(N__23638),
            .I(N__23561));
    Span4Mux_v I__5110 (
            .O(N__23635),
            .I(N__23561));
    LocalMux I__5109 (
            .O(N__23630),
            .I(N__23561));
    CascadeMux I__5108 (
            .O(N__23629),
            .I(N__23553));
    LocalMux I__5107 (
            .O(N__23624),
            .I(N__23549));
    LocalMux I__5106 (
            .O(N__23621),
            .I(N__23544));
    Span12Mux_h I__5105 (
            .O(N__23618),
            .I(N__23544));
    InMux I__5104 (
            .O(N__23617),
            .I(N__23535));
    InMux I__5103 (
            .O(N__23614),
            .I(N__23535));
    InMux I__5102 (
            .O(N__23613),
            .I(N__23535));
    InMux I__5101 (
            .O(N__23612),
            .I(N__23535));
    Span4Mux_h I__5100 (
            .O(N__23605),
            .I(N__23532));
    InMux I__5099 (
            .O(N__23602),
            .I(N__23527));
    InMux I__5098 (
            .O(N__23601),
            .I(N__23527));
    Span4Mux_v I__5097 (
            .O(N__23588),
            .I(N__23518));
    LocalMux I__5096 (
            .O(N__23575),
            .I(N__23518));
    LocalMux I__5095 (
            .O(N__23570),
            .I(N__23518));
    Span4Mux_h I__5094 (
            .O(N__23561),
            .I(N__23518));
    InMux I__5093 (
            .O(N__23560),
            .I(N__23509));
    InMux I__5092 (
            .O(N__23559),
            .I(N__23509));
    InMux I__5091 (
            .O(N__23558),
            .I(N__23509));
    InMux I__5090 (
            .O(N__23557),
            .I(N__23509));
    InMux I__5089 (
            .O(N__23556),
            .I(N__23502));
    InMux I__5088 (
            .O(N__23553),
            .I(N__23502));
    InMux I__5087 (
            .O(N__23552),
            .I(N__23502));
    Odrv4 I__5086 (
            .O(N__23549),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    Odrv12 I__5085 (
            .O(N__23544),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    LocalMux I__5084 (
            .O(N__23535),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    Odrv4 I__5083 (
            .O(N__23532),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    LocalMux I__5082 (
            .O(N__23527),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    Odrv4 I__5081 (
            .O(N__23518),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    LocalMux I__5080 (
            .O(N__23509),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    LocalMux I__5079 (
            .O(N__23502),
            .I(\ppm_encoder_1.PPM_STATE_58_d ));
    CascadeMux I__5078 (
            .O(N__23485),
            .I(N__23481));
    InMux I__5077 (
            .O(N__23484),
            .I(N__23478));
    InMux I__5076 (
            .O(N__23481),
            .I(N__23475));
    LocalMux I__5075 (
            .O(N__23478),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    LocalMux I__5074 (
            .O(N__23475),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__5073 (
            .O(N__23470),
            .I(N__23465));
    InMux I__5072 (
            .O(N__23469),
            .I(N__23462));
    InMux I__5071 (
            .O(N__23468),
            .I(N__23459));
    LocalMux I__5070 (
            .O(N__23465),
            .I(N__23456));
    LocalMux I__5069 (
            .O(N__23462),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__5068 (
            .O(N__23459),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__5067 (
            .O(N__23456),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__5066 (
            .O(N__23449),
            .I(N__23444));
    InMux I__5065 (
            .O(N__23448),
            .I(N__23441));
    InMux I__5064 (
            .O(N__23447),
            .I(N__23438));
    LocalMux I__5063 (
            .O(N__23444),
            .I(N__23435));
    LocalMux I__5062 (
            .O(N__23441),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__5061 (
            .O(N__23438),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__5060 (
            .O(N__23435),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    CascadeMux I__5059 (
            .O(N__23428),
            .I(N__23423));
    InMux I__5058 (
            .O(N__23427),
            .I(N__23420));
    InMux I__5057 (
            .O(N__23426),
            .I(N__23417));
    InMux I__5056 (
            .O(N__23423),
            .I(N__23414));
    LocalMux I__5055 (
            .O(N__23420),
            .I(N__23411));
    LocalMux I__5054 (
            .O(N__23417),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__5053 (
            .O(N__23414),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv4 I__5052 (
            .O(N__23411),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__5051 (
            .O(N__23404),
            .I(N__23399));
    InMux I__5050 (
            .O(N__23403),
            .I(N__23396));
    InMux I__5049 (
            .O(N__23402),
            .I(N__23393));
    LocalMux I__5048 (
            .O(N__23399),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__5047 (
            .O(N__23396),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__5046 (
            .O(N__23393),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__5045 (
            .O(N__23386),
            .I(N__23382));
    InMux I__5044 (
            .O(N__23385),
            .I(N__23379));
    LocalMux I__5043 (
            .O(N__23382),
            .I(N__23376));
    LocalMux I__5042 (
            .O(N__23379),
            .I(N__23373));
    Span4Mux_h I__5041 (
            .O(N__23376),
            .I(N__23370));
    Odrv4 I__5040 (
            .O(N__23373),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    Odrv4 I__5039 (
            .O(N__23370),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    InMux I__5038 (
            .O(N__23365),
            .I(N__23362));
    LocalMux I__5037 (
            .O(N__23362),
            .I(uart_input_pc_c));
    InMux I__5036 (
            .O(N__23359),
            .I(N__23356));
    LocalMux I__5035 (
            .O(N__23356),
            .I(\uart_pc_sync.aux_0__0__0_0 ));
    InMux I__5034 (
            .O(N__23353),
            .I(N__23350));
    LocalMux I__5033 (
            .O(N__23350),
            .I(N__23347));
    Odrv4 I__5032 (
            .O(N__23347),
            .I(\uart_pc_sync.aux_1__0__0_0 ));
    CascadeMux I__5031 (
            .O(N__23344),
            .I(N__23341));
    InMux I__5030 (
            .O(N__23341),
            .I(N__23335));
    InMux I__5029 (
            .O(N__23340),
            .I(N__23335));
    LocalMux I__5028 (
            .O(N__23335),
            .I(frame_decoder_OFF2data_7));
    CascadeMux I__5027 (
            .O(N__23332),
            .I(N__23329));
    InMux I__5026 (
            .O(N__23329),
            .I(N__23326));
    LocalMux I__5025 (
            .O(N__23326),
            .I(frame_decoder_OFF2data_1));
    CascadeMux I__5024 (
            .O(N__23323),
            .I(N__23320));
    InMux I__5023 (
            .O(N__23320),
            .I(N__23317));
    LocalMux I__5022 (
            .O(N__23317),
            .I(frame_decoder_OFF2data_4));
    InMux I__5021 (
            .O(N__23314),
            .I(N__23309));
    InMux I__5020 (
            .O(N__23313),
            .I(N__23306));
    InMux I__5019 (
            .O(N__23312),
            .I(N__23303));
    LocalMux I__5018 (
            .O(N__23309),
            .I(N__23300));
    LocalMux I__5017 (
            .O(N__23306),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__5016 (
            .O(N__23303),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__5015 (
            .O(N__23300),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__5014 (
            .O(N__23293),
            .I(N__23290));
    LocalMux I__5013 (
            .O(N__23290),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ));
    CascadeMux I__5012 (
            .O(N__23287),
            .I(N__23283));
    InMux I__5011 (
            .O(N__23286),
            .I(N__23279));
    InMux I__5010 (
            .O(N__23283),
            .I(N__23276));
    InMux I__5009 (
            .O(N__23282),
            .I(N__23273));
    LocalMux I__5008 (
            .O(N__23279),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5007 (
            .O(N__23276),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5006 (
            .O(N__23273),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    CascadeMux I__5005 (
            .O(N__23266),
            .I(N__23263));
    InMux I__5004 (
            .O(N__23263),
            .I(N__23260));
    LocalMux I__5003 (
            .O(N__23260),
            .I(N__23257));
    Odrv4 I__5002 (
            .O(N__23257),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__5001 (
            .O(N__23254),
            .I(N__23249));
    InMux I__5000 (
            .O(N__23253),
            .I(N__23246));
    InMux I__4999 (
            .O(N__23252),
            .I(N__23243));
    LocalMux I__4998 (
            .O(N__23249),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__4997 (
            .O(N__23246),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__4996 (
            .O(N__23243),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__4995 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__4994 (
            .O(N__23233),
            .I(N__23230));
    Odrv12 I__4993 (
            .O(N__23230),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__4992 (
            .O(N__23227),
            .I(N__23224));
    LocalMux I__4991 (
            .O(N__23224),
            .I(N__23221));
    Span4Mux_v I__4990 (
            .O(N__23221),
            .I(N__23218));
    Span4Mux_h I__4989 (
            .O(N__23218),
            .I(N__23215));
    Span4Mux_v I__4988 (
            .O(N__23215),
            .I(N__23212));
    Odrv4 I__4987 (
            .O(N__23212),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__4986 (
            .O(N__23209),
            .I(N__23206));
    LocalMux I__4985 (
            .O(N__23206),
            .I(N__23203));
    Odrv4 I__4984 (
            .O(N__23203),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__4983 (
            .O(N__23200),
            .I(N__23197));
    LocalMux I__4982 (
            .O(N__23197),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__4981 (
            .O(N__23194),
            .I(N__23191));
    LocalMux I__4980 (
            .O(N__23191),
            .I(N__23188));
    Span4Mux_s2_v I__4979 (
            .O(N__23188),
            .I(N__23185));
    Span4Mux_v I__4978 (
            .O(N__23185),
            .I(N__23182));
    Odrv4 I__4977 (
            .O(N__23182),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__4976 (
            .O(N__23179),
            .I(N__23176));
    LocalMux I__4975 (
            .O(N__23176),
            .I(N__23173));
    Odrv4 I__4974 (
            .O(N__23173),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    CascadeMux I__4973 (
            .O(N__23170),
            .I(N__23167));
    InMux I__4972 (
            .O(N__23167),
            .I(N__23164));
    LocalMux I__4971 (
            .O(N__23164),
            .I(N__23161));
    Odrv4 I__4970 (
            .O(N__23161),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__4969 (
            .O(N__23158),
            .I(N__23155));
    LocalMux I__4968 (
            .O(N__23155),
            .I(N__23152));
    Span4Mux_v I__4967 (
            .O(N__23152),
            .I(N__23149));
    Odrv4 I__4966 (
            .O(N__23149),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    InMux I__4965 (
            .O(N__23146),
            .I(N__23143));
    LocalMux I__4964 (
            .O(N__23143),
            .I(N__23140));
    Odrv4 I__4963 (
            .O(N__23140),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__4962 (
            .O(N__23137),
            .I(N__23128));
    InMux I__4961 (
            .O(N__23136),
            .I(N__23128));
    InMux I__4960 (
            .O(N__23135),
            .I(N__23128));
    LocalMux I__4959 (
            .O(N__23128),
            .I(N__23120));
    InMux I__4958 (
            .O(N__23127),
            .I(N__23117));
    InMux I__4957 (
            .O(N__23126),
            .I(N__23108));
    InMux I__4956 (
            .O(N__23125),
            .I(N__23108));
    InMux I__4955 (
            .O(N__23124),
            .I(N__23108));
    InMux I__4954 (
            .O(N__23123),
            .I(N__23108));
    Span4Mux_s3_v I__4953 (
            .O(N__23120),
            .I(N__23101));
    LocalMux I__4952 (
            .O(N__23117),
            .I(N__23101));
    LocalMux I__4951 (
            .O(N__23108),
            .I(N__23098));
    InMux I__4950 (
            .O(N__23107),
            .I(N__23088));
    InMux I__4949 (
            .O(N__23106),
            .I(N__23088));
    Span4Mux_h I__4948 (
            .O(N__23101),
            .I(N__23083));
    Span4Mux_s3_v I__4947 (
            .O(N__23098),
            .I(N__23083));
    InMux I__4946 (
            .O(N__23097),
            .I(N__23072));
    InMux I__4945 (
            .O(N__23096),
            .I(N__23072));
    InMux I__4944 (
            .O(N__23095),
            .I(N__23072));
    InMux I__4943 (
            .O(N__23094),
            .I(N__23072));
    InMux I__4942 (
            .O(N__23093),
            .I(N__23072));
    LocalMux I__4941 (
            .O(N__23088),
            .I(N__23069));
    Odrv4 I__4940 (
            .O(N__23083),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__4939 (
            .O(N__23072),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv12 I__4938 (
            .O(N__23069),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    CEMux I__4937 (
            .O(N__23062),
            .I(N__23057));
    CEMux I__4936 (
            .O(N__23061),
            .I(N__23053));
    CEMux I__4935 (
            .O(N__23060),
            .I(N__23049));
    LocalMux I__4934 (
            .O(N__23057),
            .I(N__23046));
    CEMux I__4933 (
            .O(N__23056),
            .I(N__23043));
    LocalMux I__4932 (
            .O(N__23053),
            .I(N__23040));
    CEMux I__4931 (
            .O(N__23052),
            .I(N__23037));
    LocalMux I__4930 (
            .O(N__23049),
            .I(N__23034));
    Span4Mux_h I__4929 (
            .O(N__23046),
            .I(N__23029));
    LocalMux I__4928 (
            .O(N__23043),
            .I(N__23029));
    Span4Mux_s3_v I__4927 (
            .O(N__23040),
            .I(N__23026));
    LocalMux I__4926 (
            .O(N__23037),
            .I(N__23023));
    Span4Mux_h I__4925 (
            .O(N__23034),
            .I(N__23020));
    Span4Mux_s3_v I__4924 (
            .O(N__23029),
            .I(N__23015));
    Span4Mux_h I__4923 (
            .O(N__23026),
            .I(N__23015));
    Span4Mux_h I__4922 (
            .O(N__23023),
            .I(N__23010));
    Span4Mux_s2_v I__4921 (
            .O(N__23020),
            .I(N__23010));
    Span4Mux_h I__4920 (
            .O(N__23015),
            .I(N__23007));
    Odrv4 I__4919 (
            .O(N__23010),
            .I(\ppm_encoder_1.N_590_0 ));
    Odrv4 I__4918 (
            .O(N__23007),
            .I(\ppm_encoder_1.N_590_0 ));
    InMux I__4917 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__4916 (
            .O(N__22999),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    InMux I__4915 (
            .O(N__22996),
            .I(N__22991));
    InMux I__4914 (
            .O(N__22995),
            .I(N__22988));
    InMux I__4913 (
            .O(N__22994),
            .I(N__22985));
    LocalMux I__4912 (
            .O(N__22991),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__4911 (
            .O(N__22988),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__4910 (
            .O(N__22985),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__4909 (
            .O(N__22978),
            .I(N__22975));
    LocalMux I__4908 (
            .O(N__22975),
            .I(N__22972));
    Odrv12 I__4907 (
            .O(N__22972),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__4906 (
            .O(N__22969),
            .I(N__22965));
    InMux I__4905 (
            .O(N__22968),
            .I(N__22962));
    LocalMux I__4904 (
            .O(N__22965),
            .I(N__22959));
    LocalMux I__4903 (
            .O(N__22962),
            .I(N__22956));
    Span12Mux_h I__4902 (
            .O(N__22959),
            .I(N__22952));
    Span4Mux_v I__4901 (
            .O(N__22956),
            .I(N__22949));
    InMux I__4900 (
            .O(N__22955),
            .I(N__22946));
    Odrv12 I__4899 (
            .O(N__22952),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__4898 (
            .O(N__22949),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__4897 (
            .O(N__22946),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__4896 (
            .O(N__22939),
            .I(N__22935));
    InMux I__4895 (
            .O(N__22938),
            .I(N__22932));
    LocalMux I__4894 (
            .O(N__22935),
            .I(N__22929));
    LocalMux I__4893 (
            .O(N__22932),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    Odrv12 I__4892 (
            .O(N__22929),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    InMux I__4891 (
            .O(N__22924),
            .I(N__22921));
    LocalMux I__4890 (
            .O(N__22921),
            .I(N__22918));
    Span4Mux_s2_v I__4889 (
            .O(N__22918),
            .I(N__22915));
    Span4Mux_h I__4888 (
            .O(N__22915),
            .I(N__22910));
    InMux I__4887 (
            .O(N__22914),
            .I(N__22907));
    InMux I__4886 (
            .O(N__22913),
            .I(N__22904));
    Odrv4 I__4885 (
            .O(N__22910),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__4884 (
            .O(N__22907),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__4883 (
            .O(N__22904),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__4882 (
            .O(N__22897),
            .I(N__22893));
    CascadeMux I__4881 (
            .O(N__22896),
            .I(N__22890));
    InMux I__4880 (
            .O(N__22893),
            .I(N__22887));
    InMux I__4879 (
            .O(N__22890),
            .I(N__22884));
    LocalMux I__4878 (
            .O(N__22887),
            .I(N__22881));
    LocalMux I__4877 (
            .O(N__22884),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    Odrv4 I__4876 (
            .O(N__22881),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__4875 (
            .O(N__22876),
            .I(N__22869));
    InMux I__4874 (
            .O(N__22875),
            .I(N__22869));
    InMux I__4873 (
            .O(N__22874),
            .I(N__22866));
    LocalMux I__4872 (
            .O(N__22869),
            .I(N__22863));
    LocalMux I__4871 (
            .O(N__22866),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    Odrv12 I__4870 (
            .O(N__22863),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__4869 (
            .O(N__22858),
            .I(N__22852));
    InMux I__4868 (
            .O(N__22857),
            .I(N__22843));
    InMux I__4867 (
            .O(N__22856),
            .I(N__22838));
    InMux I__4866 (
            .O(N__22855),
            .I(N__22838));
    LocalMux I__4865 (
            .O(N__22852),
            .I(N__22835));
    InMux I__4864 (
            .O(N__22851),
            .I(N__22832));
    InMux I__4863 (
            .O(N__22850),
            .I(N__22829));
    InMux I__4862 (
            .O(N__22849),
            .I(N__22823));
    InMux I__4861 (
            .O(N__22848),
            .I(N__22823));
    InMux I__4860 (
            .O(N__22847),
            .I(N__22820));
    CascadeMux I__4859 (
            .O(N__22846),
            .I(N__22817));
    LocalMux I__4858 (
            .O(N__22843),
            .I(N__22810));
    LocalMux I__4857 (
            .O(N__22838),
            .I(N__22810));
    Span4Mux_v I__4856 (
            .O(N__22835),
            .I(N__22803));
    LocalMux I__4855 (
            .O(N__22832),
            .I(N__22803));
    LocalMux I__4854 (
            .O(N__22829),
            .I(N__22803));
    InMux I__4853 (
            .O(N__22828),
            .I(N__22800));
    LocalMux I__4852 (
            .O(N__22823),
            .I(N__22795));
    LocalMux I__4851 (
            .O(N__22820),
            .I(N__22792));
    InMux I__4850 (
            .O(N__22817),
            .I(N__22785));
    InMux I__4849 (
            .O(N__22816),
            .I(N__22785));
    InMux I__4848 (
            .O(N__22815),
            .I(N__22785));
    Span4Mux_v I__4847 (
            .O(N__22810),
            .I(N__22782));
    Span4Mux_v I__4846 (
            .O(N__22803),
            .I(N__22779));
    LocalMux I__4845 (
            .O(N__22800),
            .I(N__22776));
    InMux I__4844 (
            .O(N__22799),
            .I(N__22773));
    InMux I__4843 (
            .O(N__22798),
            .I(N__22769));
    Span4Mux_v I__4842 (
            .O(N__22795),
            .I(N__22764));
    Span4Mux_h I__4841 (
            .O(N__22792),
            .I(N__22764));
    LocalMux I__4840 (
            .O(N__22785),
            .I(N__22758));
    Span4Mux_v I__4839 (
            .O(N__22782),
            .I(N__22749));
    Span4Mux_h I__4838 (
            .O(N__22779),
            .I(N__22749));
    Span4Mux_h I__4837 (
            .O(N__22776),
            .I(N__22749));
    LocalMux I__4836 (
            .O(N__22773),
            .I(N__22749));
    InMux I__4835 (
            .O(N__22772),
            .I(N__22746));
    LocalMux I__4834 (
            .O(N__22769),
            .I(N__22741));
    Span4Mux_h I__4833 (
            .O(N__22764),
            .I(N__22741));
    InMux I__4832 (
            .O(N__22763),
            .I(N__22738));
    InMux I__4831 (
            .O(N__22762),
            .I(N__22733));
    InMux I__4830 (
            .O(N__22761),
            .I(N__22733));
    Span4Mux_h I__4829 (
            .O(N__22758),
            .I(N__22730));
    Odrv4 I__4828 (
            .O(N__22749),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__4827 (
            .O(N__22746),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__4826 (
            .O(N__22741),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__4825 (
            .O(N__22738),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__4824 (
            .O(N__22733),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__4823 (
            .O(N__22730),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__4822 (
            .O(N__22717),
            .I(N__22714));
    LocalMux I__4821 (
            .O(N__22714),
            .I(N__22709));
    InMux I__4820 (
            .O(N__22713),
            .I(N__22706));
    CascadeMux I__4819 (
            .O(N__22712),
            .I(N__22703));
    Span4Mux_v I__4818 (
            .O(N__22709),
            .I(N__22700));
    LocalMux I__4817 (
            .O(N__22706),
            .I(N__22697));
    InMux I__4816 (
            .O(N__22703),
            .I(N__22694));
    Span4Mux_h I__4815 (
            .O(N__22700),
            .I(N__22689));
    Span4Mux_v I__4814 (
            .O(N__22697),
            .I(N__22689));
    LocalMux I__4813 (
            .O(N__22694),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__4812 (
            .O(N__22689),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__4811 (
            .O(N__22684),
            .I(N__22680));
    InMux I__4810 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__4809 (
            .O(N__22680),
            .I(N__22673));
    LocalMux I__4808 (
            .O(N__22677),
            .I(N__22670));
    InMux I__4807 (
            .O(N__22676),
            .I(N__22667));
    Span4Mux_v I__4806 (
            .O(N__22673),
            .I(N__22662));
    Span4Mux_h I__4805 (
            .O(N__22670),
            .I(N__22662));
    LocalMux I__4804 (
            .O(N__22667),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__4803 (
            .O(N__22662),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__4802 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__4801 (
            .O(N__22654),
            .I(\ppm_encoder_1.N_301 ));
    InMux I__4800 (
            .O(N__22651),
            .I(N__22648));
    LocalMux I__4799 (
            .O(N__22648),
            .I(N__22645));
    Span4Mux_v I__4798 (
            .O(N__22645),
            .I(N__22642));
    Odrv4 I__4797 (
            .O(N__22642),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__4796 (
            .O(N__22639),
            .I(N__22636));
    LocalMux I__4795 (
            .O(N__22636),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    InMux I__4794 (
            .O(N__22633),
            .I(N__22628));
    InMux I__4793 (
            .O(N__22632),
            .I(N__22625));
    InMux I__4792 (
            .O(N__22631),
            .I(N__22622));
    LocalMux I__4791 (
            .O(N__22628),
            .I(N__22619));
    LocalMux I__4790 (
            .O(N__22625),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__4789 (
            .O(N__22622),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    Odrv4 I__4788 (
            .O(N__22619),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__4787 (
            .O(N__22612),
            .I(N__22607));
    InMux I__4786 (
            .O(N__22611),
            .I(N__22604));
    InMux I__4785 (
            .O(N__22610),
            .I(N__22601));
    LocalMux I__4784 (
            .O(N__22607),
            .I(N__22598));
    LocalMux I__4783 (
            .O(N__22604),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__4782 (
            .O(N__22601),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__4781 (
            .O(N__22598),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__4780 (
            .O(N__22591),
            .I(N__22586));
    InMux I__4779 (
            .O(N__22590),
            .I(N__22583));
    InMux I__4778 (
            .O(N__22589),
            .I(N__22580));
    LocalMux I__4777 (
            .O(N__22586),
            .I(N__22577));
    LocalMux I__4776 (
            .O(N__22583),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__4775 (
            .O(N__22580),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv12 I__4774 (
            .O(N__22577),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__4773 (
            .O(N__22570),
            .I(N__22565));
    InMux I__4772 (
            .O(N__22569),
            .I(N__22562));
    InMux I__4771 (
            .O(N__22568),
            .I(N__22559));
    LocalMux I__4770 (
            .O(N__22565),
            .I(N__22556));
    LocalMux I__4769 (
            .O(N__22562),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__4768 (
            .O(N__22559),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__4767 (
            .O(N__22556),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    CascadeMux I__4766 (
            .O(N__22549),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ));
    InMux I__4765 (
            .O(N__22546),
            .I(N__22543));
    LocalMux I__4764 (
            .O(N__22543),
            .I(N__22540));
    Span4Mux_s2_v I__4763 (
            .O(N__22540),
            .I(N__22537));
    Odrv4 I__4762 (
            .O(N__22537),
            .I(\ppm_encoder_1.N_144_17 ));
    InMux I__4761 (
            .O(N__22534),
            .I(N__22531));
    LocalMux I__4760 (
            .O(N__22531),
            .I(N__22528));
    Odrv4 I__4759 (
            .O(N__22528),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    InMux I__4758 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__4757 (
            .O(N__22522),
            .I(N__22519));
    Span4Mux_h I__4756 (
            .O(N__22519),
            .I(N__22516));
    Odrv4 I__4755 (
            .O(N__22516),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    CascadeMux I__4754 (
            .O(N__22513),
            .I(\ppm_encoder_1.N_144_17_cascade_ ));
    InMux I__4753 (
            .O(N__22510),
            .I(N__22507));
    LocalMux I__4752 (
            .O(N__22507),
            .I(N__22504));
    Span4Mux_h I__4751 (
            .O(N__22504),
            .I(N__22501));
    Span4Mux_v I__4750 (
            .O(N__22501),
            .I(N__22498));
    Odrv4 I__4749 (
            .O(N__22498),
            .I(\ppm_encoder_1.N_144 ));
    InMux I__4748 (
            .O(N__22495),
            .I(N__22492));
    LocalMux I__4747 (
            .O(N__22492),
            .I(N__22489));
    Span4Mux_h I__4746 (
            .O(N__22489),
            .I(N__22486));
    Span4Mux_v I__4745 (
            .O(N__22486),
            .I(N__22483));
    Odrv4 I__4744 (
            .O(N__22483),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__4743 (
            .O(N__22480),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__4742 (
            .O(N__22477),
            .I(N__22474));
    LocalMux I__4741 (
            .O(N__22474),
            .I(N__22471));
    Span12Mux_s8_h I__4740 (
            .O(N__22471),
            .I(N__22468));
    Odrv12 I__4739 (
            .O(N__22468),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__4738 (
            .O(N__22465),
            .I(\ppm_encoder_1.un1_aileron_cry_7 ));
    InMux I__4737 (
            .O(N__22462),
            .I(N__22459));
    LocalMux I__4736 (
            .O(N__22459),
            .I(N__22456));
    Odrv4 I__4735 (
            .O(N__22456),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__4734 (
            .O(N__22453),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__4733 (
            .O(N__22450),
            .I(N__22447));
    LocalMux I__4732 (
            .O(N__22447),
            .I(N__22444));
    Span4Mux_h I__4731 (
            .O(N__22444),
            .I(N__22441));
    Odrv4 I__4730 (
            .O(N__22441),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__4729 (
            .O(N__22438),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__4728 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__4727 (
            .O(N__22432),
            .I(N__22429));
    Span4Mux_v I__4726 (
            .O(N__22429),
            .I(N__22426));
    Odrv4 I__4725 (
            .O(N__22426),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__4724 (
            .O(N__22423),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__4723 (
            .O(N__22420),
            .I(N__22417));
    LocalMux I__4722 (
            .O(N__22417),
            .I(N__22414));
    Span4Mux_h I__4721 (
            .O(N__22414),
            .I(N__22411));
    Span4Mux_h I__4720 (
            .O(N__22411),
            .I(N__22408));
    Odrv4 I__4719 (
            .O(N__22408),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__4718 (
            .O(N__22405),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__4717 (
            .O(N__22402),
            .I(N__22399));
    LocalMux I__4716 (
            .O(N__22399),
            .I(N__22396));
    Odrv4 I__4715 (
            .O(N__22396),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__4714 (
            .O(N__22393),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__4713 (
            .O(N__22390),
            .I(bfn_8_20_0_));
    InMux I__4712 (
            .O(N__22387),
            .I(N__22383));
    InMux I__4711 (
            .O(N__22386),
            .I(N__22380));
    LocalMux I__4710 (
            .O(N__22383),
            .I(N__22377));
    LocalMux I__4709 (
            .O(N__22380),
            .I(N__22374));
    Span4Mux_h I__4708 (
            .O(N__22377),
            .I(N__22371));
    Span4Mux_v I__4707 (
            .O(N__22374),
            .I(N__22368));
    Span4Mux_v I__4706 (
            .O(N__22371),
            .I(N__22365));
    Odrv4 I__4705 (
            .O(N__22368),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    Odrv4 I__4704 (
            .O(N__22365),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    InMux I__4703 (
            .O(N__22360),
            .I(N__22357));
    LocalMux I__4702 (
            .O(N__22357),
            .I(N__22354));
    Span4Mux_h I__4701 (
            .O(N__22354),
            .I(N__22351));
    Odrv4 I__4700 (
            .O(N__22351),
            .I(\Commands_frame_decoder.state_1_RNO_4Z0Z_0 ));
    CascadeMux I__4699 (
            .O(N__22348),
            .I(N__22345));
    InMux I__4698 (
            .O(N__22345),
            .I(N__22342));
    LocalMux I__4697 (
            .O(N__22342),
            .I(N__22339));
    Span4Mux_h I__4696 (
            .O(N__22339),
            .I(N__22334));
    InMux I__4695 (
            .O(N__22338),
            .I(N__22331));
    InMux I__4694 (
            .O(N__22337),
            .I(N__22327));
    Span4Mux_h I__4693 (
            .O(N__22334),
            .I(N__22324));
    LocalMux I__4692 (
            .O(N__22331),
            .I(N__22321));
    InMux I__4691 (
            .O(N__22330),
            .I(N__22318));
    LocalMux I__4690 (
            .O(N__22327),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__4689 (
            .O(N__22324),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__4688 (
            .O(N__22321),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4687 (
            .O(N__22318),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__4686 (
            .O(N__22309),
            .I(N__22306));
    LocalMux I__4685 (
            .O(N__22306),
            .I(N__22302));
    InMux I__4684 (
            .O(N__22305),
            .I(N__22299));
    Span4Mux_v I__4683 (
            .O(N__22302),
            .I(N__22295));
    LocalMux I__4682 (
            .O(N__22299),
            .I(N__22292));
    InMux I__4681 (
            .O(N__22298),
            .I(N__22289));
    Odrv4 I__4680 (
            .O(N__22295),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    Odrv4 I__4679 (
            .O(N__22292),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    LocalMux I__4678 (
            .O(N__22289),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    InMux I__4677 (
            .O(N__22282),
            .I(N__22279));
    LocalMux I__4676 (
            .O(N__22279),
            .I(N__22276));
    Odrv12 I__4675 (
            .O(N__22276),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__4674 (
            .O(N__22273),
            .I(N__22268));
    InMux I__4673 (
            .O(N__22272),
            .I(N__22265));
    InMux I__4672 (
            .O(N__22271),
            .I(N__22262));
    LocalMux I__4671 (
            .O(N__22268),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__4670 (
            .O(N__22265),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__4669 (
            .O(N__22262),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__4668 (
            .O(N__22255),
            .I(N__22252));
    LocalMux I__4667 (
            .O(N__22252),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    InMux I__4666 (
            .O(N__22249),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__4665 (
            .O(N__22246),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__4664 (
            .O(N__22243),
            .I(N__22232));
    InMux I__4663 (
            .O(N__22242),
            .I(N__22232));
    InMux I__4662 (
            .O(N__22241),
            .I(N__22227));
    CascadeMux I__4661 (
            .O(N__22240),
            .I(N__22224));
    CascadeMux I__4660 (
            .O(N__22239),
            .I(N__22221));
    CascadeMux I__4659 (
            .O(N__22238),
            .I(N__22218));
    CascadeMux I__4658 (
            .O(N__22237),
            .I(N__22215));
    LocalMux I__4657 (
            .O(N__22232),
            .I(N__22212));
    InMux I__4656 (
            .O(N__22231),
            .I(N__22207));
    InMux I__4655 (
            .O(N__22230),
            .I(N__22207));
    LocalMux I__4654 (
            .O(N__22227),
            .I(N__22204));
    InMux I__4653 (
            .O(N__22224),
            .I(N__22199));
    InMux I__4652 (
            .O(N__22221),
            .I(N__22199));
    InMux I__4651 (
            .O(N__22218),
            .I(N__22194));
    InMux I__4650 (
            .O(N__22215),
            .I(N__22194));
    Odrv4 I__4649 (
            .O(N__22212),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4648 (
            .O(N__22207),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__4647 (
            .O(N__22204),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4646 (
            .O(N__22199),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4645 (
            .O(N__22194),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__4644 (
            .O(N__22183),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__4643 (
            .O(N__22180),
            .I(N__22177));
    LocalMux I__4642 (
            .O(N__22177),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    CascadeMux I__4641 (
            .O(N__22174),
            .I(N__22170));
    CascadeMux I__4640 (
            .O(N__22173),
            .I(N__22166));
    InMux I__4639 (
            .O(N__22170),
            .I(N__22162));
    InMux I__4638 (
            .O(N__22169),
            .I(N__22155));
    InMux I__4637 (
            .O(N__22166),
            .I(N__22155));
    InMux I__4636 (
            .O(N__22165),
            .I(N__22155));
    LocalMux I__4635 (
            .O(N__22162),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4634 (
            .O(N__22155),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__4633 (
            .O(N__22150),
            .I(N__22144));
    InMux I__4632 (
            .O(N__22149),
            .I(N__22144));
    LocalMux I__4631 (
            .O(N__22144),
            .I(N__22141));
    Odrv4 I__4630 (
            .O(N__22141),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    CascadeMux I__4629 (
            .O(N__22138),
            .I(N__22135));
    InMux I__4628 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__4627 (
            .O(N__22132),
            .I(N__22129));
    Odrv4 I__4626 (
            .O(N__22129),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1 ));
    InMux I__4625 (
            .O(N__22126),
            .I(N__22123));
    LocalMux I__4624 (
            .O(N__22123),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    InMux I__4623 (
            .O(N__22120),
            .I(N__22113));
    InMux I__4622 (
            .O(N__22119),
            .I(N__22110));
    InMux I__4621 (
            .O(N__22118),
            .I(N__22107));
    InMux I__4620 (
            .O(N__22117),
            .I(N__22102));
    InMux I__4619 (
            .O(N__22116),
            .I(N__22102));
    LocalMux I__4618 (
            .O(N__22113),
            .I(\uart_pc.N_143 ));
    LocalMux I__4617 (
            .O(N__22110),
            .I(\uart_pc.N_143 ));
    LocalMux I__4616 (
            .O(N__22107),
            .I(\uart_pc.N_143 ));
    LocalMux I__4615 (
            .O(N__22102),
            .I(\uart_pc.N_143 ));
    CascadeMux I__4614 (
            .O(N__22093),
            .I(N__22088));
    CascadeMux I__4613 (
            .O(N__22092),
            .I(N__22085));
    InMux I__4612 (
            .O(N__22091),
            .I(N__22080));
    InMux I__4611 (
            .O(N__22088),
            .I(N__22077));
    InMux I__4610 (
            .O(N__22085),
            .I(N__22074));
    InMux I__4609 (
            .O(N__22084),
            .I(N__22069));
    InMux I__4608 (
            .O(N__22083),
            .I(N__22069));
    LocalMux I__4607 (
            .O(N__22080),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4606 (
            .O(N__22077),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4605 (
            .O(N__22074),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4604 (
            .O(N__22069),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__4603 (
            .O(N__22060),
            .I(N__22057));
    LocalMux I__4602 (
            .O(N__22057),
            .I(N__22047));
    InMux I__4601 (
            .O(N__22056),
            .I(N__22044));
    InMux I__4600 (
            .O(N__22055),
            .I(N__22035));
    InMux I__4599 (
            .O(N__22054),
            .I(N__22035));
    InMux I__4598 (
            .O(N__22053),
            .I(N__22035));
    InMux I__4597 (
            .O(N__22052),
            .I(N__22035));
    InMux I__4596 (
            .O(N__22051),
            .I(N__22030));
    InMux I__4595 (
            .O(N__22050),
            .I(N__22030));
    Odrv4 I__4594 (
            .O(N__22047),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4593 (
            .O(N__22044),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4592 (
            .O(N__22035),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4591 (
            .O(N__22030),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__4590 (
            .O(N__22021),
            .I(N__22016));
    InMux I__4589 (
            .O(N__22020),
            .I(N__22011));
    InMux I__4588 (
            .O(N__22019),
            .I(N__22008));
    LocalMux I__4587 (
            .O(N__22016),
            .I(N__22005));
    InMux I__4586 (
            .O(N__22015),
            .I(N__22000));
    InMux I__4585 (
            .O(N__22014),
            .I(N__22000));
    LocalMux I__4584 (
            .O(N__22011),
            .I(N__21995));
    LocalMux I__4583 (
            .O(N__22008),
            .I(N__21992));
    Span4Mux_v I__4582 (
            .O(N__22005),
            .I(N__21986));
    LocalMux I__4581 (
            .O(N__22000),
            .I(N__21986));
    CascadeMux I__4580 (
            .O(N__21999),
            .I(N__21982));
    InMux I__4579 (
            .O(N__21998),
            .I(N__21979));
    Span4Mux_h I__4578 (
            .O(N__21995),
            .I(N__21976));
    Span4Mux_h I__4577 (
            .O(N__21992),
            .I(N__21973));
    InMux I__4576 (
            .O(N__21991),
            .I(N__21970));
    Span4Mux_h I__4575 (
            .O(N__21986),
            .I(N__21967));
    InMux I__4574 (
            .O(N__21985),
            .I(N__21962));
    InMux I__4573 (
            .O(N__21982),
            .I(N__21962));
    LocalMux I__4572 (
            .O(N__21979),
            .I(N__21959));
    Odrv4 I__4571 (
            .O(N__21976),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__4570 (
            .O(N__21973),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__4569 (
            .O(N__21970),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__4568 (
            .O(N__21967),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__4567 (
            .O(N__21962),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv12 I__4566 (
            .O(N__21959),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__4565 (
            .O(N__21946),
            .I(N__21938));
    InMux I__4564 (
            .O(N__21945),
            .I(N__21938));
    InMux I__4563 (
            .O(N__21944),
            .I(N__21935));
    InMux I__4562 (
            .O(N__21943),
            .I(N__21932));
    LocalMux I__4561 (
            .O(N__21938),
            .I(N__21928));
    LocalMux I__4560 (
            .O(N__21935),
            .I(N__21923));
    LocalMux I__4559 (
            .O(N__21932),
            .I(N__21923));
    InMux I__4558 (
            .O(N__21931),
            .I(N__21919));
    Span4Mux_h I__4557 (
            .O(N__21928),
            .I(N__21914));
    Span4Mux_h I__4556 (
            .O(N__21923),
            .I(N__21911));
    InMux I__4555 (
            .O(N__21922),
            .I(N__21908));
    LocalMux I__4554 (
            .O(N__21919),
            .I(N__21905));
    InMux I__4553 (
            .O(N__21918),
            .I(N__21900));
    InMux I__4552 (
            .O(N__21917),
            .I(N__21900));
    Odrv4 I__4551 (
            .O(N__21914),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__4550 (
            .O(N__21911),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__4549 (
            .O(N__21908),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv12 I__4548 (
            .O(N__21905),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__4547 (
            .O(N__21900),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__4546 (
            .O(N__21889),
            .I(N__21882));
    InMux I__4545 (
            .O(N__21888),
            .I(N__21882));
    InMux I__4544 (
            .O(N__21887),
            .I(N__21877));
    LocalMux I__4543 (
            .O(N__21882),
            .I(N__21873));
    InMux I__4542 (
            .O(N__21881),
            .I(N__21870));
    InMux I__4541 (
            .O(N__21880),
            .I(N__21867));
    LocalMux I__4540 (
            .O(N__21877),
            .I(N__21864));
    InMux I__4539 (
            .O(N__21876),
            .I(N__21861));
    Span4Mux_h I__4538 (
            .O(N__21873),
            .I(N__21858));
    LocalMux I__4537 (
            .O(N__21870),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__4536 (
            .O(N__21867),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__4535 (
            .O(N__21864),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__4534 (
            .O(N__21861),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__4533 (
            .O(N__21858),
            .I(\uart_drone.stateZ0Z_4 ));
    InMux I__4532 (
            .O(N__21847),
            .I(N__21844));
    LocalMux I__4531 (
            .O(N__21844),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__4530 (
            .O(N__21841),
            .I(N__21837));
    CascadeMux I__4529 (
            .O(N__21840),
            .I(N__21834));
    LocalMux I__4528 (
            .O(N__21837),
            .I(N__21831));
    InMux I__4527 (
            .O(N__21834),
            .I(N__21828));
    Odrv12 I__4526 (
            .O(N__21831),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__4525 (
            .O(N__21828),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    InMux I__4524 (
            .O(N__21823),
            .I(N__21820));
    LocalMux I__4523 (
            .O(N__21820),
            .I(N__21817));
    Odrv12 I__4522 (
            .O(N__21817),
            .I(\uart_drone.data_Auxce_0_3 ));
    InMux I__4521 (
            .O(N__21814),
            .I(N__21810));
    CascadeMux I__4520 (
            .O(N__21813),
            .I(N__21807));
    LocalMux I__4519 (
            .O(N__21810),
            .I(N__21804));
    InMux I__4518 (
            .O(N__21807),
            .I(N__21801));
    Odrv12 I__4517 (
            .O(N__21804),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__4516 (
            .O(N__21801),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__4515 (
            .O(N__21796),
            .I(N__21781));
    InMux I__4514 (
            .O(N__21795),
            .I(N__21781));
    InMux I__4513 (
            .O(N__21794),
            .I(N__21781));
    InMux I__4512 (
            .O(N__21793),
            .I(N__21781));
    InMux I__4511 (
            .O(N__21792),
            .I(N__21781));
    LocalMux I__4510 (
            .O(N__21781),
            .I(N__21778));
    Span4Mux_h I__4509 (
            .O(N__21778),
            .I(N__21772));
    InMux I__4508 (
            .O(N__21777),
            .I(N__21765));
    InMux I__4507 (
            .O(N__21776),
            .I(N__21765));
    InMux I__4506 (
            .O(N__21775),
            .I(N__21765));
    Odrv4 I__4505 (
            .O(N__21772),
            .I(\uart_drone.un1_state_2_0 ));
    LocalMux I__4504 (
            .O(N__21765),
            .I(\uart_drone.un1_state_2_0 ));
    InMux I__4503 (
            .O(N__21760),
            .I(N__21757));
    LocalMux I__4502 (
            .O(N__21757),
            .I(N__21751));
    InMux I__4501 (
            .O(N__21756),
            .I(N__21743));
    InMux I__4500 (
            .O(N__21755),
            .I(N__21733));
    InMux I__4499 (
            .O(N__21754),
            .I(N__21733));
    Span4Mux_v I__4498 (
            .O(N__21751),
            .I(N__21730));
    InMux I__4497 (
            .O(N__21750),
            .I(N__21727));
    IoInMux I__4496 (
            .O(N__21749),
            .I(N__21724));
    InMux I__4495 (
            .O(N__21748),
            .I(N__21721));
    InMux I__4494 (
            .O(N__21747),
            .I(N__21716));
    InMux I__4493 (
            .O(N__21746),
            .I(N__21716));
    LocalMux I__4492 (
            .O(N__21743),
            .I(N__21713));
    InMux I__4491 (
            .O(N__21742),
            .I(N__21706));
    InMux I__4490 (
            .O(N__21741),
            .I(N__21706));
    InMux I__4489 (
            .O(N__21740),
            .I(N__21706));
    InMux I__4488 (
            .O(N__21739),
            .I(N__21701));
    InMux I__4487 (
            .O(N__21738),
            .I(N__21701));
    LocalMux I__4486 (
            .O(N__21733),
            .I(N__21694));
    Span4Mux_h I__4485 (
            .O(N__21730),
            .I(N__21694));
    LocalMux I__4484 (
            .O(N__21727),
            .I(N__21694));
    LocalMux I__4483 (
            .O(N__21724),
            .I(N__21691));
    LocalMux I__4482 (
            .O(N__21721),
            .I(N__21686));
    LocalMux I__4481 (
            .O(N__21716),
            .I(N__21686));
    Span4Mux_h I__4480 (
            .O(N__21713),
            .I(N__21683));
    LocalMux I__4479 (
            .O(N__21706),
            .I(N__21676));
    LocalMux I__4478 (
            .O(N__21701),
            .I(N__21676));
    Sp12to4 I__4477 (
            .O(N__21694),
            .I(N__21676));
    Span4Mux_s1_v I__4476 (
            .O(N__21691),
            .I(N__21673));
    Span12Mux_v I__4475 (
            .O(N__21686),
            .I(N__21668));
    Sp12to4 I__4474 (
            .O(N__21683),
            .I(N__21668));
    Span12Mux_v I__4473 (
            .O(N__21676),
            .I(N__21665));
    Sp12to4 I__4472 (
            .O(N__21673),
            .I(N__21660));
    Span12Mux_v I__4471 (
            .O(N__21668),
            .I(N__21660));
    Odrv12 I__4470 (
            .O(N__21665),
            .I(uart_drone_input_debug_c));
    Odrv12 I__4469 (
            .O(N__21660),
            .I(uart_drone_input_debug_c));
    InMux I__4468 (
            .O(N__21655),
            .I(N__21651));
    CascadeMux I__4467 (
            .O(N__21654),
            .I(N__21648));
    LocalMux I__4466 (
            .O(N__21651),
            .I(N__21645));
    InMux I__4465 (
            .O(N__21648),
            .I(N__21642));
    Odrv12 I__4464 (
            .O(N__21645),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__4463 (
            .O(N__21642),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    InMux I__4462 (
            .O(N__21637),
            .I(N__21634));
    LocalMux I__4461 (
            .O(N__21634),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__4460 (
            .O(N__21631),
            .I(N__21626));
    CascadeMux I__4459 (
            .O(N__21630),
            .I(N__21623));
    CascadeMux I__4458 (
            .O(N__21629),
            .I(N__21620));
    LocalMux I__4457 (
            .O(N__21626),
            .I(N__21616));
    InMux I__4456 (
            .O(N__21623),
            .I(N__21611));
    InMux I__4455 (
            .O(N__21620),
            .I(N__21611));
    InMux I__4454 (
            .O(N__21619),
            .I(N__21608));
    Span4Mux_h I__4453 (
            .O(N__21616),
            .I(N__21603));
    LocalMux I__4452 (
            .O(N__21611),
            .I(N__21603));
    LocalMux I__4451 (
            .O(N__21608),
            .I(\uart_drone.stateZ0Z_2 ));
    Odrv4 I__4450 (
            .O(N__21603),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__4449 (
            .O(N__21598),
            .I(N__21595));
    InMux I__4448 (
            .O(N__21595),
            .I(N__21592));
    LocalMux I__4447 (
            .O(N__21592),
            .I(N__21589));
    Odrv4 I__4446 (
            .O(N__21589),
            .I(\uart_drone.N_145 ));
    SRMux I__4445 (
            .O(N__21586),
            .I(N__21583));
    LocalMux I__4444 (
            .O(N__21583),
            .I(N__21580));
    Span4Mux_h I__4443 (
            .O(N__21580),
            .I(N__21577));
    Span4Mux_h I__4442 (
            .O(N__21577),
            .I(N__21573));
    SRMux I__4441 (
            .O(N__21576),
            .I(N__21570));
    Odrv4 I__4440 (
            .O(N__21573),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    LocalMux I__4439 (
            .O(N__21570),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__4438 (
            .O(N__21565),
            .I(N__21561));
    CascadeMux I__4437 (
            .O(N__21564),
            .I(N__21558));
    LocalMux I__4436 (
            .O(N__21561),
            .I(N__21554));
    InMux I__4435 (
            .O(N__21558),
            .I(N__21547));
    InMux I__4434 (
            .O(N__21557),
            .I(N__21547));
    Span4Mux_h I__4433 (
            .O(N__21554),
            .I(N__21544));
    InMux I__4432 (
            .O(N__21553),
            .I(N__21539));
    InMux I__4431 (
            .O(N__21552),
            .I(N__21539));
    LocalMux I__4430 (
            .O(N__21547),
            .I(\uart_drone.N_143 ));
    Odrv4 I__4429 (
            .O(N__21544),
            .I(\uart_drone.N_143 ));
    LocalMux I__4428 (
            .O(N__21539),
            .I(\uart_drone.N_143 ));
    InMux I__4427 (
            .O(N__21532),
            .I(N__21526));
    InMux I__4426 (
            .O(N__21531),
            .I(N__21526));
    LocalMux I__4425 (
            .O(N__21526),
            .I(N__21523));
    Odrv4 I__4424 (
            .O(N__21523),
            .I(\uart_drone.N_144_1 ));
    InMux I__4423 (
            .O(N__21520),
            .I(N__21517));
    LocalMux I__4422 (
            .O(N__21517),
            .I(N__21514));
    Odrv4 I__4421 (
            .O(N__21514),
            .I(\scaler_2.N_521_i_l_ofxZ0 ));
    InMux I__4420 (
            .O(N__21511),
            .I(bfn_8_14_0_));
    InMux I__4419 (
            .O(N__21508),
            .I(\scaler_2.un3_source_data_0_cry_8 ));
    InMux I__4418 (
            .O(N__21505),
            .I(N__21501));
    CascadeMux I__4417 (
            .O(N__21504),
            .I(N__21498));
    LocalMux I__4416 (
            .O(N__21501),
            .I(N__21495));
    InMux I__4415 (
            .O(N__21498),
            .I(N__21492));
    Odrv12 I__4414 (
            .O(N__21495),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__4413 (
            .O(N__21492),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    InMux I__4412 (
            .O(N__21487),
            .I(N__21484));
    LocalMux I__4411 (
            .O(N__21484),
            .I(N__21480));
    CascadeMux I__4410 (
            .O(N__21483),
            .I(N__21477));
    Span4Mux_h I__4409 (
            .O(N__21480),
            .I(N__21474));
    InMux I__4408 (
            .O(N__21477),
            .I(N__21471));
    Odrv4 I__4407 (
            .O(N__21474),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__4406 (
            .O(N__21471),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    InMux I__4405 (
            .O(N__21466),
            .I(N__21463));
    LocalMux I__4404 (
            .O(N__21463),
            .I(N__21460));
    Odrv4 I__4403 (
            .O(N__21460),
            .I(frame_decoder_CH2data_1));
    InMux I__4402 (
            .O(N__21457),
            .I(\scaler_2.un3_source_data_0_cry_0 ));
    InMux I__4401 (
            .O(N__21454),
            .I(N__21451));
    LocalMux I__4400 (
            .O(N__21451),
            .I(frame_decoder_CH2data_2));
    InMux I__4399 (
            .O(N__21448),
            .I(\scaler_2.un3_source_data_0_cry_1 ));
    InMux I__4398 (
            .O(N__21445),
            .I(N__21442));
    LocalMux I__4397 (
            .O(N__21442),
            .I(frame_decoder_CH2data_3));
    CascadeMux I__4396 (
            .O(N__21439),
            .I(N__21436));
    InMux I__4395 (
            .O(N__21436),
            .I(N__21433));
    LocalMux I__4394 (
            .O(N__21433),
            .I(frame_decoder_OFF2data_3));
    InMux I__4393 (
            .O(N__21430),
            .I(\scaler_2.un3_source_data_0_cry_2 ));
    InMux I__4392 (
            .O(N__21427),
            .I(N__21424));
    LocalMux I__4391 (
            .O(N__21424),
            .I(N__21421));
    Odrv4 I__4390 (
            .O(N__21421),
            .I(frame_decoder_CH2data_4));
    InMux I__4389 (
            .O(N__21418),
            .I(\scaler_2.un3_source_data_0_cry_3 ));
    InMux I__4388 (
            .O(N__21415),
            .I(N__21412));
    LocalMux I__4387 (
            .O(N__21412),
            .I(frame_decoder_CH2data_5));
    CascadeMux I__4386 (
            .O(N__21409),
            .I(N__21406));
    InMux I__4385 (
            .O(N__21406),
            .I(N__21403));
    LocalMux I__4384 (
            .O(N__21403),
            .I(frame_decoder_OFF2data_5));
    InMux I__4383 (
            .O(N__21400),
            .I(\scaler_2.un3_source_data_0_cry_4 ));
    InMux I__4382 (
            .O(N__21397),
            .I(N__21394));
    LocalMux I__4381 (
            .O(N__21394),
            .I(frame_decoder_CH2data_6));
    CascadeMux I__4380 (
            .O(N__21391),
            .I(N__21388));
    InMux I__4379 (
            .O(N__21388),
            .I(N__21385));
    LocalMux I__4378 (
            .O(N__21385),
            .I(N__21382));
    Odrv4 I__4377 (
            .O(N__21382),
            .I(frame_decoder_OFF2data_6));
    InMux I__4376 (
            .O(N__21379),
            .I(\scaler_2.un3_source_data_0_cry_5 ));
    InMux I__4375 (
            .O(N__21376),
            .I(N__21373));
    LocalMux I__4374 (
            .O(N__21373),
            .I(N__21370));
    Odrv4 I__4373 (
            .O(N__21370),
            .I(\scaler_2.un3_source_data_0_axb_7 ));
    InMux I__4372 (
            .O(N__21367),
            .I(\scaler_2.un3_source_data_0_cry_6 ));
    InMux I__4371 (
            .O(N__21364),
            .I(N__21361));
    LocalMux I__4370 (
            .O(N__21361),
            .I(\uart_drone_sync.aux_0__0_Z0Z_0 ));
    InMux I__4369 (
            .O(N__21358),
            .I(N__21355));
    LocalMux I__4368 (
            .O(N__21355),
            .I(\uart_drone_sync.aux_1__0_Z0Z_0 ));
    InMux I__4367 (
            .O(N__21352),
            .I(N__21349));
    LocalMux I__4366 (
            .O(N__21349),
            .I(\uart_drone_sync.aux_2__0_Z0Z_0 ));
    InMux I__4365 (
            .O(N__21346),
            .I(N__21343));
    LocalMux I__4364 (
            .O(N__21343),
            .I(\uart_drone_sync.aux_3__0_Z0Z_0 ));
    CEMux I__4363 (
            .O(N__21340),
            .I(N__21335));
    CEMux I__4362 (
            .O(N__21339),
            .I(N__21332));
    CEMux I__4361 (
            .O(N__21338),
            .I(N__21329));
    LocalMux I__4360 (
            .O(N__21335),
            .I(N__21326));
    LocalMux I__4359 (
            .O(N__21332),
            .I(N__21321));
    LocalMux I__4358 (
            .O(N__21329),
            .I(N__21321));
    Span4Mux_h I__4357 (
            .O(N__21326),
            .I(N__21318));
    Span4Mux_v I__4356 (
            .O(N__21321),
            .I(N__21315));
    Odrv4 I__4355 (
            .O(N__21318),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    Odrv4 I__4354 (
            .O(N__21315),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__4353 (
            .O(N__21310),
            .I(N__21304));
    InMux I__4352 (
            .O(N__21309),
            .I(N__21304));
    LocalMux I__4351 (
            .O(N__21304),
            .I(frame_decoder_CH2data_7));
    CascadeMux I__4350 (
            .O(N__21301),
            .I(N__21298));
    InMux I__4349 (
            .O(N__21298),
            .I(N__21291));
    InMux I__4348 (
            .O(N__21297),
            .I(N__21291));
    InMux I__4347 (
            .O(N__21296),
            .I(N__21288));
    LocalMux I__4346 (
            .O(N__21291),
            .I(N__21285));
    LocalMux I__4345 (
            .O(N__21288),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv12 I__4344 (
            .O(N__21285),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__4343 (
            .O(N__21280),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__4342 (
            .O(N__21277),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__4341 (
            .O(N__21274),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__4340 (
            .O(N__21271),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__4339 (
            .O(N__21268),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__4338 (
            .O(N__21265),
            .I(bfn_7_30_0_));
    InMux I__4337 (
            .O(N__21262),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__4336 (
            .O(N__21259),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__4335 (
            .O(N__21256),
            .I(N__21247));
    SRMux I__4334 (
            .O(N__21255),
            .I(N__21247));
    SRMux I__4333 (
            .O(N__21254),
            .I(N__21247));
    GlobalMux I__4332 (
            .O(N__21247),
            .I(N__21244));
    gio2CtrlBuf I__4331 (
            .O(N__21244),
            .I(\ppm_encoder_1.N_168_g ));
    InMux I__4330 (
            .O(N__21241),
            .I(N__21238));
    LocalMux I__4329 (
            .O(N__21238),
            .I(uart_input_drone_c));
    InMux I__4328 (
            .O(N__21235),
            .I(N__21232));
    LocalMux I__4327 (
            .O(N__21232),
            .I(N__21226));
    InMux I__4326 (
            .O(N__21231),
            .I(N__21221));
    InMux I__4325 (
            .O(N__21230),
            .I(N__21221));
    InMux I__4324 (
            .O(N__21229),
            .I(N__21218));
    Span4Mux_h I__4323 (
            .O(N__21226),
            .I(N__21215));
    LocalMux I__4322 (
            .O(N__21221),
            .I(N__21212));
    LocalMux I__4321 (
            .O(N__21218),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    Odrv4 I__4320 (
            .O(N__21215),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    Odrv4 I__4319 (
            .O(N__21212),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__4318 (
            .O(N__21205),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    CascadeMux I__4317 (
            .O(N__21202),
            .I(N__21199));
    InMux I__4316 (
            .O(N__21199),
            .I(N__21195));
    CascadeMux I__4315 (
            .O(N__21198),
            .I(N__21192));
    LocalMux I__4314 (
            .O(N__21195),
            .I(N__21187));
    InMux I__4313 (
            .O(N__21192),
            .I(N__21182));
    InMux I__4312 (
            .O(N__21191),
            .I(N__21182));
    InMux I__4311 (
            .O(N__21190),
            .I(N__21179));
    Span4Mux_h I__4310 (
            .O(N__21187),
            .I(N__21176));
    LocalMux I__4309 (
            .O(N__21182),
            .I(N__21173));
    LocalMux I__4308 (
            .O(N__21179),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    Odrv4 I__4307 (
            .O(N__21176),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    Odrv4 I__4306 (
            .O(N__21173),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__4305 (
            .O(N__21166),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__4304 (
            .O(N__21163),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__4303 (
            .O(N__21160),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__4302 (
            .O(N__21157),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__4301 (
            .O(N__21154),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__4300 (
            .O(N__21151),
            .I(bfn_7_29_0_));
    InMux I__4299 (
            .O(N__21148),
            .I(N__21143));
    InMux I__4298 (
            .O(N__21147),
            .I(N__21140));
    InMux I__4297 (
            .O(N__21146),
            .I(N__21137));
    LocalMux I__4296 (
            .O(N__21143),
            .I(N__21132));
    LocalMux I__4295 (
            .O(N__21140),
            .I(N__21132));
    LocalMux I__4294 (
            .O(N__21137),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv12 I__4293 (
            .O(N__21132),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__4292 (
            .O(N__21127),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__4291 (
            .O(N__21124),
            .I(N__21117));
    InMux I__4290 (
            .O(N__21123),
            .I(N__21117));
    InMux I__4289 (
            .O(N__21122),
            .I(N__21114));
    LocalMux I__4288 (
            .O(N__21117),
            .I(N__21111));
    LocalMux I__4287 (
            .O(N__21114),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__4286 (
            .O(N__21111),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__4285 (
            .O(N__21106),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__4284 (
            .O(N__21103),
            .I(N__21099));
    InMux I__4283 (
            .O(N__21102),
            .I(N__21096));
    LocalMux I__4282 (
            .O(N__21099),
            .I(N__21093));
    LocalMux I__4281 (
            .O(N__21096),
            .I(N__21090));
    Span4Mux_v I__4280 (
            .O(N__21093),
            .I(N__21084));
    Span4Mux_v I__4279 (
            .O(N__21090),
            .I(N__21084));
    InMux I__4278 (
            .O(N__21089),
            .I(N__21081));
    Odrv4 I__4277 (
            .O(N__21084),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__4276 (
            .O(N__21081),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    CascadeMux I__4275 (
            .O(N__21076),
            .I(N__21073));
    InMux I__4274 (
            .O(N__21073),
            .I(N__21069));
    InMux I__4273 (
            .O(N__21072),
            .I(N__21066));
    LocalMux I__4272 (
            .O(N__21069),
            .I(N__21062));
    LocalMux I__4271 (
            .O(N__21066),
            .I(N__21059));
    InMux I__4270 (
            .O(N__21065),
            .I(N__21056));
    Span4Mux_h I__4269 (
            .O(N__21062),
            .I(N__21053));
    Span4Mux_h I__4268 (
            .O(N__21059),
            .I(N__21050));
    LocalMux I__4267 (
            .O(N__21056),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__4266 (
            .O(N__21053),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__4265 (
            .O(N__21050),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__4264 (
            .O(N__21043),
            .I(N__21039));
    InMux I__4263 (
            .O(N__21042),
            .I(N__21036));
    LocalMux I__4262 (
            .O(N__21039),
            .I(N__21033));
    LocalMux I__4261 (
            .O(N__21036),
            .I(N__21029));
    Span4Mux_h I__4260 (
            .O(N__21033),
            .I(N__21026));
    InMux I__4259 (
            .O(N__21032),
            .I(N__21023));
    Odrv12 I__4258 (
            .O(N__21029),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__4257 (
            .O(N__21026),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__4256 (
            .O(N__21023),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__4255 (
            .O(N__21016),
            .I(N__21011));
    CascadeMux I__4254 (
            .O(N__21015),
            .I(N__21008));
    InMux I__4253 (
            .O(N__21014),
            .I(N__21005));
    LocalMux I__4252 (
            .O(N__21011),
            .I(N__21002));
    InMux I__4251 (
            .O(N__21008),
            .I(N__20999));
    LocalMux I__4250 (
            .O(N__21005),
            .I(N__20996));
    Span4Mux_s3_h I__4249 (
            .O(N__21002),
            .I(N__20993));
    LocalMux I__4248 (
            .O(N__20999),
            .I(N__20990));
    Span4Mux_v I__4247 (
            .O(N__20996),
            .I(N__20985));
    Span4Mux_h I__4246 (
            .O(N__20993),
            .I(N__20985));
    Odrv4 I__4245 (
            .O(N__20990),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__4244 (
            .O(N__20985),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    CascadeMux I__4243 (
            .O(N__20980),
            .I(N__20976));
    CascadeMux I__4242 (
            .O(N__20979),
            .I(N__20973));
    InMux I__4241 (
            .O(N__20976),
            .I(N__20969));
    InMux I__4240 (
            .O(N__20973),
            .I(N__20966));
    CascadeMux I__4239 (
            .O(N__20972),
            .I(N__20963));
    LocalMux I__4238 (
            .O(N__20969),
            .I(N__20952));
    LocalMux I__4237 (
            .O(N__20966),
            .I(N__20952));
    InMux I__4236 (
            .O(N__20963),
            .I(N__20949));
    InMux I__4235 (
            .O(N__20962),
            .I(N__20944));
    InMux I__4234 (
            .O(N__20961),
            .I(N__20939));
    InMux I__4233 (
            .O(N__20960),
            .I(N__20939));
    InMux I__4232 (
            .O(N__20959),
            .I(N__20935));
    InMux I__4231 (
            .O(N__20958),
            .I(N__20928));
    InMux I__4230 (
            .O(N__20957),
            .I(N__20925));
    Span4Mux_v I__4229 (
            .O(N__20952),
            .I(N__20915));
    LocalMux I__4228 (
            .O(N__20949),
            .I(N__20915));
    InMux I__4227 (
            .O(N__20948),
            .I(N__20912));
    InMux I__4226 (
            .O(N__20947),
            .I(N__20909));
    LocalMux I__4225 (
            .O(N__20944),
            .I(N__20904));
    LocalMux I__4224 (
            .O(N__20939),
            .I(N__20904));
    InMux I__4223 (
            .O(N__20938),
            .I(N__20901));
    LocalMux I__4222 (
            .O(N__20935),
            .I(N__20898));
    InMux I__4221 (
            .O(N__20934),
            .I(N__20895));
    InMux I__4220 (
            .O(N__20933),
            .I(N__20892));
    InMux I__4219 (
            .O(N__20932),
            .I(N__20889));
    CascadeMux I__4218 (
            .O(N__20931),
            .I(N__20886));
    LocalMux I__4217 (
            .O(N__20928),
            .I(N__20882));
    LocalMux I__4216 (
            .O(N__20925),
            .I(N__20879));
    InMux I__4215 (
            .O(N__20924),
            .I(N__20872));
    InMux I__4214 (
            .O(N__20923),
            .I(N__20872));
    InMux I__4213 (
            .O(N__20922),
            .I(N__20872));
    InMux I__4212 (
            .O(N__20921),
            .I(N__20869));
    InMux I__4211 (
            .O(N__20920),
            .I(N__20866));
    Span4Mux_h I__4210 (
            .O(N__20915),
            .I(N__20861));
    LocalMux I__4209 (
            .O(N__20912),
            .I(N__20861));
    LocalMux I__4208 (
            .O(N__20909),
            .I(N__20856));
    Span4Mux_v I__4207 (
            .O(N__20904),
            .I(N__20856));
    LocalMux I__4206 (
            .O(N__20901),
            .I(N__20849));
    Span4Mux_h I__4205 (
            .O(N__20898),
            .I(N__20849));
    LocalMux I__4204 (
            .O(N__20895),
            .I(N__20849));
    LocalMux I__4203 (
            .O(N__20892),
            .I(N__20844));
    LocalMux I__4202 (
            .O(N__20889),
            .I(N__20844));
    InMux I__4201 (
            .O(N__20886),
            .I(N__20839));
    InMux I__4200 (
            .O(N__20885),
            .I(N__20839));
    Span12Mux_v I__4199 (
            .O(N__20882),
            .I(N__20828));
    Span12Mux_s3_v I__4198 (
            .O(N__20879),
            .I(N__20828));
    LocalMux I__4197 (
            .O(N__20872),
            .I(N__20828));
    LocalMux I__4196 (
            .O(N__20869),
            .I(N__20828));
    LocalMux I__4195 (
            .O(N__20866),
            .I(N__20828));
    Span4Mux_v I__4194 (
            .O(N__20861),
            .I(N__20825));
    Span4Mux_h I__4193 (
            .O(N__20856),
            .I(N__20820));
    Span4Mux_v I__4192 (
            .O(N__20849),
            .I(N__20820));
    Odrv4 I__4191 (
            .O(N__20844),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__4190 (
            .O(N__20839),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv12 I__4189 (
            .O(N__20828),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__4188 (
            .O(N__20825),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__4187 (
            .O(N__20820),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    CascadeMux I__4186 (
            .O(N__20809),
            .I(N__20803));
    InMux I__4185 (
            .O(N__20808),
            .I(N__20800));
    CascadeMux I__4184 (
            .O(N__20807),
            .I(N__20794));
    CascadeMux I__4183 (
            .O(N__20806),
            .I(N__20787));
    InMux I__4182 (
            .O(N__20803),
            .I(N__20770));
    LocalMux I__4181 (
            .O(N__20800),
            .I(N__20767));
    InMux I__4180 (
            .O(N__20799),
            .I(N__20760));
    InMux I__4179 (
            .O(N__20798),
            .I(N__20760));
    InMux I__4178 (
            .O(N__20797),
            .I(N__20760));
    InMux I__4177 (
            .O(N__20794),
            .I(N__20756));
    InMux I__4176 (
            .O(N__20793),
            .I(N__20747));
    InMux I__4175 (
            .O(N__20792),
            .I(N__20747));
    InMux I__4174 (
            .O(N__20791),
            .I(N__20747));
    InMux I__4173 (
            .O(N__20790),
            .I(N__20747));
    InMux I__4172 (
            .O(N__20787),
            .I(N__20738));
    InMux I__4171 (
            .O(N__20786),
            .I(N__20738));
    InMux I__4170 (
            .O(N__20785),
            .I(N__20738));
    InMux I__4169 (
            .O(N__20784),
            .I(N__20738));
    InMux I__4168 (
            .O(N__20783),
            .I(N__20731));
    InMux I__4167 (
            .O(N__20782),
            .I(N__20731));
    InMux I__4166 (
            .O(N__20781),
            .I(N__20731));
    InMux I__4165 (
            .O(N__20780),
            .I(N__20722));
    InMux I__4164 (
            .O(N__20779),
            .I(N__20722));
    InMux I__4163 (
            .O(N__20778),
            .I(N__20722));
    InMux I__4162 (
            .O(N__20777),
            .I(N__20722));
    InMux I__4161 (
            .O(N__20776),
            .I(N__20715));
    InMux I__4160 (
            .O(N__20775),
            .I(N__20715));
    InMux I__4159 (
            .O(N__20774),
            .I(N__20715));
    InMux I__4158 (
            .O(N__20773),
            .I(N__20710));
    LocalMux I__4157 (
            .O(N__20770),
            .I(N__20703));
    Span4Mux_h I__4156 (
            .O(N__20767),
            .I(N__20703));
    LocalMux I__4155 (
            .O(N__20760),
            .I(N__20703));
    InMux I__4154 (
            .O(N__20759),
            .I(N__20699));
    LocalMux I__4153 (
            .O(N__20756),
            .I(N__20694));
    LocalMux I__4152 (
            .O(N__20747),
            .I(N__20694));
    LocalMux I__4151 (
            .O(N__20738),
            .I(N__20682));
    LocalMux I__4150 (
            .O(N__20731),
            .I(N__20679));
    LocalMux I__4149 (
            .O(N__20722),
            .I(N__20676));
    LocalMux I__4148 (
            .O(N__20715),
            .I(N__20673));
    InMux I__4147 (
            .O(N__20714),
            .I(N__20668));
    InMux I__4146 (
            .O(N__20713),
            .I(N__20668));
    LocalMux I__4145 (
            .O(N__20710),
            .I(N__20663));
    Span4Mux_h I__4144 (
            .O(N__20703),
            .I(N__20660));
    InMux I__4143 (
            .O(N__20702),
            .I(N__20657));
    LocalMux I__4142 (
            .O(N__20699),
            .I(N__20652));
    Span4Mux_s2_v I__4141 (
            .O(N__20694),
            .I(N__20652));
    InMux I__4140 (
            .O(N__20693),
            .I(N__20641));
    InMux I__4139 (
            .O(N__20692),
            .I(N__20641));
    InMux I__4138 (
            .O(N__20691),
            .I(N__20641));
    InMux I__4137 (
            .O(N__20690),
            .I(N__20641));
    InMux I__4136 (
            .O(N__20689),
            .I(N__20641));
    InMux I__4135 (
            .O(N__20688),
            .I(N__20638));
    InMux I__4134 (
            .O(N__20687),
            .I(N__20635));
    InMux I__4133 (
            .O(N__20686),
            .I(N__20630));
    InMux I__4132 (
            .O(N__20685),
            .I(N__20630));
    Span4Mux_v I__4131 (
            .O(N__20682),
            .I(N__20619));
    Span4Mux_v I__4130 (
            .O(N__20679),
            .I(N__20619));
    Span4Mux_h I__4129 (
            .O(N__20676),
            .I(N__20619));
    Span4Mux_v I__4128 (
            .O(N__20673),
            .I(N__20619));
    LocalMux I__4127 (
            .O(N__20668),
            .I(N__20619));
    InMux I__4126 (
            .O(N__20667),
            .I(N__20614));
    InMux I__4125 (
            .O(N__20666),
            .I(N__20614));
    Odrv12 I__4124 (
            .O(N__20663),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__4123 (
            .O(N__20660),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4122 (
            .O(N__20657),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__4121 (
            .O(N__20652),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4120 (
            .O(N__20641),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4119 (
            .O(N__20638),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4118 (
            .O(N__20635),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4117 (
            .O(N__20630),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__4116 (
            .O(N__20619),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4115 (
            .O(N__20614),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    CascadeMux I__4114 (
            .O(N__20593),
            .I(N__20590));
    InMux I__4113 (
            .O(N__20590),
            .I(N__20587));
    LocalMux I__4112 (
            .O(N__20587),
            .I(N__20584));
    Span4Mux_s3_h I__4111 (
            .O(N__20584),
            .I(N__20581));
    Span4Mux_h I__4110 (
            .O(N__20581),
            .I(N__20578));
    Odrv4 I__4109 (
            .O(N__20578),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    CascadeMux I__4108 (
            .O(N__20575),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ));
    CascadeMux I__4107 (
            .O(N__20572),
            .I(N__20565));
    InMux I__4106 (
            .O(N__20571),
            .I(N__20560));
    InMux I__4105 (
            .O(N__20570),
            .I(N__20560));
    InMux I__4104 (
            .O(N__20569),
            .I(N__20556));
    InMux I__4103 (
            .O(N__20568),
            .I(N__20546));
    InMux I__4102 (
            .O(N__20565),
            .I(N__20546));
    LocalMux I__4101 (
            .O(N__20560),
            .I(N__20541));
    InMux I__4100 (
            .O(N__20559),
            .I(N__20538));
    LocalMux I__4099 (
            .O(N__20556),
            .I(N__20534));
    InMux I__4098 (
            .O(N__20555),
            .I(N__20531));
    InMux I__4097 (
            .O(N__20554),
            .I(N__20528));
    InMux I__4096 (
            .O(N__20553),
            .I(N__20521));
    InMux I__4095 (
            .O(N__20552),
            .I(N__20521));
    InMux I__4094 (
            .O(N__20551),
            .I(N__20521));
    LocalMux I__4093 (
            .O(N__20546),
            .I(N__20518));
    CascadeMux I__4092 (
            .O(N__20545),
            .I(N__20510));
    InMux I__4091 (
            .O(N__20544),
            .I(N__20507));
    Span4Mux_s2_v I__4090 (
            .O(N__20541),
            .I(N__20504));
    LocalMux I__4089 (
            .O(N__20538),
            .I(N__20501));
    InMux I__4088 (
            .O(N__20537),
            .I(N__20498));
    Span4Mux_v I__4087 (
            .O(N__20534),
            .I(N__20491));
    LocalMux I__4086 (
            .O(N__20531),
            .I(N__20491));
    LocalMux I__4085 (
            .O(N__20528),
            .I(N__20491));
    LocalMux I__4084 (
            .O(N__20521),
            .I(N__20486));
    Span4Mux_h I__4083 (
            .O(N__20518),
            .I(N__20486));
    InMux I__4082 (
            .O(N__20517),
            .I(N__20483));
    InMux I__4081 (
            .O(N__20516),
            .I(N__20478));
    InMux I__4080 (
            .O(N__20515),
            .I(N__20478));
    InMux I__4079 (
            .O(N__20514),
            .I(N__20475));
    InMux I__4078 (
            .O(N__20513),
            .I(N__20470));
    InMux I__4077 (
            .O(N__20510),
            .I(N__20470));
    LocalMux I__4076 (
            .O(N__20507),
            .I(N__20467));
    Span4Mux_h I__4075 (
            .O(N__20504),
            .I(N__20462));
    Span4Mux_h I__4074 (
            .O(N__20501),
            .I(N__20462));
    LocalMux I__4073 (
            .O(N__20498),
            .I(N__20455));
    Span4Mux_h I__4072 (
            .O(N__20491),
            .I(N__20455));
    Span4Mux_v I__4071 (
            .O(N__20486),
            .I(N__20455));
    LocalMux I__4070 (
            .O(N__20483),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__4069 (
            .O(N__20478),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__4068 (
            .O(N__20475),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__4067 (
            .O(N__20470),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__4066 (
            .O(N__20467),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__4065 (
            .O(N__20462),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__4064 (
            .O(N__20455),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__4063 (
            .O(N__20440),
            .I(N__20435));
    InMux I__4062 (
            .O(N__20439),
            .I(N__20430));
    InMux I__4061 (
            .O(N__20438),
            .I(N__20430));
    LocalMux I__4060 (
            .O(N__20435),
            .I(N__20427));
    LocalMux I__4059 (
            .O(N__20430),
            .I(N__20424));
    Span4Mux_h I__4058 (
            .O(N__20427),
            .I(N__20419));
    Span4Mux_h I__4057 (
            .O(N__20424),
            .I(N__20419));
    Odrv4 I__4056 (
            .O(N__20419),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    CascadeMux I__4055 (
            .O(N__20416),
            .I(N__20413));
    InMux I__4054 (
            .O(N__20413),
            .I(N__20409));
    CascadeMux I__4053 (
            .O(N__20412),
            .I(N__20405));
    LocalMux I__4052 (
            .O(N__20409),
            .I(N__20402));
    InMux I__4051 (
            .O(N__20408),
            .I(N__20399));
    InMux I__4050 (
            .O(N__20405),
            .I(N__20396));
    Span4Mux_v I__4049 (
            .O(N__20402),
            .I(N__20393));
    LocalMux I__4048 (
            .O(N__20399),
            .I(N__20390));
    LocalMux I__4047 (
            .O(N__20396),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__4046 (
            .O(N__20393),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv12 I__4045 (
            .O(N__20390),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    CascadeMux I__4044 (
            .O(N__20383),
            .I(N__20376));
    CascadeMux I__4043 (
            .O(N__20382),
            .I(N__20373));
    CascadeMux I__4042 (
            .O(N__20381),
            .I(N__20370));
    CascadeMux I__4041 (
            .O(N__20380),
            .I(N__20366));
    CascadeMux I__4040 (
            .O(N__20379),
            .I(N__20362));
    InMux I__4039 (
            .O(N__20376),
            .I(N__20355));
    InMux I__4038 (
            .O(N__20373),
            .I(N__20355));
    InMux I__4037 (
            .O(N__20370),
            .I(N__20352));
    InMux I__4036 (
            .O(N__20369),
            .I(N__20346));
    InMux I__4035 (
            .O(N__20366),
            .I(N__20346));
    InMux I__4034 (
            .O(N__20365),
            .I(N__20340));
    InMux I__4033 (
            .O(N__20362),
            .I(N__20340));
    InMux I__4032 (
            .O(N__20361),
            .I(N__20337));
    InMux I__4031 (
            .O(N__20360),
            .I(N__20334));
    LocalMux I__4030 (
            .O(N__20355),
            .I(N__20331));
    LocalMux I__4029 (
            .O(N__20352),
            .I(N__20328));
    CascadeMux I__4028 (
            .O(N__20351),
            .I(N__20324));
    LocalMux I__4027 (
            .O(N__20346),
            .I(N__20318));
    InMux I__4026 (
            .O(N__20345),
            .I(N__20315));
    LocalMux I__4025 (
            .O(N__20340),
            .I(N__20312));
    LocalMux I__4024 (
            .O(N__20337),
            .I(N__20309));
    LocalMux I__4023 (
            .O(N__20334),
            .I(N__20302));
    Span4Mux_s3_v I__4022 (
            .O(N__20331),
            .I(N__20302));
    Span4Mux_s2_h I__4021 (
            .O(N__20328),
            .I(N__20302));
    InMux I__4020 (
            .O(N__20327),
            .I(N__20293));
    InMux I__4019 (
            .O(N__20324),
            .I(N__20293));
    InMux I__4018 (
            .O(N__20323),
            .I(N__20293));
    InMux I__4017 (
            .O(N__20322),
            .I(N__20293));
    InMux I__4016 (
            .O(N__20321),
            .I(N__20290));
    Span4Mux_v I__4015 (
            .O(N__20318),
            .I(N__20285));
    LocalMux I__4014 (
            .O(N__20315),
            .I(N__20285));
    Span4Mux_h I__4013 (
            .O(N__20312),
            .I(N__20282));
    Span4Mux_h I__4012 (
            .O(N__20309),
            .I(N__20277));
    Span4Mux_h I__4011 (
            .O(N__20302),
            .I(N__20277));
    LocalMux I__4010 (
            .O(N__20293),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__4009 (
            .O(N__20290),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__4008 (
            .O(N__20285),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__4007 (
            .O(N__20282),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__4006 (
            .O(N__20277),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    InMux I__4005 (
            .O(N__20266),
            .I(N__20262));
    CascadeMux I__4004 (
            .O(N__20265),
            .I(N__20259));
    LocalMux I__4003 (
            .O(N__20262),
            .I(N__20256));
    InMux I__4002 (
            .O(N__20259),
            .I(N__20253));
    Odrv4 I__4001 (
            .O(N__20256),
            .I(\ppm_encoder_1.N_590_i ));
    LocalMux I__4000 (
            .O(N__20253),
            .I(\ppm_encoder_1.N_590_i ));
    InMux I__3999 (
            .O(N__20248),
            .I(N__20245));
    LocalMux I__3998 (
            .O(N__20245),
            .I(N__20240));
    InMux I__3997 (
            .O(N__20244),
            .I(N__20237));
    InMux I__3996 (
            .O(N__20243),
            .I(N__20234));
    Span4Mux_s2_v I__3995 (
            .O(N__20240),
            .I(N__20229));
    LocalMux I__3994 (
            .O(N__20237),
            .I(N__20229));
    LocalMux I__3993 (
            .O(N__20234),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__3992 (
            .O(N__20229),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__3991 (
            .O(N__20224),
            .I(N__20221));
    LocalMux I__3990 (
            .O(N__20221),
            .I(N__20215));
    InMux I__3989 (
            .O(N__20220),
            .I(N__20210));
    InMux I__3988 (
            .O(N__20219),
            .I(N__20210));
    InMux I__3987 (
            .O(N__20218),
            .I(N__20207));
    Span4Mux_h I__3986 (
            .O(N__20215),
            .I(N__20204));
    LocalMux I__3985 (
            .O(N__20210),
            .I(N__20201));
    LocalMux I__3984 (
            .O(N__20207),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__3983 (
            .O(N__20204),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__3982 (
            .O(N__20201),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__3981 (
            .O(N__20194),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__3980 (
            .O(N__20191),
            .I(N__20188));
    LocalMux I__3979 (
            .O(N__20188),
            .I(N__20185));
    Span4Mux_h I__3978 (
            .O(N__20185),
            .I(N__20181));
    InMux I__3977 (
            .O(N__20184),
            .I(N__20178));
    Span4Mux_h I__3976 (
            .O(N__20181),
            .I(N__20173));
    LocalMux I__3975 (
            .O(N__20178),
            .I(N__20173));
    Odrv4 I__3974 (
            .O(N__20173),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__3973 (
            .O(N__20170),
            .I(\ppm_encoder_1.N_305_cascade_ ));
    InMux I__3972 (
            .O(N__20167),
            .I(N__20164));
    LocalMux I__3971 (
            .O(N__20164),
            .I(N__20161));
    Span4Mux_h I__3970 (
            .O(N__20161),
            .I(N__20158));
    Odrv4 I__3969 (
            .O(N__20158),
            .I(\ppm_encoder_1.N_298 ));
    InMux I__3968 (
            .O(N__20155),
            .I(N__20152));
    LocalMux I__3967 (
            .O(N__20152),
            .I(N__20147));
    InMux I__3966 (
            .O(N__20151),
            .I(N__20142));
    InMux I__3965 (
            .O(N__20150),
            .I(N__20142));
    Odrv12 I__3964 (
            .O(N__20147),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    LocalMux I__3963 (
            .O(N__20142),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__3962 (
            .O(N__20137),
            .I(N__20133));
    CascadeMux I__3961 (
            .O(N__20136),
            .I(N__20130));
    LocalMux I__3960 (
            .O(N__20133),
            .I(N__20126));
    InMux I__3959 (
            .O(N__20130),
            .I(N__20123));
    CascadeMux I__3958 (
            .O(N__20129),
            .I(N__20120));
    Span4Mux_v I__3957 (
            .O(N__20126),
            .I(N__20117));
    LocalMux I__3956 (
            .O(N__20123),
            .I(N__20114));
    InMux I__3955 (
            .O(N__20120),
            .I(N__20111));
    Span4Mux_h I__3954 (
            .O(N__20117),
            .I(N__20108));
    Span4Mux_v I__3953 (
            .O(N__20114),
            .I(N__20105));
    LocalMux I__3952 (
            .O(N__20111),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__3951 (
            .O(N__20108),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__3950 (
            .O(N__20105),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    CascadeMux I__3949 (
            .O(N__20098),
            .I(\ppm_encoder_1.N_304_cascade_ ));
    InMux I__3948 (
            .O(N__20095),
            .I(N__20092));
    LocalMux I__3947 (
            .O(N__20092),
            .I(N__20088));
    InMux I__3946 (
            .O(N__20091),
            .I(N__20084));
    Span4Mux_s3_h I__3945 (
            .O(N__20088),
            .I(N__20081));
    InMux I__3944 (
            .O(N__20087),
            .I(N__20078));
    LocalMux I__3943 (
            .O(N__20084),
            .I(N__20073));
    Span4Mux_h I__3942 (
            .O(N__20081),
            .I(N__20073));
    LocalMux I__3941 (
            .O(N__20078),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    Odrv4 I__3940 (
            .O(N__20073),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__3939 (
            .O(N__20068),
            .I(N__20063));
    InMux I__3938 (
            .O(N__20067),
            .I(N__20058));
    InMux I__3937 (
            .O(N__20066),
            .I(N__20058));
    LocalMux I__3936 (
            .O(N__20063),
            .I(N__20055));
    LocalMux I__3935 (
            .O(N__20058),
            .I(N__20052));
    Span4Mux_h I__3934 (
            .O(N__20055),
            .I(N__20049));
    Span4Mux_h I__3933 (
            .O(N__20052),
            .I(N__20046));
    Odrv4 I__3932 (
            .O(N__20049),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    Odrv4 I__3931 (
            .O(N__20046),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__3930 (
            .O(N__20041),
            .I(N__20036));
    InMux I__3929 (
            .O(N__20040),
            .I(N__20033));
    InMux I__3928 (
            .O(N__20039),
            .I(N__20030));
    LocalMux I__3927 (
            .O(N__20036),
            .I(N__20027));
    LocalMux I__3926 (
            .O(N__20033),
            .I(N__20024));
    LocalMux I__3925 (
            .O(N__20030),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__3924 (
            .O(N__20027),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv12 I__3923 (
            .O(N__20024),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__3922 (
            .O(N__20017),
            .I(N__20014));
    InMux I__3921 (
            .O(N__20014),
            .I(N__20011));
    LocalMux I__3920 (
            .O(N__20011),
            .I(N__20006));
    CascadeMux I__3919 (
            .O(N__20010),
            .I(N__20001));
    InMux I__3918 (
            .O(N__20009),
            .I(N__19998));
    Span4Mux_h I__3917 (
            .O(N__20006),
            .I(N__19995));
    InMux I__3916 (
            .O(N__20005),
            .I(N__19988));
    InMux I__3915 (
            .O(N__20004),
            .I(N__19988));
    InMux I__3914 (
            .O(N__20001),
            .I(N__19988));
    LocalMux I__3913 (
            .O(N__19998),
            .I(N__19985));
    Odrv4 I__3912 (
            .O(N__19995),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    LocalMux I__3911 (
            .O(N__19988),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__3910 (
            .O(N__19985),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    CascadeMux I__3909 (
            .O(N__19978),
            .I(\ppm_encoder_1.N_319_cascade_ ));
    InMux I__3908 (
            .O(N__19975),
            .I(N__19972));
    LocalMux I__3907 (
            .O(N__19972),
            .I(N__19969));
    Span4Mux_v I__3906 (
            .O(N__19969),
            .I(N__19966));
    Odrv4 I__3905 (
            .O(N__19966),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    CascadeMux I__3904 (
            .O(N__19963),
            .I(N__19959));
    InMux I__3903 (
            .O(N__19962),
            .I(N__19956));
    InMux I__3902 (
            .O(N__19959),
            .I(N__19953));
    LocalMux I__3901 (
            .O(N__19956),
            .I(N__19949));
    LocalMux I__3900 (
            .O(N__19953),
            .I(N__19946));
    InMux I__3899 (
            .O(N__19952),
            .I(N__19943));
    Span4Mux_v I__3898 (
            .O(N__19949),
            .I(N__19938));
    Span4Mux_h I__3897 (
            .O(N__19946),
            .I(N__19938));
    LocalMux I__3896 (
            .O(N__19943),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__3895 (
            .O(N__19938),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__3894 (
            .O(N__19933),
            .I(N__19930));
    LocalMux I__3893 (
            .O(N__19930),
            .I(N__19927));
    Span4Mux_s3_v I__3892 (
            .O(N__19927),
            .I(N__19924));
    Span4Mux_h I__3891 (
            .O(N__19924),
            .I(N__19921));
    Odrv4 I__3890 (
            .O(N__19921),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__3889 (
            .O(N__19918),
            .I(N__19915));
    LocalMux I__3888 (
            .O(N__19915),
            .I(N__19910));
    InMux I__3887 (
            .O(N__19914),
            .I(N__19905));
    InMux I__3886 (
            .O(N__19913),
            .I(N__19905));
    Odrv4 I__3885 (
            .O(N__19910),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    LocalMux I__3884 (
            .O(N__19905),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__3883 (
            .O(N__19900),
            .I(N__19897));
    LocalMux I__3882 (
            .O(N__19897),
            .I(N__19893));
    InMux I__3881 (
            .O(N__19896),
            .I(N__19890));
    Span4Mux_v I__3880 (
            .O(N__19893),
            .I(N__19887));
    LocalMux I__3879 (
            .O(N__19890),
            .I(N__19884));
    Span4Mux_h I__3878 (
            .O(N__19887),
            .I(N__19881));
    Odrv12 I__3877 (
            .O(N__19884),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv4 I__3876 (
            .O(N__19881),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__3875 (
            .O(N__19876),
            .I(N__19871));
    InMux I__3874 (
            .O(N__19875),
            .I(N__19868));
    CascadeMux I__3873 (
            .O(N__19874),
            .I(N__19865));
    LocalMux I__3872 (
            .O(N__19871),
            .I(N__19862));
    LocalMux I__3871 (
            .O(N__19868),
            .I(N__19859));
    InMux I__3870 (
            .O(N__19865),
            .I(N__19856));
    Span4Mux_v I__3869 (
            .O(N__19862),
            .I(N__19853));
    Span4Mux_h I__3868 (
            .O(N__19859),
            .I(N__19850));
    LocalMux I__3867 (
            .O(N__19856),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__3866 (
            .O(N__19853),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__3865 (
            .O(N__19850),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    InMux I__3864 (
            .O(N__19843),
            .I(N__19840));
    LocalMux I__3863 (
            .O(N__19840),
            .I(N__19837));
    Odrv4 I__3862 (
            .O(N__19837),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__3861 (
            .O(N__19834),
            .I(N__19831));
    LocalMux I__3860 (
            .O(N__19831),
            .I(N__19827));
    CascadeMux I__3859 (
            .O(N__19830),
            .I(N__19824));
    Span4Mux_s3_v I__3858 (
            .O(N__19827),
            .I(N__19821));
    InMux I__3857 (
            .O(N__19824),
            .I(N__19818));
    Span4Mux_v I__3856 (
            .O(N__19821),
            .I(N__19812));
    LocalMux I__3855 (
            .O(N__19818),
            .I(N__19812));
    InMux I__3854 (
            .O(N__19817),
            .I(N__19809));
    Span4Mux_h I__3853 (
            .O(N__19812),
            .I(N__19806));
    LocalMux I__3852 (
            .O(N__19809),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__3851 (
            .O(N__19806),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    InMux I__3850 (
            .O(N__19801),
            .I(N__19798));
    LocalMux I__3849 (
            .O(N__19798),
            .I(N__19793));
    InMux I__3848 (
            .O(N__19797),
            .I(N__19790));
    CascadeMux I__3847 (
            .O(N__19796),
            .I(N__19787));
    Span4Mux_s3_h I__3846 (
            .O(N__19793),
            .I(N__19784));
    LocalMux I__3845 (
            .O(N__19790),
            .I(N__19781));
    InMux I__3844 (
            .O(N__19787),
            .I(N__19778));
    Span4Mux_h I__3843 (
            .O(N__19784),
            .I(N__19775));
    Span4Mux_h I__3842 (
            .O(N__19781),
            .I(N__19772));
    LocalMux I__3841 (
            .O(N__19778),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__3840 (
            .O(N__19775),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__3839 (
            .O(N__19772),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__3838 (
            .O(N__19765),
            .I(N__19762));
    LocalMux I__3837 (
            .O(N__19762),
            .I(N__19759));
    Odrv12 I__3836 (
            .O(N__19759),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__3835 (
            .O(N__19756),
            .I(N__19753));
    LocalMux I__3834 (
            .O(N__19753),
            .I(N__19750));
    Span4Mux_s3_v I__3833 (
            .O(N__19750),
            .I(N__19745));
    InMux I__3832 (
            .O(N__19749),
            .I(N__19742));
    CascadeMux I__3831 (
            .O(N__19748),
            .I(N__19739));
    Span4Mux_h I__3830 (
            .O(N__19745),
            .I(N__19736));
    LocalMux I__3829 (
            .O(N__19742),
            .I(N__19733));
    InMux I__3828 (
            .O(N__19739),
            .I(N__19730));
    Span4Mux_v I__3827 (
            .O(N__19736),
            .I(N__19725));
    Span4Mux_h I__3826 (
            .O(N__19733),
            .I(N__19725));
    LocalMux I__3825 (
            .O(N__19730),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__3824 (
            .O(N__19725),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__3823 (
            .O(N__19720),
            .I(N__19717));
    LocalMux I__3822 (
            .O(N__19717),
            .I(N__19714));
    Odrv4 I__3821 (
            .O(N__19714),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__3820 (
            .O(N__19711),
            .I(N__19704));
    InMux I__3819 (
            .O(N__19710),
            .I(N__19704));
    CascadeMux I__3818 (
            .O(N__19709),
            .I(N__19701));
    LocalMux I__3817 (
            .O(N__19704),
            .I(N__19698));
    InMux I__3816 (
            .O(N__19701),
            .I(N__19695));
    Span4Mux_v I__3815 (
            .O(N__19698),
            .I(N__19692));
    LocalMux I__3814 (
            .O(N__19695),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__3813 (
            .O(N__19692),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__3812 (
            .O(N__19687),
            .I(N__19684));
    LocalMux I__3811 (
            .O(N__19684),
            .I(N__19681));
    Odrv4 I__3810 (
            .O(N__19681),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__3809 (
            .O(N__19678),
            .I(N__19675));
    LocalMux I__3808 (
            .O(N__19675),
            .I(N__19672));
    Odrv4 I__3807 (
            .O(N__19672),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    InMux I__3806 (
            .O(N__19669),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__3805 (
            .O(N__19666),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__3804 (
            .O(N__19663),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__3803 (
            .O(N__19660),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__3802 (
            .O(N__19657),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__3801 (
            .O(N__19654),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__3800 (
            .O(N__19651),
            .I(bfn_7_20_0_));
    InMux I__3799 (
            .O(N__19648),
            .I(N__19645));
    LocalMux I__3798 (
            .O(N__19645),
            .I(N__19642));
    Odrv4 I__3797 (
            .O(N__19642),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__3796 (
            .O(N__19639),
            .I(N__19632));
    InMux I__3795 (
            .O(N__19638),
            .I(N__19632));
    CascadeMux I__3794 (
            .O(N__19637),
            .I(N__19629));
    LocalMux I__3793 (
            .O(N__19632),
            .I(N__19626));
    InMux I__3792 (
            .O(N__19629),
            .I(N__19623));
    Span4Mux_v I__3791 (
            .O(N__19626),
            .I(N__19620));
    LocalMux I__3790 (
            .O(N__19623),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__3789 (
            .O(N__19620),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__3788 (
            .O(N__19615),
            .I(N__19610));
    InMux I__3787 (
            .O(N__19614),
            .I(N__19607));
    CascadeMux I__3786 (
            .O(N__19613),
            .I(N__19604));
    LocalMux I__3785 (
            .O(N__19610),
            .I(N__19599));
    LocalMux I__3784 (
            .O(N__19607),
            .I(N__19599));
    InMux I__3783 (
            .O(N__19604),
            .I(N__19596));
    Span4Mux_v I__3782 (
            .O(N__19599),
            .I(N__19593));
    LocalMux I__3781 (
            .O(N__19596),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    Odrv4 I__3780 (
            .O(N__19593),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    CascadeMux I__3779 (
            .O(N__19588),
            .I(\uart_pc.N_143_cascade_ ));
    SRMux I__3778 (
            .O(N__19585),
            .I(N__19582));
    LocalMux I__3777 (
            .O(N__19582),
            .I(N__19578));
    SRMux I__3776 (
            .O(N__19581),
            .I(N__19575));
    Span4Mux_h I__3775 (
            .O(N__19578),
            .I(N__19572));
    LocalMux I__3774 (
            .O(N__19575),
            .I(N__19569));
    Span4Mux_h I__3773 (
            .O(N__19572),
            .I(N__19566));
    Span12Mux_s7_h I__3772 (
            .O(N__19569),
            .I(N__19563));
    Odrv4 I__3771 (
            .O(N__19566),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv12 I__3770 (
            .O(N__19563),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__3769 (
            .O(N__19558),
            .I(N__19552));
    InMux I__3768 (
            .O(N__19557),
            .I(N__19547));
    InMux I__3767 (
            .O(N__19556),
            .I(N__19547));
    InMux I__3766 (
            .O(N__19555),
            .I(N__19544));
    LocalMux I__3765 (
            .O(N__19552),
            .I(N__19541));
    LocalMux I__3764 (
            .O(N__19547),
            .I(N__19536));
    LocalMux I__3763 (
            .O(N__19544),
            .I(N__19536));
    Span4Mux_h I__3762 (
            .O(N__19541),
            .I(N__19531));
    Span4Mux_v I__3761 (
            .O(N__19536),
            .I(N__19531));
    Odrv4 I__3760 (
            .O(N__19531),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__3759 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__3758 (
            .O(N__19525),
            .I(N__19521));
    InMux I__3757 (
            .O(N__19524),
            .I(N__19518));
    Odrv4 I__3756 (
            .O(N__19521),
            .I(\uart_pc.N_126_li ));
    LocalMux I__3755 (
            .O(N__19518),
            .I(\uart_pc.N_126_li ));
    InMux I__3754 (
            .O(N__19513),
            .I(N__19505));
    InMux I__3753 (
            .O(N__19512),
            .I(N__19496));
    InMux I__3752 (
            .O(N__19511),
            .I(N__19496));
    InMux I__3751 (
            .O(N__19510),
            .I(N__19496));
    InMux I__3750 (
            .O(N__19509),
            .I(N__19496));
    InMux I__3749 (
            .O(N__19508),
            .I(N__19493));
    LocalMux I__3748 (
            .O(N__19505),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__3747 (
            .O(N__19496),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__3746 (
            .O(N__19493),
            .I(\uart_pc.stateZ0Z_4 ));
    InMux I__3745 (
            .O(N__19486),
            .I(N__19483));
    LocalMux I__3744 (
            .O(N__19483),
            .I(N__19479));
    InMux I__3743 (
            .O(N__19482),
            .I(N__19476));
    Span4Mux_v I__3742 (
            .O(N__19479),
            .I(N__19466));
    LocalMux I__3741 (
            .O(N__19476),
            .I(N__19466));
    InMux I__3740 (
            .O(N__19475),
            .I(N__19458));
    InMux I__3739 (
            .O(N__19474),
            .I(N__19458));
    InMux I__3738 (
            .O(N__19473),
            .I(N__19458));
    InMux I__3737 (
            .O(N__19472),
            .I(N__19453));
    InMux I__3736 (
            .O(N__19471),
            .I(N__19453));
    Span4Mux_h I__3735 (
            .O(N__19466),
            .I(N__19450));
    InMux I__3734 (
            .O(N__19465),
            .I(N__19447));
    LocalMux I__3733 (
            .O(N__19458),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__3732 (
            .O(N__19453),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__3731 (
            .O(N__19450),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__3730 (
            .O(N__19447),
            .I(\uart_pc.stateZ0Z_3 ));
    CascadeMux I__3729 (
            .O(N__19438),
            .I(\uart_pc.N_126_li_cascade_ ));
    InMux I__3728 (
            .O(N__19435),
            .I(N__19425));
    InMux I__3727 (
            .O(N__19434),
            .I(N__19410));
    InMux I__3726 (
            .O(N__19433),
            .I(N__19410));
    InMux I__3725 (
            .O(N__19432),
            .I(N__19410));
    InMux I__3724 (
            .O(N__19431),
            .I(N__19410));
    InMux I__3723 (
            .O(N__19430),
            .I(N__19410));
    InMux I__3722 (
            .O(N__19429),
            .I(N__19410));
    InMux I__3721 (
            .O(N__19428),
            .I(N__19410));
    LocalMux I__3720 (
            .O(N__19425),
            .I(N__19407));
    LocalMux I__3719 (
            .O(N__19410),
            .I(N__19404));
    Span4Mux_h I__3718 (
            .O(N__19407),
            .I(N__19401));
    Span4Mux_h I__3717 (
            .O(N__19404),
            .I(N__19398));
    Odrv4 I__3716 (
            .O(N__19401),
            .I(\uart_pc.un1_state_2_0 ));
    Odrv4 I__3715 (
            .O(N__19398),
            .I(\uart_pc.un1_state_2_0 ));
    InMux I__3714 (
            .O(N__19393),
            .I(N__19390));
    LocalMux I__3713 (
            .O(N__19390),
            .I(N__19387));
    Span4Mux_v I__3712 (
            .O(N__19387),
            .I(N__19384));
    Odrv4 I__3711 (
            .O(N__19384),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__3710 (
            .O(N__19381),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__3709 (
            .O(N__19378),
            .I(N__19374));
    InMux I__3708 (
            .O(N__19377),
            .I(N__19371));
    LocalMux I__3707 (
            .O(N__19374),
            .I(N__19367));
    LocalMux I__3706 (
            .O(N__19371),
            .I(N__19364));
    InMux I__3705 (
            .O(N__19370),
            .I(N__19361));
    Span4Mux_v I__3704 (
            .O(N__19367),
            .I(N__19358));
    Span4Mux_h I__3703 (
            .O(N__19364),
            .I(N__19355));
    LocalMux I__3702 (
            .O(N__19361),
            .I(\uart_pc.N_152 ));
    Odrv4 I__3701 (
            .O(N__19358),
            .I(\uart_pc.N_152 ));
    Odrv4 I__3700 (
            .O(N__19355),
            .I(\uart_pc.N_152 ));
    InMux I__3699 (
            .O(N__19348),
            .I(N__19345));
    LocalMux I__3698 (
            .O(N__19345),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__3697 (
            .O(N__19342),
            .I(\uart_pc.N_144_1_cascade_ ));
    InMux I__3696 (
            .O(N__19339),
            .I(N__19335));
    InMux I__3695 (
            .O(N__19338),
            .I(N__19332));
    LocalMux I__3694 (
            .O(N__19335),
            .I(N__19329));
    LocalMux I__3693 (
            .O(N__19332),
            .I(N__19324));
    Span4Mux_h I__3692 (
            .O(N__19329),
            .I(N__19321));
    InMux I__3691 (
            .O(N__19328),
            .I(N__19316));
    InMux I__3690 (
            .O(N__19327),
            .I(N__19316));
    Span4Mux_h I__3689 (
            .O(N__19324),
            .I(N__19313));
    Span4Mux_v I__3688 (
            .O(N__19321),
            .I(N__19310));
    LocalMux I__3687 (
            .O(N__19316),
            .I(N__19307));
    Odrv4 I__3686 (
            .O(N__19313),
            .I(\uart_pc.state_1_sqmuxa ));
    Odrv4 I__3685 (
            .O(N__19310),
            .I(\uart_pc.state_1_sqmuxa ));
    Odrv4 I__3684 (
            .O(N__19307),
            .I(\uart_pc.state_1_sqmuxa ));
    CascadeMux I__3683 (
            .O(N__19300),
            .I(N__19297));
    InMux I__3682 (
            .O(N__19297),
            .I(N__19294));
    LocalMux I__3681 (
            .O(N__19294),
            .I(\uart_pc.N_145 ));
    CascadeMux I__3680 (
            .O(N__19291),
            .I(N__19286));
    InMux I__3679 (
            .O(N__19290),
            .I(N__19279));
    InMux I__3678 (
            .O(N__19289),
            .I(N__19279));
    InMux I__3677 (
            .O(N__19286),
            .I(N__19279));
    LocalMux I__3676 (
            .O(N__19279),
            .I(N__19275));
    CascadeMux I__3675 (
            .O(N__19278),
            .I(N__19271));
    Span4Mux_v I__3674 (
            .O(N__19275),
            .I(N__19268));
    InMux I__3673 (
            .O(N__19274),
            .I(N__19263));
    InMux I__3672 (
            .O(N__19271),
            .I(N__19263));
    Sp12to4 I__3671 (
            .O(N__19268),
            .I(N__19260));
    LocalMux I__3670 (
            .O(N__19263),
            .I(N__19257));
    Odrv12 I__3669 (
            .O(N__19260),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__3668 (
            .O(N__19257),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__3667 (
            .O(N__19252),
            .I(N__19246));
    CascadeMux I__3666 (
            .O(N__19251),
            .I(N__19243));
    InMux I__3665 (
            .O(N__19250),
            .I(N__19240));
    InMux I__3664 (
            .O(N__19249),
            .I(N__19233));
    InMux I__3663 (
            .O(N__19246),
            .I(N__19233));
    InMux I__3662 (
            .O(N__19243),
            .I(N__19233));
    LocalMux I__3661 (
            .O(N__19240),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__3660 (
            .O(N__19233),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__3659 (
            .O(N__19228),
            .I(N__19225));
    LocalMux I__3658 (
            .O(N__19225),
            .I(N__19222));
    Span4Mux_h I__3657 (
            .O(N__19222),
            .I(N__19219));
    Odrv4 I__3656 (
            .O(N__19219),
            .I(\uart_drone.data_Auxce_0_6 ));
    CascadeMux I__3655 (
            .O(N__19216),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__3654 (
            .O(N__19213),
            .I(N__19210));
    InMux I__3653 (
            .O(N__19210),
            .I(N__19206));
    InMux I__3652 (
            .O(N__19209),
            .I(N__19203));
    LocalMux I__3651 (
            .O(N__19206),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__3650 (
            .O(N__19203),
            .I(\uart_pc.stateZ0Z_0 ));
    InMux I__3649 (
            .O(N__19198),
            .I(N__19195));
    LocalMux I__3648 (
            .O(N__19195),
            .I(N__19192));
    Span4Mux_h I__3647 (
            .O(N__19192),
            .I(N__19188));
    InMux I__3646 (
            .O(N__19191),
            .I(N__19185));
    Odrv4 I__3645 (
            .O(N__19188),
            .I(\uart_drone.N_126_li ));
    LocalMux I__3644 (
            .O(N__19185),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__3643 (
            .O(N__19180),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__3642 (
            .O(N__19177),
            .I(N__19173));
    InMux I__3641 (
            .O(N__19176),
            .I(N__19170));
    LocalMux I__3640 (
            .O(N__19173),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__3639 (
            .O(N__19170),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__3638 (
            .O(N__19165),
            .I(N__19162));
    LocalMux I__3637 (
            .O(N__19162),
            .I(N__19159));
    Odrv4 I__3636 (
            .O(N__19159),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__3635 (
            .O(N__19156),
            .I(N__19148));
    CascadeMux I__3634 (
            .O(N__19155),
            .I(N__19145));
    CascadeMux I__3633 (
            .O(N__19154),
            .I(N__19142));
    CascadeMux I__3632 (
            .O(N__19153),
            .I(N__19138));
    CascadeMux I__3631 (
            .O(N__19152),
            .I(N__19134));
    IoInMux I__3630 (
            .O(N__19151),
            .I(N__19129));
    LocalMux I__3629 (
            .O(N__19148),
            .I(N__19126));
    InMux I__3628 (
            .O(N__19145),
            .I(N__19111));
    InMux I__3627 (
            .O(N__19142),
            .I(N__19111));
    InMux I__3626 (
            .O(N__19141),
            .I(N__19111));
    InMux I__3625 (
            .O(N__19138),
            .I(N__19111));
    InMux I__3624 (
            .O(N__19137),
            .I(N__19111));
    InMux I__3623 (
            .O(N__19134),
            .I(N__19111));
    InMux I__3622 (
            .O(N__19133),
            .I(N__19111));
    InMux I__3621 (
            .O(N__19132),
            .I(N__19108));
    LocalMux I__3620 (
            .O(N__19129),
            .I(N__19105));
    Span4Mux_v I__3619 (
            .O(N__19126),
            .I(N__19101));
    LocalMux I__3618 (
            .O(N__19111),
            .I(N__19098));
    LocalMux I__3617 (
            .O(N__19108),
            .I(N__19095));
    IoSpan4Mux I__3616 (
            .O(N__19105),
            .I(N__19089));
    InMux I__3615 (
            .O(N__19104),
            .I(N__19086));
    Sp12to4 I__3614 (
            .O(N__19101),
            .I(N__19083));
    Span4Mux_h I__3613 (
            .O(N__19098),
            .I(N__19080));
    Span4Mux_h I__3612 (
            .O(N__19095),
            .I(N__19077));
    InMux I__3611 (
            .O(N__19094),
            .I(N__19072));
    InMux I__3610 (
            .O(N__19093),
            .I(N__19072));
    InMux I__3609 (
            .O(N__19092),
            .I(N__19069));
    Span4Mux_s1_v I__3608 (
            .O(N__19089),
            .I(N__19066));
    LocalMux I__3607 (
            .O(N__19086),
            .I(N__19055));
    Span12Mux_h I__3606 (
            .O(N__19083),
            .I(N__19055));
    Sp12to4 I__3605 (
            .O(N__19080),
            .I(N__19055));
    Sp12to4 I__3604 (
            .O(N__19077),
            .I(N__19055));
    LocalMux I__3603 (
            .O(N__19072),
            .I(N__19055));
    LocalMux I__3602 (
            .O(N__19069),
            .I(N__19052));
    Span4Mux_h I__3601 (
            .O(N__19066),
            .I(N__19049));
    Span12Mux_v I__3600 (
            .O(N__19055),
            .I(N__19044));
    Span12Mux_s7_h I__3599 (
            .O(N__19052),
            .I(N__19044));
    Odrv4 I__3598 (
            .O(N__19049),
            .I(uart_commands_input_debug_c));
    Odrv12 I__3597 (
            .O(N__19044),
            .I(uart_commands_input_debug_c));
    CascadeMux I__3596 (
            .O(N__19039),
            .I(N__19034));
    InMux I__3595 (
            .O(N__19038),
            .I(N__19031));
    InMux I__3594 (
            .O(N__19037),
            .I(N__19026));
    InMux I__3593 (
            .O(N__19034),
            .I(N__19026));
    LocalMux I__3592 (
            .O(N__19031),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__3591 (
            .O(N__19026),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__3590 (
            .O(N__19021),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    InMux I__3589 (
            .O(N__19018),
            .I(N__19015));
    LocalMux I__3588 (
            .O(N__19015),
            .I(N__19012));
    Odrv4 I__3587 (
            .O(N__19012),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__3586 (
            .O(N__19009),
            .I(N__19006));
    LocalMux I__3585 (
            .O(N__19006),
            .I(N__19003));
    Span4Mux_h I__3584 (
            .O(N__19003),
            .I(N__19000));
    Odrv4 I__3583 (
            .O(N__19000),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__3582 (
            .O(N__18997),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__3581 (
            .O(N__18994),
            .I(N__18989));
    InMux I__3580 (
            .O(N__18993),
            .I(N__18986));
    InMux I__3579 (
            .O(N__18992),
            .I(N__18981));
    InMux I__3578 (
            .O(N__18989),
            .I(N__18981));
    LocalMux I__3577 (
            .O(N__18986),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__3576 (
            .O(N__18981),
            .I(\uart_drone.stateZ0Z_1 ));
    InMux I__3575 (
            .O(N__18976),
            .I(N__18973));
    LocalMux I__3574 (
            .O(N__18973),
            .I(N__18970));
    Span4Mux_v I__3573 (
            .O(N__18970),
            .I(N__18965));
    InMux I__3572 (
            .O(N__18969),
            .I(N__18962));
    InMux I__3571 (
            .O(N__18968),
            .I(N__18959));
    Span4Mux_v I__3570 (
            .O(N__18965),
            .I(N__18955));
    LocalMux I__3569 (
            .O(N__18962),
            .I(N__18950));
    LocalMux I__3568 (
            .O(N__18959),
            .I(N__18950));
    InMux I__3567 (
            .O(N__18958),
            .I(N__18947));
    Odrv4 I__3566 (
            .O(N__18955),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv12 I__3565 (
            .O(N__18950),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__3564 (
            .O(N__18947),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    CascadeMux I__3563 (
            .O(N__18940),
            .I(\ppm_encoder_1.N_237_cascade_ ));
    InMux I__3562 (
            .O(N__18937),
            .I(N__18932));
    InMux I__3561 (
            .O(N__18936),
            .I(N__18929));
    InMux I__3560 (
            .O(N__18935),
            .I(N__18925));
    LocalMux I__3559 (
            .O(N__18932),
            .I(N__18922));
    LocalMux I__3558 (
            .O(N__18929),
            .I(N__18919));
    InMux I__3557 (
            .O(N__18928),
            .I(N__18916));
    LocalMux I__3556 (
            .O(N__18925),
            .I(N__18913));
    Span4Mux_v I__3555 (
            .O(N__18922),
            .I(N__18910));
    Span4Mux_s2_v I__3554 (
            .O(N__18919),
            .I(N__18905));
    LocalMux I__3553 (
            .O(N__18916),
            .I(N__18905));
    Span4Mux_v I__3552 (
            .O(N__18913),
            .I(N__18895));
    Span4Mux_h I__3551 (
            .O(N__18910),
            .I(N__18895));
    Span4Mux_v I__3550 (
            .O(N__18905),
            .I(N__18895));
    InMux I__3549 (
            .O(N__18904),
            .I(N__18888));
    InMux I__3548 (
            .O(N__18903),
            .I(N__18888));
    InMux I__3547 (
            .O(N__18902),
            .I(N__18888));
    Odrv4 I__3546 (
            .O(N__18895),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__3545 (
            .O(N__18888),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    IoInMux I__3544 (
            .O(N__18883),
            .I(N__18880));
    LocalMux I__3543 (
            .O(N__18880),
            .I(N__18877));
    Span4Mux_s1_v I__3542 (
            .O(N__18877),
            .I(N__18874));
    Span4Mux_h I__3541 (
            .O(N__18874),
            .I(N__18871));
    Odrv4 I__3540 (
            .O(N__18871),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__3539 (
            .O(N__18868),
            .I(N__18864));
    InMux I__3538 (
            .O(N__18867),
            .I(N__18861));
    LocalMux I__3537 (
            .O(N__18864),
            .I(N__18858));
    LocalMux I__3536 (
            .O(N__18861),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    Odrv12 I__3535 (
            .O(N__18858),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__3534 (
            .O(N__18853),
            .I(N__18850));
    LocalMux I__3533 (
            .O(N__18850),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__3532 (
            .O(N__18847),
            .I(N__18844));
    LocalMux I__3531 (
            .O(N__18844),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__3530 (
            .O(N__18841),
            .I(N__18838));
    LocalMux I__3529 (
            .O(N__18838),
            .I(\uart_pc_sync.aux_2__0__0_0 ));
    InMux I__3528 (
            .O(N__18835),
            .I(N__18832));
    LocalMux I__3527 (
            .O(N__18832),
            .I(\uart_pc_sync.aux_3__0__0_0 ));
    InMux I__3526 (
            .O(N__18829),
            .I(N__18826));
    LocalMux I__3525 (
            .O(N__18826),
            .I(N__18823));
    Odrv4 I__3524 (
            .O(N__18823),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    InMux I__3523 (
            .O(N__18820),
            .I(N__18817));
    LocalMux I__3522 (
            .O(N__18817),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    CascadeMux I__3521 (
            .O(N__18814),
            .I(N__18811));
    InMux I__3520 (
            .O(N__18811),
            .I(N__18808));
    LocalMux I__3519 (
            .O(N__18808),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    CascadeMux I__3518 (
            .O(N__18805),
            .I(N__18802));
    InMux I__3517 (
            .O(N__18802),
            .I(N__18799));
    LocalMux I__3516 (
            .O(N__18799),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    InMux I__3515 (
            .O(N__18796),
            .I(N__18793));
    LocalMux I__3514 (
            .O(N__18793),
            .I(N__18790));
    Span4Mux_h I__3513 (
            .O(N__18790),
            .I(N__18787));
    Odrv4 I__3512 (
            .O(N__18787),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__3511 (
            .O(N__18784),
            .I(N__18781));
    LocalMux I__3510 (
            .O(N__18781),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__3509 (
            .O(N__18778),
            .I(N__18775));
    LocalMux I__3508 (
            .O(N__18775),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__3507 (
            .O(N__18772),
            .I(N__18769));
    LocalMux I__3506 (
            .O(N__18769),
            .I(N__18766));
    Span4Mux_v I__3505 (
            .O(N__18766),
            .I(N__18763));
    Odrv4 I__3504 (
            .O(N__18763),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    InMux I__3503 (
            .O(N__18760),
            .I(N__18757));
    LocalMux I__3502 (
            .O(N__18757),
            .I(N__18754));
    Span4Mux_v I__3501 (
            .O(N__18754),
            .I(N__18751));
    Odrv4 I__3500 (
            .O(N__18751),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    CascadeMux I__3499 (
            .O(N__18748),
            .I(N__18745));
    InMux I__3498 (
            .O(N__18745),
            .I(N__18742));
    LocalMux I__3497 (
            .O(N__18742),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__3496 (
            .O(N__18739),
            .I(N__18736));
    LocalMux I__3495 (
            .O(N__18736),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    CascadeMux I__3494 (
            .O(N__18733),
            .I(N__18730));
    InMux I__3493 (
            .O(N__18730),
            .I(N__18727));
    LocalMux I__3492 (
            .O(N__18727),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__3491 (
            .O(N__18724),
            .I(N__18721));
    LocalMux I__3490 (
            .O(N__18721),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__3489 (
            .O(N__18718),
            .I(N__18715));
    LocalMux I__3488 (
            .O(N__18715),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    InMux I__3487 (
            .O(N__18712),
            .I(N__18709));
    LocalMux I__3486 (
            .O(N__18709),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__3485 (
            .O(N__18706),
            .I(N__18703));
    LocalMux I__3484 (
            .O(N__18703),
            .I(N__18700));
    Odrv12 I__3483 (
            .O(N__18700),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    CascadeMux I__3482 (
            .O(N__18697),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ));
    InMux I__3481 (
            .O(N__18694),
            .I(N__18688));
    InMux I__3480 (
            .O(N__18693),
            .I(N__18688));
    LocalMux I__3479 (
            .O(N__18688),
            .I(N__18685));
    Span4Mux_h I__3478 (
            .O(N__18685),
            .I(N__18682));
    Span4Mux_v I__3477 (
            .O(N__18682),
            .I(N__18679));
    Odrv4 I__3476 (
            .O(N__18679),
            .I(\ppm_encoder_1.N_237 ));
    InMux I__3475 (
            .O(N__18676),
            .I(N__18670));
    InMux I__3474 (
            .O(N__18675),
            .I(N__18670));
    LocalMux I__3473 (
            .O(N__18670),
            .I(N__18667));
    Span4Mux_v I__3472 (
            .O(N__18667),
            .I(N__18663));
    InMux I__3471 (
            .O(N__18666),
            .I(N__18660));
    Odrv4 I__3470 (
            .O(N__18663),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__3469 (
            .O(N__18660),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__3468 (
            .O(N__18655),
            .I(N__18651));
    InMux I__3467 (
            .O(N__18654),
            .I(N__18648));
    LocalMux I__3466 (
            .O(N__18651),
            .I(N__18643));
    LocalMux I__3465 (
            .O(N__18648),
            .I(N__18643));
    Span4Mux_h I__3464 (
            .O(N__18643),
            .I(N__18640));
    Odrv4 I__3463 (
            .O(N__18640),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    InMux I__3462 (
            .O(N__18637),
            .I(N__18634));
    LocalMux I__3461 (
            .O(N__18634),
            .I(N__18631));
    Span4Mux_v I__3460 (
            .O(N__18631),
            .I(N__18626));
    InMux I__3459 (
            .O(N__18630),
            .I(N__18621));
    InMux I__3458 (
            .O(N__18629),
            .I(N__18621));
    Odrv4 I__3457 (
            .O(N__18626),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    LocalMux I__3456 (
            .O(N__18621),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__3455 (
            .O(N__18616),
            .I(N__18613));
    LocalMux I__3454 (
            .O(N__18613),
            .I(N__18609));
    InMux I__3453 (
            .O(N__18612),
            .I(N__18606));
    Span4Mux_h I__3452 (
            .O(N__18609),
            .I(N__18600));
    LocalMux I__3451 (
            .O(N__18606),
            .I(N__18600));
    InMux I__3450 (
            .O(N__18605),
            .I(N__18597));
    Span4Mux_v I__3449 (
            .O(N__18600),
            .I(N__18594));
    LocalMux I__3448 (
            .O(N__18597),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__3447 (
            .O(N__18594),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    InMux I__3446 (
            .O(N__18589),
            .I(N__18586));
    LocalMux I__3445 (
            .O(N__18586),
            .I(N__18583));
    Span4Mux_v I__3444 (
            .O(N__18583),
            .I(N__18579));
    InMux I__3443 (
            .O(N__18582),
            .I(N__18576));
    Odrv4 I__3442 (
            .O(N__18579),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    LocalMux I__3441 (
            .O(N__18576),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    InMux I__3440 (
            .O(N__18571),
            .I(N__18567));
    CascadeMux I__3439 (
            .O(N__18570),
            .I(N__18564));
    LocalMux I__3438 (
            .O(N__18567),
            .I(N__18558));
    InMux I__3437 (
            .O(N__18564),
            .I(N__18555));
    InMux I__3436 (
            .O(N__18563),
            .I(N__18552));
    InMux I__3435 (
            .O(N__18562),
            .I(N__18547));
    InMux I__3434 (
            .O(N__18561),
            .I(N__18547));
    Span4Mux_h I__3433 (
            .O(N__18558),
            .I(N__18542));
    LocalMux I__3432 (
            .O(N__18555),
            .I(N__18542));
    LocalMux I__3431 (
            .O(N__18552),
            .I(N__18539));
    LocalMux I__3430 (
            .O(N__18547),
            .I(N__18532));
    Span4Mux_v I__3429 (
            .O(N__18542),
            .I(N__18532));
    Span4Mux_h I__3428 (
            .O(N__18539),
            .I(N__18529));
    InMux I__3427 (
            .O(N__18538),
            .I(N__18524));
    InMux I__3426 (
            .O(N__18537),
            .I(N__18524));
    Odrv4 I__3425 (
            .O(N__18532),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__3424 (
            .O(N__18529),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__3423 (
            .O(N__18524),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__3422 (
            .O(N__18517),
            .I(\ppm_encoder_1.N_296_cascade_ ));
    InMux I__3421 (
            .O(N__18514),
            .I(N__18511));
    LocalMux I__3420 (
            .O(N__18511),
            .I(N__18508));
    Span4Mux_v I__3419 (
            .O(N__18508),
            .I(N__18504));
    InMux I__3418 (
            .O(N__18507),
            .I(N__18501));
    Odrv4 I__3417 (
            .O(N__18504),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    LocalMux I__3416 (
            .O(N__18501),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__3415 (
            .O(N__18496),
            .I(N__18493));
    LocalMux I__3414 (
            .O(N__18493),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    InMux I__3413 (
            .O(N__18490),
            .I(N__18487));
    LocalMux I__3412 (
            .O(N__18487),
            .I(N__18481));
    InMux I__3411 (
            .O(N__18486),
            .I(N__18474));
    InMux I__3410 (
            .O(N__18485),
            .I(N__18474));
    InMux I__3409 (
            .O(N__18484),
            .I(N__18474));
    Odrv12 I__3408 (
            .O(N__18481),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    LocalMux I__3407 (
            .O(N__18474),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    InMux I__3406 (
            .O(N__18469),
            .I(N__18466));
    LocalMux I__3405 (
            .O(N__18466),
            .I(N__18463));
    Span4Mux_h I__3404 (
            .O(N__18463),
            .I(N__18457));
    InMux I__3403 (
            .O(N__18462),
            .I(N__18450));
    InMux I__3402 (
            .O(N__18461),
            .I(N__18450));
    InMux I__3401 (
            .O(N__18460),
            .I(N__18450));
    Odrv4 I__3400 (
            .O(N__18457),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__3399 (
            .O(N__18450),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__3398 (
            .O(N__18445),
            .I(N__18442));
    LocalMux I__3397 (
            .O(N__18442),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__3396 (
            .O(N__18439),
            .I(N__18436));
    LocalMux I__3395 (
            .O(N__18436),
            .I(N__18433));
    Span4Mux_h I__3394 (
            .O(N__18433),
            .I(N__18430));
    Odrv4 I__3393 (
            .O(N__18430),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__3392 (
            .O(N__18427),
            .I(N__18424));
    LocalMux I__3391 (
            .O(N__18424),
            .I(N__18421));
    Span4Mux_s3_v I__3390 (
            .O(N__18421),
            .I(N__18418));
    Odrv4 I__3389 (
            .O(N__18418),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    InMux I__3388 (
            .O(N__18415),
            .I(N__18412));
    LocalMux I__3387 (
            .O(N__18412),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CascadeMux I__3386 (
            .O(N__18409),
            .I(N__18406));
    InMux I__3385 (
            .O(N__18406),
            .I(N__18397));
    InMux I__3384 (
            .O(N__18405),
            .I(N__18397));
    InMux I__3383 (
            .O(N__18404),
            .I(N__18397));
    LocalMux I__3382 (
            .O(N__18397),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__3381 (
            .O(N__18394),
            .I(N__18391));
    LocalMux I__3380 (
            .O(N__18391),
            .I(N__18388));
    Odrv4 I__3379 (
            .O(N__18388),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__3378 (
            .O(N__18385),
            .I(N__18382));
    LocalMux I__3377 (
            .O(N__18382),
            .I(N__18379));
    Span4Mux_h I__3376 (
            .O(N__18379),
            .I(N__18376));
    Span4Mux_h I__3375 (
            .O(N__18376),
            .I(N__18373));
    Odrv4 I__3374 (
            .O(N__18373),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__3373 (
            .O(N__18370),
            .I(N__18367));
    LocalMux I__3372 (
            .O(N__18367),
            .I(N__18364));
    Odrv4 I__3371 (
            .O(N__18364),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__3370 (
            .O(N__18361),
            .I(N__18358));
    LocalMux I__3369 (
            .O(N__18358),
            .I(N__18354));
    InMux I__3368 (
            .O(N__18357),
            .I(N__18351));
    Span4Mux_h I__3367 (
            .O(N__18354),
            .I(N__18348));
    LocalMux I__3366 (
            .O(N__18351),
            .I(N__18345));
    Odrv4 I__3365 (
            .O(N__18348),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    Odrv4 I__3364 (
            .O(N__18345),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    InMux I__3363 (
            .O(N__18340),
            .I(N__18337));
    LocalMux I__3362 (
            .O(N__18337),
            .I(N__18334));
    Span4Mux_h I__3361 (
            .O(N__18334),
            .I(N__18331));
    Odrv4 I__3360 (
            .O(N__18331),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    CascadeMux I__3359 (
            .O(N__18328),
            .I(N__18325));
    InMux I__3358 (
            .O(N__18325),
            .I(N__18322));
    LocalMux I__3357 (
            .O(N__18322),
            .I(N__18319));
    Odrv4 I__3356 (
            .O(N__18319),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__3355 (
            .O(N__18316),
            .I(N__18313));
    LocalMux I__3354 (
            .O(N__18313),
            .I(N__18310));
    Span4Mux_h I__3353 (
            .O(N__18310),
            .I(N__18307));
    Odrv4 I__3352 (
            .O(N__18307),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__3351 (
            .O(N__18304),
            .I(N__18301));
    LocalMux I__3350 (
            .O(N__18301),
            .I(N__18298));
    Odrv4 I__3349 (
            .O(N__18298),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__3348 (
            .O(N__18295),
            .I(N__18291));
    InMux I__3347 (
            .O(N__18294),
            .I(N__18288));
    LocalMux I__3346 (
            .O(N__18291),
            .I(N__18285));
    LocalMux I__3345 (
            .O(N__18288),
            .I(N__18282));
    Odrv4 I__3344 (
            .O(N__18285),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    Odrv4 I__3343 (
            .O(N__18282),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    InMux I__3342 (
            .O(N__18277),
            .I(N__18274));
    LocalMux I__3341 (
            .O(N__18274),
            .I(N__18271));
    Span4Mux_h I__3340 (
            .O(N__18271),
            .I(N__18268));
    Odrv4 I__3339 (
            .O(N__18268),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    CascadeMux I__3338 (
            .O(N__18265),
            .I(N__18262));
    InMux I__3337 (
            .O(N__18262),
            .I(N__18259));
    LocalMux I__3336 (
            .O(N__18259),
            .I(N__18256));
    Span4Mux_v I__3335 (
            .O(N__18256),
            .I(N__18253));
    Odrv4 I__3334 (
            .O(N__18253),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__3333 (
            .O(N__18250),
            .I(N__18245));
    InMux I__3332 (
            .O(N__18249),
            .I(N__18238));
    InMux I__3331 (
            .O(N__18248),
            .I(N__18238));
    LocalMux I__3330 (
            .O(N__18245),
            .I(N__18235));
    InMux I__3329 (
            .O(N__18244),
            .I(N__18232));
    InMux I__3328 (
            .O(N__18243),
            .I(N__18228));
    LocalMux I__3327 (
            .O(N__18238),
            .I(N__18224));
    Span4Mux_v I__3326 (
            .O(N__18235),
            .I(N__18221));
    LocalMux I__3325 (
            .O(N__18232),
            .I(N__18218));
    InMux I__3324 (
            .O(N__18231),
            .I(N__18215));
    LocalMux I__3323 (
            .O(N__18228),
            .I(N__18212));
    InMux I__3322 (
            .O(N__18227),
            .I(N__18206));
    Span4Mux_v I__3321 (
            .O(N__18224),
            .I(N__18195));
    Span4Mux_h I__3320 (
            .O(N__18221),
            .I(N__18192));
    Span4Mux_h I__3319 (
            .O(N__18218),
            .I(N__18187));
    LocalMux I__3318 (
            .O(N__18215),
            .I(N__18187));
    Span4Mux_h I__3317 (
            .O(N__18212),
            .I(N__18184));
    InMux I__3316 (
            .O(N__18211),
            .I(N__18177));
    InMux I__3315 (
            .O(N__18210),
            .I(N__18177));
    InMux I__3314 (
            .O(N__18209),
            .I(N__18177));
    LocalMux I__3313 (
            .O(N__18206),
            .I(N__18174));
    InMux I__3312 (
            .O(N__18205),
            .I(N__18171));
    InMux I__3311 (
            .O(N__18204),
            .I(N__18166));
    InMux I__3310 (
            .O(N__18203),
            .I(N__18166));
    InMux I__3309 (
            .O(N__18202),
            .I(N__18161));
    InMux I__3308 (
            .O(N__18201),
            .I(N__18161));
    InMux I__3307 (
            .O(N__18200),
            .I(N__18158));
    InMux I__3306 (
            .O(N__18199),
            .I(N__18153));
    InMux I__3305 (
            .O(N__18198),
            .I(N__18153));
    Odrv4 I__3304 (
            .O(N__18195),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__3303 (
            .O(N__18192),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__3302 (
            .O(N__18187),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__3301 (
            .O(N__18184),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3300 (
            .O(N__18177),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv12 I__3299 (
            .O(N__18174),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3298 (
            .O(N__18171),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3297 (
            .O(N__18166),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3296 (
            .O(N__18161),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3295 (
            .O(N__18158),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3294 (
            .O(N__18153),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__3293 (
            .O(N__18130),
            .I(N__18127));
    LocalMux I__3292 (
            .O(N__18127),
            .I(N__18124));
    Span4Mux_h I__3291 (
            .O(N__18124),
            .I(N__18121));
    Span4Mux_s2_h I__3290 (
            .O(N__18121),
            .I(N__18118));
    Odrv4 I__3289 (
            .O(N__18118),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    CascadeMux I__3288 (
            .O(N__18115),
            .I(N__18104));
    CascadeMux I__3287 (
            .O(N__18114),
            .I(N__18101));
    CascadeMux I__3286 (
            .O(N__18113),
            .I(N__18098));
    CascadeMux I__3285 (
            .O(N__18112),
            .I(N__18095));
    CascadeMux I__3284 (
            .O(N__18111),
            .I(N__18091));
    CascadeMux I__3283 (
            .O(N__18110),
            .I(N__18087));
    CascadeMux I__3282 (
            .O(N__18109),
            .I(N__18084));
    CascadeMux I__3281 (
            .O(N__18108),
            .I(N__18081));
    InMux I__3280 (
            .O(N__18107),
            .I(N__18072));
    InMux I__3279 (
            .O(N__18104),
            .I(N__18072));
    InMux I__3278 (
            .O(N__18101),
            .I(N__18072));
    InMux I__3277 (
            .O(N__18098),
            .I(N__18067));
    InMux I__3276 (
            .O(N__18095),
            .I(N__18067));
    CascadeMux I__3275 (
            .O(N__18094),
            .I(N__18064));
    InMux I__3274 (
            .O(N__18091),
            .I(N__18055));
    InMux I__3273 (
            .O(N__18090),
            .I(N__18055));
    InMux I__3272 (
            .O(N__18087),
            .I(N__18055));
    InMux I__3271 (
            .O(N__18084),
            .I(N__18050));
    InMux I__3270 (
            .O(N__18081),
            .I(N__18050));
    CascadeMux I__3269 (
            .O(N__18080),
            .I(N__18046));
    CascadeMux I__3268 (
            .O(N__18079),
            .I(N__18042));
    LocalMux I__3267 (
            .O(N__18072),
            .I(N__18039));
    LocalMux I__3266 (
            .O(N__18067),
            .I(N__18036));
    InMux I__3265 (
            .O(N__18064),
            .I(N__18033));
    InMux I__3264 (
            .O(N__18063),
            .I(N__18030));
    CascadeMux I__3263 (
            .O(N__18062),
            .I(N__18027));
    LocalMux I__3262 (
            .O(N__18055),
            .I(N__18023));
    LocalMux I__3261 (
            .O(N__18050),
            .I(N__18020));
    InMux I__3260 (
            .O(N__18049),
            .I(N__18011));
    InMux I__3259 (
            .O(N__18046),
            .I(N__18011));
    InMux I__3258 (
            .O(N__18045),
            .I(N__18011));
    InMux I__3257 (
            .O(N__18042),
            .I(N__18011));
    Span4Mux_v I__3256 (
            .O(N__18039),
            .I(N__18001));
    Span4Mux_s2_v I__3255 (
            .O(N__18036),
            .I(N__18001));
    LocalMux I__3254 (
            .O(N__18033),
            .I(N__18001));
    LocalMux I__3253 (
            .O(N__18030),
            .I(N__18001));
    InMux I__3252 (
            .O(N__18027),
            .I(N__17998));
    CascadeMux I__3251 (
            .O(N__18026),
            .I(N__17995));
    Span4Mux_v I__3250 (
            .O(N__18023),
            .I(N__17988));
    Span4Mux_h I__3249 (
            .O(N__18020),
            .I(N__17988));
    LocalMux I__3248 (
            .O(N__18011),
            .I(N__17988));
    InMux I__3247 (
            .O(N__18010),
            .I(N__17985));
    Span4Mux_h I__3246 (
            .O(N__18001),
            .I(N__17980));
    LocalMux I__3245 (
            .O(N__17998),
            .I(N__17980));
    InMux I__3244 (
            .O(N__17995),
            .I(N__17977));
    Odrv4 I__3243 (
            .O(N__17988),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__3242 (
            .O(N__17985),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__3241 (
            .O(N__17980),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__3240 (
            .O(N__17977),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__3239 (
            .O(N__17968),
            .I(N__17965));
    LocalMux I__3238 (
            .O(N__17965),
            .I(N__17962));
    Span4Mux_v I__3237 (
            .O(N__17962),
            .I(N__17959));
    Odrv4 I__3236 (
            .O(N__17959),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__3235 (
            .O(N__17956),
            .I(N__17953));
    LocalMux I__3234 (
            .O(N__17953),
            .I(N__17948));
    InMux I__3233 (
            .O(N__17952),
            .I(N__17945));
    CascadeMux I__3232 (
            .O(N__17951),
            .I(N__17942));
    Span4Mux_h I__3231 (
            .O(N__17948),
            .I(N__17938));
    LocalMux I__3230 (
            .O(N__17945),
            .I(N__17935));
    InMux I__3229 (
            .O(N__17942),
            .I(N__17930));
    InMux I__3228 (
            .O(N__17941),
            .I(N__17930));
    Odrv4 I__3227 (
            .O(N__17938),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv12 I__3226 (
            .O(N__17935),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__3225 (
            .O(N__17930),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__3224 (
            .O(N__17923),
            .I(N__17920));
    LocalMux I__3223 (
            .O(N__17920),
            .I(N__17915));
    InMux I__3222 (
            .O(N__17919),
            .I(N__17912));
    InMux I__3221 (
            .O(N__17918),
            .I(N__17909));
    Span4Mux_h I__3220 (
            .O(N__17915),
            .I(N__17904));
    LocalMux I__3219 (
            .O(N__17912),
            .I(N__17904));
    LocalMux I__3218 (
            .O(N__17909),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    Odrv4 I__3217 (
            .O(N__17904),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    CascadeMux I__3216 (
            .O(N__17899),
            .I(N__17895));
    CascadeMux I__3215 (
            .O(N__17898),
            .I(N__17891));
    InMux I__3214 (
            .O(N__17895),
            .I(N__17888));
    InMux I__3213 (
            .O(N__17894),
            .I(N__17885));
    InMux I__3212 (
            .O(N__17891),
            .I(N__17882));
    LocalMux I__3211 (
            .O(N__17888),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    LocalMux I__3210 (
            .O(N__17885),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    LocalMux I__3209 (
            .O(N__17882),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    CascadeMux I__3208 (
            .O(N__17875),
            .I(\ppm_encoder_1.N_302_cascade_ ));
    InMux I__3207 (
            .O(N__17872),
            .I(N__17869));
    LocalMux I__3206 (
            .O(N__17869),
            .I(N__17866));
    Span4Mux_s3_v I__3205 (
            .O(N__17866),
            .I(N__17863));
    Odrv4 I__3204 (
            .O(N__17863),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__3203 (
            .O(N__17860),
            .I(N__17852));
    InMux I__3202 (
            .O(N__17859),
            .I(N__17852));
    InMux I__3201 (
            .O(N__17858),
            .I(N__17847));
    InMux I__3200 (
            .O(N__17857),
            .I(N__17847));
    LocalMux I__3199 (
            .O(N__17852),
            .I(N__17844));
    LocalMux I__3198 (
            .O(N__17847),
            .I(N__17839));
    Span4Mux_h I__3197 (
            .O(N__17844),
            .I(N__17836));
    InMux I__3196 (
            .O(N__17843),
            .I(N__17831));
    InMux I__3195 (
            .O(N__17842),
            .I(N__17831));
    Odrv4 I__3194 (
            .O(N__17839),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__3193 (
            .O(N__17836),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__3192 (
            .O(N__17831),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__3191 (
            .O(N__17824),
            .I(N__17820));
    InMux I__3190 (
            .O(N__17823),
            .I(N__17815));
    InMux I__3189 (
            .O(N__17820),
            .I(N__17810));
    InMux I__3188 (
            .O(N__17819),
            .I(N__17810));
    InMux I__3187 (
            .O(N__17818),
            .I(N__17805));
    LocalMux I__3186 (
            .O(N__17815),
            .I(N__17802));
    LocalMux I__3185 (
            .O(N__17810),
            .I(N__17798));
    InMux I__3184 (
            .O(N__17809),
            .I(N__17793));
    InMux I__3183 (
            .O(N__17808),
            .I(N__17793));
    LocalMux I__3182 (
            .O(N__17805),
            .I(N__17788));
    Span4Mux_v I__3181 (
            .O(N__17802),
            .I(N__17788));
    InMux I__3180 (
            .O(N__17801),
            .I(N__17785));
    Span4Mux_h I__3179 (
            .O(N__17798),
            .I(N__17780));
    LocalMux I__3178 (
            .O(N__17793),
            .I(N__17780));
    Odrv4 I__3177 (
            .O(N__17788),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__3176 (
            .O(N__17785),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__3175 (
            .O(N__17780),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__3174 (
            .O(N__17773),
            .I(N__17770));
    LocalMux I__3173 (
            .O(N__17770),
            .I(N__17767));
    Span4Mux_v I__3172 (
            .O(N__17767),
            .I(N__17764));
    Odrv4 I__3171 (
            .O(N__17764),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__3170 (
            .O(N__17761),
            .I(N__17758));
    LocalMux I__3169 (
            .O(N__17758),
            .I(N__17755));
    Odrv4 I__3168 (
            .O(N__17755),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__3167 (
            .O(N__17752),
            .I(N__17749));
    LocalMux I__3166 (
            .O(N__17749),
            .I(N__17746));
    Span4Mux_v I__3165 (
            .O(N__17746),
            .I(N__17742));
    InMux I__3164 (
            .O(N__17745),
            .I(N__17739));
    Sp12to4 I__3163 (
            .O(N__17742),
            .I(N__17734));
    LocalMux I__3162 (
            .O(N__17739),
            .I(N__17734));
    Odrv12 I__3161 (
            .O(N__17734),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__3160 (
            .O(N__17731),
            .I(N__17728));
    LocalMux I__3159 (
            .O(N__17728),
            .I(N__17725));
    Span4Mux_h I__3158 (
            .O(N__17725),
            .I(N__17722));
    Odrv4 I__3157 (
            .O(N__17722),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__3156 (
            .O(N__17719),
            .I(N__17716));
    LocalMux I__3155 (
            .O(N__17716),
            .I(N__17712));
    InMux I__3154 (
            .O(N__17715),
            .I(N__17709));
    Odrv4 I__3153 (
            .O(N__17712),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    LocalMux I__3152 (
            .O(N__17709),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__3151 (
            .O(N__17704),
            .I(N__17701));
    LocalMux I__3150 (
            .O(N__17701),
            .I(\uart_pc.data_Auxce_0_3 ));
    CascadeMux I__3149 (
            .O(N__17698),
            .I(N__17695));
    InMux I__3148 (
            .O(N__17695),
            .I(N__17692));
    LocalMux I__3147 (
            .O(N__17692),
            .I(N__17689));
    Span4Mux_h I__3146 (
            .O(N__17689),
            .I(N__17685));
    InMux I__3145 (
            .O(N__17688),
            .I(N__17682));
    Odrv4 I__3144 (
            .O(N__17685),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__3143 (
            .O(N__17682),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__3142 (
            .O(N__17677),
            .I(N__17674));
    LocalMux I__3141 (
            .O(N__17674),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__3140 (
            .O(N__17671),
            .I(N__17667));
    CascadeMux I__3139 (
            .O(N__17670),
            .I(N__17664));
    LocalMux I__3138 (
            .O(N__17667),
            .I(N__17661));
    InMux I__3137 (
            .O(N__17664),
            .I(N__17658));
    Odrv4 I__3136 (
            .O(N__17661),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__3135 (
            .O(N__17658),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__3134 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__3133 (
            .O(N__17650),
            .I(\uart_pc.data_Auxce_0_5 ));
    CascadeMux I__3132 (
            .O(N__17647),
            .I(N__17644));
    InMux I__3131 (
            .O(N__17644),
            .I(N__17641));
    LocalMux I__3130 (
            .O(N__17641),
            .I(N__17638));
    Span4Mux_v I__3129 (
            .O(N__17638),
            .I(N__17634));
    InMux I__3128 (
            .O(N__17637),
            .I(N__17631));
    Odrv4 I__3127 (
            .O(N__17634),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__3126 (
            .O(N__17631),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__3125 (
            .O(N__17626),
            .I(N__17623));
    InMux I__3124 (
            .O(N__17623),
            .I(N__17620));
    LocalMux I__3123 (
            .O(N__17620),
            .I(N__17617));
    Span4Mux_h I__3122 (
            .O(N__17617),
            .I(N__17613));
    InMux I__3121 (
            .O(N__17616),
            .I(N__17610));
    Odrv4 I__3120 (
            .O(N__17613),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__3119 (
            .O(N__17610),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    InMux I__3118 (
            .O(N__17605),
            .I(N__17602));
    LocalMux I__3117 (
            .O(N__17602),
            .I(N__17599));
    Span4Mux_v I__3116 (
            .O(N__17599),
            .I(N__17596));
    Odrv4 I__3115 (
            .O(N__17596),
            .I(\uart_pc.data_Auxce_0_6 ));
    CascadeMux I__3114 (
            .O(N__17593),
            .I(N__17590));
    InMux I__3113 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__3112 (
            .O(N__17587),
            .I(N__17583));
    CascadeMux I__3111 (
            .O(N__17586),
            .I(N__17580));
    Span4Mux_v I__3110 (
            .O(N__17583),
            .I(N__17577));
    InMux I__3109 (
            .O(N__17580),
            .I(N__17574));
    Odrv4 I__3108 (
            .O(N__17577),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__3107 (
            .O(N__17574),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    CascadeMux I__3106 (
            .O(N__17569),
            .I(N__17566));
    InMux I__3105 (
            .O(N__17566),
            .I(N__17562));
    InMux I__3104 (
            .O(N__17565),
            .I(N__17559));
    LocalMux I__3103 (
            .O(N__17562),
            .I(N__17556));
    LocalMux I__3102 (
            .O(N__17559),
            .I(N__17553));
    Span4Mux_h I__3101 (
            .O(N__17556),
            .I(N__17549));
    Span4Mux_h I__3100 (
            .O(N__17553),
            .I(N__17546));
    InMux I__3099 (
            .O(N__17552),
            .I(N__17543));
    Odrv4 I__3098 (
            .O(N__17549),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__3097 (
            .O(N__17546),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__3096 (
            .O(N__17543),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__3095 (
            .O(N__17536),
            .I(N__17532));
    InMux I__3094 (
            .O(N__17535),
            .I(N__17529));
    LocalMux I__3093 (
            .O(N__17532),
            .I(N__17526));
    LocalMux I__3092 (
            .O(N__17529),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    Odrv4 I__3091 (
            .O(N__17526),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    CascadeMux I__3090 (
            .O(N__17521),
            .I(N__17517));
    InMux I__3089 (
            .O(N__17520),
            .I(N__17510));
    InMux I__3088 (
            .O(N__17517),
            .I(N__17510));
    InMux I__3087 (
            .O(N__17516),
            .I(N__17505));
    InMux I__3086 (
            .O(N__17515),
            .I(N__17505));
    LocalMux I__3085 (
            .O(N__17510),
            .I(N__17502));
    LocalMux I__3084 (
            .O(N__17505),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    Odrv4 I__3083 (
            .O(N__17502),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__3082 (
            .O(N__17497),
            .I(N__17494));
    InMux I__3081 (
            .O(N__17494),
            .I(N__17491));
    LocalMux I__3080 (
            .O(N__17491),
            .I(N__17488));
    Odrv4 I__3079 (
            .O(N__17488),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    InMux I__3078 (
            .O(N__17485),
            .I(N__17480));
    InMux I__3077 (
            .O(N__17484),
            .I(N__17475));
    InMux I__3076 (
            .O(N__17483),
            .I(N__17475));
    LocalMux I__3075 (
            .O(N__17480),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__3074 (
            .O(N__17475),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__3073 (
            .O(N__17470),
            .I(N__17467));
    LocalMux I__3072 (
            .O(N__17467),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__3071 (
            .O(N__17464),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__3070 (
            .O(N__17461),
            .I(N__17458));
    LocalMux I__3069 (
            .O(N__17458),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__3068 (
            .O(N__17455),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__3067 (
            .O(N__17452),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__3066 (
            .O(N__17449),
            .I(N__17446));
    LocalMux I__3065 (
            .O(N__17446),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    CascadeMux I__3064 (
            .O(N__17443),
            .I(N__17440));
    InMux I__3063 (
            .O(N__17440),
            .I(N__17433));
    InMux I__3062 (
            .O(N__17439),
            .I(N__17433));
    InMux I__3061 (
            .O(N__17438),
            .I(N__17429));
    LocalMux I__3060 (
            .O(N__17433),
            .I(N__17426));
    InMux I__3059 (
            .O(N__17432),
            .I(N__17423));
    LocalMux I__3058 (
            .O(N__17429),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__3057 (
            .O(N__17426),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__3056 (
            .O(N__17423),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    InMux I__3055 (
            .O(N__17416),
            .I(N__17412));
    CascadeMux I__3054 (
            .O(N__17415),
            .I(N__17409));
    LocalMux I__3053 (
            .O(N__17412),
            .I(N__17406));
    InMux I__3052 (
            .O(N__17409),
            .I(N__17403));
    Odrv4 I__3051 (
            .O(N__17406),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__3050 (
            .O(N__17403),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__3049 (
            .O(N__17398),
            .I(N__17394));
    InMux I__3048 (
            .O(N__17397),
            .I(N__17391));
    LocalMux I__3047 (
            .O(N__17394),
            .I(N__17381));
    LocalMux I__3046 (
            .O(N__17391),
            .I(N__17381));
    InMux I__3045 (
            .O(N__17390),
            .I(N__17372));
    InMux I__3044 (
            .O(N__17389),
            .I(N__17372));
    InMux I__3043 (
            .O(N__17388),
            .I(N__17372));
    InMux I__3042 (
            .O(N__17387),
            .I(N__17372));
    InMux I__3041 (
            .O(N__17386),
            .I(N__17367));
    Span4Mux_v I__3040 (
            .O(N__17381),
            .I(N__17362));
    LocalMux I__3039 (
            .O(N__17372),
            .I(N__17362));
    InMux I__3038 (
            .O(N__17371),
            .I(N__17357));
    InMux I__3037 (
            .O(N__17370),
            .I(N__17357));
    LocalMux I__3036 (
            .O(N__17367),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    Odrv4 I__3035 (
            .O(N__17362),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__3034 (
            .O(N__17357),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__3033 (
            .O(N__17350),
            .I(N__17345));
    InMux I__3032 (
            .O(N__17349),
            .I(N__17342));
    CascadeMux I__3031 (
            .O(N__17348),
            .I(N__17336));
    LocalMux I__3030 (
            .O(N__17345),
            .I(N__17333));
    LocalMux I__3029 (
            .O(N__17342),
            .I(N__17330));
    CascadeMux I__3028 (
            .O(N__17341),
            .I(N__17327));
    CascadeMux I__3027 (
            .O(N__17340),
            .I(N__17323));
    InMux I__3026 (
            .O(N__17339),
            .I(N__17315));
    InMux I__3025 (
            .O(N__17336),
            .I(N__17315));
    Span4Mux_v I__3024 (
            .O(N__17333),
            .I(N__17312));
    Span4Mux_h I__3023 (
            .O(N__17330),
            .I(N__17309));
    InMux I__3022 (
            .O(N__17327),
            .I(N__17300));
    InMux I__3021 (
            .O(N__17326),
            .I(N__17300));
    InMux I__3020 (
            .O(N__17323),
            .I(N__17300));
    InMux I__3019 (
            .O(N__17322),
            .I(N__17300));
    InMux I__3018 (
            .O(N__17321),
            .I(N__17295));
    InMux I__3017 (
            .O(N__17320),
            .I(N__17295));
    LocalMux I__3016 (
            .O(N__17315),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv4 I__3015 (
            .O(N__17312),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv4 I__3014 (
            .O(N__17309),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__3013 (
            .O(N__17300),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__3012 (
            .O(N__17295),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__3011 (
            .O(N__17284),
            .I(N__17274));
    CascadeMux I__3010 (
            .O(N__17283),
            .I(N__17270));
    InMux I__3009 (
            .O(N__17282),
            .I(N__17265));
    InMux I__3008 (
            .O(N__17281),
            .I(N__17265));
    InMux I__3007 (
            .O(N__17280),
            .I(N__17256));
    InMux I__3006 (
            .O(N__17279),
            .I(N__17256));
    InMux I__3005 (
            .O(N__17278),
            .I(N__17256));
    InMux I__3004 (
            .O(N__17277),
            .I(N__17256));
    LocalMux I__3003 (
            .O(N__17274),
            .I(N__17253));
    InMux I__3002 (
            .O(N__17273),
            .I(N__17250));
    InMux I__3001 (
            .O(N__17270),
            .I(N__17245));
    LocalMux I__3000 (
            .O(N__17265),
            .I(N__17240));
    LocalMux I__2999 (
            .O(N__17256),
            .I(N__17240));
    Span4Mux_v I__2998 (
            .O(N__17253),
            .I(N__17235));
    LocalMux I__2997 (
            .O(N__17250),
            .I(N__17235));
    InMux I__2996 (
            .O(N__17249),
            .I(N__17230));
    InMux I__2995 (
            .O(N__17248),
            .I(N__17230));
    LocalMux I__2994 (
            .O(N__17245),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv4 I__2993 (
            .O(N__17240),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv4 I__2992 (
            .O(N__17235),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__2991 (
            .O(N__17230),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    InMux I__2990 (
            .O(N__17221),
            .I(N__17218));
    LocalMux I__2989 (
            .O(N__17218),
            .I(N__17215));
    Odrv4 I__2988 (
            .O(N__17215),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    InMux I__2987 (
            .O(N__17212),
            .I(N__17208));
    CascadeMux I__2986 (
            .O(N__17211),
            .I(N__17205));
    LocalMux I__2985 (
            .O(N__17208),
            .I(N__17202));
    InMux I__2984 (
            .O(N__17205),
            .I(N__17199));
    Odrv12 I__2983 (
            .O(N__17202),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__2982 (
            .O(N__17199),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    InMux I__2981 (
            .O(N__17194),
            .I(N__17191));
    LocalMux I__2980 (
            .O(N__17191),
            .I(\uart_pc.data_Auxce_0_1 ));
    InMux I__2979 (
            .O(N__17188),
            .I(N__17185));
    LocalMux I__2978 (
            .O(N__17185),
            .I(N__17182));
    Span4Mux_h I__2977 (
            .O(N__17182),
            .I(N__17178));
    InMux I__2976 (
            .O(N__17181),
            .I(N__17175));
    Odrv4 I__2975 (
            .O(N__17178),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__2974 (
            .O(N__17175),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__2973 (
            .O(N__17170),
            .I(N__17167));
    LocalMux I__2972 (
            .O(N__17167),
            .I(N__17164));
    Span4Mux_h I__2971 (
            .O(N__17164),
            .I(N__17161));
    Odrv4 I__2970 (
            .O(N__17161),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    CascadeMux I__2969 (
            .O(N__17158),
            .I(N__17155));
    InMux I__2968 (
            .O(N__17155),
            .I(N__17151));
    CascadeMux I__2967 (
            .O(N__17154),
            .I(N__17148));
    LocalMux I__2966 (
            .O(N__17151),
            .I(N__17145));
    InMux I__2965 (
            .O(N__17148),
            .I(N__17142));
    Odrv12 I__2964 (
            .O(N__17145),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__2963 (
            .O(N__17142),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    InMux I__2962 (
            .O(N__17137),
            .I(N__17132));
    InMux I__2961 (
            .O(N__17136),
            .I(N__17127));
    InMux I__2960 (
            .O(N__17135),
            .I(N__17127));
    LocalMux I__2959 (
            .O(N__17132),
            .I(N__17124));
    LocalMux I__2958 (
            .O(N__17127),
            .I(N__17121));
    Odrv4 I__2957 (
            .O(N__17124),
            .I(\uart_drone.state_1_sqmuxa ));
    Odrv4 I__2956 (
            .O(N__17121),
            .I(\uart_drone.state_1_sqmuxa ));
    SRMux I__2955 (
            .O(N__17116),
            .I(N__17113));
    LocalMux I__2954 (
            .O(N__17113),
            .I(N__17109));
    SRMux I__2953 (
            .O(N__17112),
            .I(N__17106));
    Sp12to4 I__2952 (
            .O(N__17109),
            .I(N__17103));
    LocalMux I__2951 (
            .O(N__17106),
            .I(N__17100));
    Odrv12 I__2950 (
            .O(N__17103),
            .I(\Commands_frame_decoder.un1_state49_iZ0 ));
    Odrv12 I__2949 (
            .O(N__17100),
            .I(\Commands_frame_decoder.un1_state49_iZ0 ));
    CascadeMux I__2948 (
            .O(N__17095),
            .I(\uart_drone.N_126_li_cascade_ ));
    CascadeMux I__2947 (
            .O(N__17092),
            .I(\uart_drone.N_143_cascade_ ));
    CascadeMux I__2946 (
            .O(N__17089),
            .I(N__17085));
    InMux I__2945 (
            .O(N__17088),
            .I(N__17082));
    InMux I__2944 (
            .O(N__17085),
            .I(N__17079));
    LocalMux I__2943 (
            .O(N__17082),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__2942 (
            .O(N__17079),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__2941 (
            .O(N__17074),
            .I(N__17070));
    InMux I__2940 (
            .O(N__17073),
            .I(N__17067));
    InMux I__2939 (
            .O(N__17070),
            .I(N__17064));
    LocalMux I__2938 (
            .O(N__17067),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__2937 (
            .O(N__17064),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__2936 (
            .O(N__17059),
            .I(N__17055));
    InMux I__2935 (
            .O(N__17058),
            .I(N__17052));
    InMux I__2934 (
            .O(N__17055),
            .I(N__17049));
    LocalMux I__2933 (
            .O(N__17052),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__2932 (
            .O(N__17049),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CascadeMux I__2931 (
            .O(N__17044),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    InMux I__2930 (
            .O(N__17041),
            .I(N__17038));
    LocalMux I__2929 (
            .O(N__17038),
            .I(N__17033));
    InMux I__2928 (
            .O(N__17037),
            .I(N__17030));
    InMux I__2927 (
            .O(N__17036),
            .I(N__17027));
    Span4Mux_h I__2926 (
            .O(N__17033),
            .I(N__17019));
    LocalMux I__2925 (
            .O(N__17030),
            .I(N__17019));
    LocalMux I__2924 (
            .O(N__17027),
            .I(N__17016));
    InMux I__2923 (
            .O(N__17026),
            .I(N__17011));
    InMux I__2922 (
            .O(N__17025),
            .I(N__17011));
    InMux I__2921 (
            .O(N__17024),
            .I(N__17008));
    Odrv4 I__2920 (
            .O(N__17019),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    Odrv4 I__2919 (
            .O(N__17016),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__2918 (
            .O(N__17011),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__2917 (
            .O(N__17008),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__2916 (
            .O(N__16999),
            .I(N__16996));
    LocalMux I__2915 (
            .O(N__16996),
            .I(N__16988));
    InMux I__2914 (
            .O(N__16995),
            .I(N__16982));
    InMux I__2913 (
            .O(N__16994),
            .I(N__16982));
    InMux I__2912 (
            .O(N__16993),
            .I(N__16975));
    InMux I__2911 (
            .O(N__16992),
            .I(N__16975));
    InMux I__2910 (
            .O(N__16991),
            .I(N__16975));
    Span4Mux_v I__2909 (
            .O(N__16988),
            .I(N__16972));
    InMux I__2908 (
            .O(N__16987),
            .I(N__16968));
    LocalMux I__2907 (
            .O(N__16982),
            .I(N__16963));
    LocalMux I__2906 (
            .O(N__16975),
            .I(N__16963));
    Span4Mux_h I__2905 (
            .O(N__16972),
            .I(N__16960));
    InMux I__2904 (
            .O(N__16971),
            .I(N__16957));
    LocalMux I__2903 (
            .O(N__16968),
            .I(N__16952));
    Span4Mux_v I__2902 (
            .O(N__16963),
            .I(N__16952));
    Odrv4 I__2901 (
            .O(N__16960),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__2900 (
            .O(N__16957),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__2899 (
            .O(N__16952),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    InMux I__2898 (
            .O(N__16945),
            .I(N__16939));
    InMux I__2897 (
            .O(N__16944),
            .I(N__16939));
    LocalMux I__2896 (
            .O(N__16939),
            .I(\Commands_frame_decoder.state_1Z0Z_5 ));
    InMux I__2895 (
            .O(N__16936),
            .I(N__16933));
    LocalMux I__2894 (
            .O(N__16933),
            .I(N__16930));
    Odrv4 I__2893 (
            .O(N__16930),
            .I(\Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0 ));
    InMux I__2892 (
            .O(N__16927),
            .I(N__16924));
    LocalMux I__2891 (
            .O(N__16924),
            .I(\Commands_frame_decoder.state_1_ns_0_a4_0_3_2 ));
    CascadeMux I__2890 (
            .O(N__16921),
            .I(\Commands_frame_decoder.N_323_cascade_ ));
    CEMux I__2889 (
            .O(N__16918),
            .I(N__16915));
    LocalMux I__2888 (
            .O(N__16915),
            .I(N__16912));
    Span4Mux_h I__2887 (
            .O(N__16912),
            .I(N__16909));
    Odrv4 I__2886 (
            .O(N__16909),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__2885 (
            .O(N__16906),
            .I(N__16902));
    InMux I__2884 (
            .O(N__16905),
            .I(N__16899));
    LocalMux I__2883 (
            .O(N__16902),
            .I(\Commands_frame_decoder.state_1Z0Z_2 ));
    LocalMux I__2882 (
            .O(N__16899),
            .I(\Commands_frame_decoder.state_1Z0Z_2 ));
    InMux I__2881 (
            .O(N__16894),
            .I(N__16882));
    InMux I__2880 (
            .O(N__16893),
            .I(N__16882));
    InMux I__2879 (
            .O(N__16892),
            .I(N__16882));
    InMux I__2878 (
            .O(N__16891),
            .I(N__16882));
    LocalMux I__2877 (
            .O(N__16882),
            .I(N__16879));
    Span4Mux_h I__2876 (
            .O(N__16879),
            .I(N__16875));
    InMux I__2875 (
            .O(N__16878),
            .I(N__16872));
    Odrv4 I__2874 (
            .O(N__16875),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    LocalMux I__2873 (
            .O(N__16872),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    CascadeMux I__2872 (
            .O(N__16867),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ));
    InMux I__2871 (
            .O(N__16864),
            .I(N__16858));
    InMux I__2870 (
            .O(N__16863),
            .I(N__16858));
    LocalMux I__2869 (
            .O(N__16858),
            .I(\Commands_frame_decoder.state_1Z0Z_3 ));
    CascadeMux I__2868 (
            .O(N__16855),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ));
    InMux I__2867 (
            .O(N__16852),
            .I(N__16848));
    InMux I__2866 (
            .O(N__16851),
            .I(N__16845));
    LocalMux I__2865 (
            .O(N__16848),
            .I(N__16842));
    LocalMux I__2864 (
            .O(N__16845),
            .I(\Commands_frame_decoder.state_1Z0Z_4 ));
    Odrv12 I__2863 (
            .O(N__16842),
            .I(\Commands_frame_decoder.state_1Z0Z_4 ));
    InMux I__2862 (
            .O(N__16837),
            .I(N__16833));
    InMux I__2861 (
            .O(N__16836),
            .I(N__16830));
    LocalMux I__2860 (
            .O(N__16833),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__2859 (
            .O(N__16830),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__2858 (
            .O(N__16825),
            .I(N__16821));
    InMux I__2857 (
            .O(N__16824),
            .I(N__16818));
    LocalMux I__2856 (
            .O(N__16821),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__2855 (
            .O(N__16818),
            .I(\reset_module_System.countZ0Z_3 ));
    CascadeMux I__2854 (
            .O(N__16813),
            .I(N__16810));
    InMux I__2853 (
            .O(N__16810),
            .I(N__16806));
    InMux I__2852 (
            .O(N__16809),
            .I(N__16803));
    LocalMux I__2851 (
            .O(N__16806),
            .I(N__16800));
    LocalMux I__2850 (
            .O(N__16803),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__2849 (
            .O(N__16800),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__2848 (
            .O(N__16795),
            .I(N__16791));
    InMux I__2847 (
            .O(N__16794),
            .I(N__16788));
    LocalMux I__2846 (
            .O(N__16791),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__2845 (
            .O(N__16788),
            .I(\reset_module_System.countZ0Z_2 ));
    CascadeMux I__2844 (
            .O(N__16783),
            .I(N__16778));
    InMux I__2843 (
            .O(N__16782),
            .I(N__16774));
    InMux I__2842 (
            .O(N__16781),
            .I(N__16771));
    InMux I__2841 (
            .O(N__16778),
            .I(N__16766));
    InMux I__2840 (
            .O(N__16777),
            .I(N__16766));
    LocalMux I__2839 (
            .O(N__16774),
            .I(N__16761));
    LocalMux I__2838 (
            .O(N__16771),
            .I(N__16761));
    LocalMux I__2837 (
            .O(N__16766),
            .I(\reset_module_System.reset6_15 ));
    Odrv4 I__2836 (
            .O(N__16761),
            .I(\reset_module_System.reset6_15 ));
    InMux I__2835 (
            .O(N__16756),
            .I(N__16753));
    LocalMux I__2834 (
            .O(N__16753),
            .I(N__16749));
    InMux I__2833 (
            .O(N__16752),
            .I(N__16746));
    Odrv4 I__2832 (
            .O(N__16749),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__2831 (
            .O(N__16746),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__2830 (
            .O(N__16741),
            .I(N__16737));
    InMux I__2829 (
            .O(N__16740),
            .I(N__16734));
    LocalMux I__2828 (
            .O(N__16737),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__2827 (
            .O(N__16734),
            .I(\reset_module_System.countZ0Z_10 ));
    CascadeMux I__2826 (
            .O(N__16729),
            .I(N__16726));
    InMux I__2825 (
            .O(N__16726),
            .I(N__16722));
    InMux I__2824 (
            .O(N__16725),
            .I(N__16719));
    LocalMux I__2823 (
            .O(N__16722),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__2822 (
            .O(N__16719),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__2821 (
            .O(N__16714),
            .I(N__16710));
    InMux I__2820 (
            .O(N__16713),
            .I(N__16707));
    LocalMux I__2819 (
            .O(N__16710),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__2818 (
            .O(N__16707),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__2817 (
            .O(N__16702),
            .I(N__16696));
    InMux I__2816 (
            .O(N__16701),
            .I(N__16691));
    InMux I__2815 (
            .O(N__16700),
            .I(N__16691));
    InMux I__2814 (
            .O(N__16699),
            .I(N__16688));
    LocalMux I__2813 (
            .O(N__16696),
            .I(N__16681));
    LocalMux I__2812 (
            .O(N__16691),
            .I(N__16681));
    LocalMux I__2811 (
            .O(N__16688),
            .I(N__16681));
    Odrv4 I__2810 (
            .O(N__16681),
            .I(\reset_module_System.reset6_14 ));
    CascadeMux I__2809 (
            .O(N__16678),
            .I(N__16673));
    CascadeMux I__2808 (
            .O(N__16677),
            .I(N__16669));
    CascadeMux I__2807 (
            .O(N__16676),
            .I(N__16666));
    InMux I__2806 (
            .O(N__16673),
            .I(N__16654));
    InMux I__2805 (
            .O(N__16672),
            .I(N__16654));
    InMux I__2804 (
            .O(N__16669),
            .I(N__16654));
    InMux I__2803 (
            .O(N__16666),
            .I(N__16654));
    InMux I__2802 (
            .O(N__16665),
            .I(N__16651));
    InMux I__2801 (
            .O(N__16664),
            .I(N__16646));
    InMux I__2800 (
            .O(N__16663),
            .I(N__16646));
    LocalMux I__2799 (
            .O(N__16654),
            .I(N__16639));
    LocalMux I__2798 (
            .O(N__16651),
            .I(N__16639));
    LocalMux I__2797 (
            .O(N__16646),
            .I(N__16639));
    Span4Mux_v I__2796 (
            .O(N__16639),
            .I(N__16636));
    Odrv4 I__2795 (
            .O(N__16636),
            .I(\Commands_frame_decoder.state_1_RNIVM1OZ0Z_6 ));
    CascadeMux I__2794 (
            .O(N__16633),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    InMux I__2793 (
            .O(N__16630),
            .I(N__16627));
    LocalMux I__2792 (
            .O(N__16627),
            .I(N__16624));
    Span4Mux_v I__2791 (
            .O(N__16624),
            .I(N__16620));
    InMux I__2790 (
            .O(N__16623),
            .I(N__16617));
    Span4Mux_h I__2789 (
            .O(N__16620),
            .I(N__16614));
    LocalMux I__2788 (
            .O(N__16617),
            .I(alt_kp_4));
    Odrv4 I__2787 (
            .O(N__16614),
            .I(alt_kp_4));
    InMux I__2786 (
            .O(N__16609),
            .I(N__16606));
    LocalMux I__2785 (
            .O(N__16606),
            .I(N__16603));
    Odrv4 I__2784 (
            .O(N__16603),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__2783 (
            .O(N__16600),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__2782 (
            .O(N__16597),
            .I(N__16592));
    InMux I__2781 (
            .O(N__16596),
            .I(N__16589));
    InMux I__2780 (
            .O(N__16595),
            .I(N__16586));
    LocalMux I__2779 (
            .O(N__16592),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__2778 (
            .O(N__16589),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__2777 (
            .O(N__16586),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__2776 (
            .O(N__16579),
            .I(N__16576));
    InMux I__2775 (
            .O(N__16576),
            .I(N__16573));
    LocalMux I__2774 (
            .O(N__16573),
            .I(N__16570));
    Odrv4 I__2773 (
            .O(N__16570),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__2772 (
            .O(N__16567),
            .I(N__16564));
    LocalMux I__2771 (
            .O(N__16564),
            .I(N__16561));
    Span4Mux_h I__2770 (
            .O(N__16561),
            .I(N__16558));
    Odrv4 I__2769 (
            .O(N__16558),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__2768 (
            .O(N__16555),
            .I(N__16552));
    LocalMux I__2767 (
            .O(N__16552),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    CascadeMux I__2766 (
            .O(N__16549),
            .I(N__16546));
    InMux I__2765 (
            .O(N__16546),
            .I(N__16543));
    LocalMux I__2764 (
            .O(N__16543),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__2763 (
            .O(N__16540),
            .I(N__16537));
    LocalMux I__2762 (
            .O(N__16537),
            .I(N__16534));
    Odrv12 I__2761 (
            .O(N__16534),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__2760 (
            .O(N__16531),
            .I(N__16528));
    LocalMux I__2759 (
            .O(N__16528),
            .I(N__16525));
    Odrv4 I__2758 (
            .O(N__16525),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    InMux I__2757 (
            .O(N__16522),
            .I(N__16519));
    LocalMux I__2756 (
            .O(N__16519),
            .I(N__16516));
    Span4Mux_v I__2755 (
            .O(N__16516),
            .I(N__16513));
    Odrv4 I__2754 (
            .O(N__16513),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__2753 (
            .O(N__16510),
            .I(N__16507));
    LocalMux I__2752 (
            .O(N__16507),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__2751 (
            .O(N__16504),
            .I(N__16501));
    LocalMux I__2750 (
            .O(N__16501),
            .I(N__16498));
    Span4Mux_v I__2749 (
            .O(N__16498),
            .I(N__16495));
    Odrv4 I__2748 (
            .O(N__16495),
            .I(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ));
    CascadeMux I__2747 (
            .O(N__16492),
            .I(N__16489));
    InMux I__2746 (
            .O(N__16489),
            .I(N__16486));
    LocalMux I__2745 (
            .O(N__16486),
            .I(N__16483));
    Span4Mux_h I__2744 (
            .O(N__16483),
            .I(N__16480));
    Odrv4 I__2743 (
            .O(N__16480),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__2742 (
            .O(N__16477),
            .I(N__16474));
    LocalMux I__2741 (
            .O(N__16474),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__2740 (
            .O(N__16471),
            .I(N__16468));
    LocalMux I__2739 (
            .O(N__16468),
            .I(N__16465));
    Span4Mux_s3_v I__2738 (
            .O(N__16465),
            .I(N__16462));
    Odrv4 I__2737 (
            .O(N__16462),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__2736 (
            .O(N__16459),
            .I(N__16452));
    InMux I__2735 (
            .O(N__16458),
            .I(N__16452));
    InMux I__2734 (
            .O(N__16457),
            .I(N__16449));
    LocalMux I__2733 (
            .O(N__16452),
            .I(N__16444));
    LocalMux I__2732 (
            .O(N__16449),
            .I(N__16437));
    InMux I__2731 (
            .O(N__16448),
            .I(N__16432));
    InMux I__2730 (
            .O(N__16447),
            .I(N__16432));
    Span4Mux_h I__2729 (
            .O(N__16444),
            .I(N__16429));
    InMux I__2728 (
            .O(N__16443),
            .I(N__16426));
    InMux I__2727 (
            .O(N__16442),
            .I(N__16419));
    InMux I__2726 (
            .O(N__16441),
            .I(N__16419));
    InMux I__2725 (
            .O(N__16440),
            .I(N__16419));
    Span4Mux_s3_v I__2724 (
            .O(N__16437),
            .I(N__16414));
    LocalMux I__2723 (
            .O(N__16432),
            .I(N__16414));
    Odrv4 I__2722 (
            .O(N__16429),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__2721 (
            .O(N__16426),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__2720 (
            .O(N__16419),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    Odrv4 I__2719 (
            .O(N__16414),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    InMux I__2718 (
            .O(N__16405),
            .I(N__16402));
    LocalMux I__2717 (
            .O(N__16402),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__2716 (
            .O(N__16399),
            .I(N__16396));
    LocalMux I__2715 (
            .O(N__16396),
            .I(N__16393));
    Span4Mux_h I__2714 (
            .O(N__16393),
            .I(N__16390));
    Odrv4 I__2713 (
            .O(N__16390),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__2712 (
            .O(N__16387),
            .I(N__16384));
    LocalMux I__2711 (
            .O(N__16384),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    CascadeMux I__2710 (
            .O(N__16381),
            .I(N__16378));
    InMux I__2709 (
            .O(N__16378),
            .I(N__16375));
    LocalMux I__2708 (
            .O(N__16375),
            .I(N__16372));
    Odrv4 I__2707 (
            .O(N__16372),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ));
    InMux I__2706 (
            .O(N__16369),
            .I(N__16366));
    LocalMux I__2705 (
            .O(N__16366),
            .I(N__16363));
    Span4Mux_h I__2704 (
            .O(N__16363),
            .I(N__16360));
    Odrv4 I__2703 (
            .O(N__16360),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__2702 (
            .O(N__16357),
            .I(N__16354));
    LocalMux I__2701 (
            .O(N__16354),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__2700 (
            .O(N__16351),
            .I(N__16348));
    LocalMux I__2699 (
            .O(N__16348),
            .I(N__16345));
    Span4Mux_h I__2698 (
            .O(N__16345),
            .I(N__16341));
    InMux I__2697 (
            .O(N__16344),
            .I(N__16338));
    Odrv4 I__2696 (
            .O(N__16341),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    LocalMux I__2695 (
            .O(N__16338),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    CascadeMux I__2694 (
            .O(N__16333),
            .I(N__16330));
    InMux I__2693 (
            .O(N__16330),
            .I(N__16327));
    LocalMux I__2692 (
            .O(N__16327),
            .I(N__16323));
    InMux I__2691 (
            .O(N__16326),
            .I(N__16320));
    Span4Mux_v I__2690 (
            .O(N__16323),
            .I(N__16314));
    LocalMux I__2689 (
            .O(N__16320),
            .I(N__16314));
    CascadeMux I__2688 (
            .O(N__16319),
            .I(N__16308));
    Span4Mux_h I__2687 (
            .O(N__16314),
            .I(N__16305));
    InMux I__2686 (
            .O(N__16313),
            .I(N__16302));
    InMux I__2685 (
            .O(N__16312),
            .I(N__16295));
    InMux I__2684 (
            .O(N__16311),
            .I(N__16295));
    InMux I__2683 (
            .O(N__16308),
            .I(N__16295));
    Odrv4 I__2682 (
            .O(N__16305),
            .I(\ppm_encoder_1.N_226 ));
    LocalMux I__2681 (
            .O(N__16302),
            .I(\ppm_encoder_1.N_226 ));
    LocalMux I__2680 (
            .O(N__16295),
            .I(\ppm_encoder_1.N_226 ));
    CascadeMux I__2679 (
            .O(N__16288),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ));
    InMux I__2678 (
            .O(N__16285),
            .I(N__16282));
    LocalMux I__2677 (
            .O(N__16282),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    CascadeMux I__2676 (
            .O(N__16279),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ));
    InMux I__2675 (
            .O(N__16276),
            .I(N__16273));
    LocalMux I__2674 (
            .O(N__16273),
            .I(N__16270));
    Span4Mux_h I__2673 (
            .O(N__16270),
            .I(N__16267));
    Odrv4 I__2672 (
            .O(N__16267),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__2671 (
            .O(N__16264),
            .I(N__16261));
    LocalMux I__2670 (
            .O(N__16261),
            .I(N__16257));
    InMux I__2669 (
            .O(N__16260),
            .I(N__16254));
    Span4Mux_v I__2668 (
            .O(N__16257),
            .I(N__16251));
    LocalMux I__2667 (
            .O(N__16254),
            .I(N__16248));
    Odrv4 I__2666 (
            .O(N__16251),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    Odrv4 I__2665 (
            .O(N__16248),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    InMux I__2664 (
            .O(N__16243),
            .I(N__16240));
    LocalMux I__2663 (
            .O(N__16240),
            .I(N__16235));
    InMux I__2662 (
            .O(N__16239),
            .I(N__16230));
    InMux I__2661 (
            .O(N__16238),
            .I(N__16230));
    Odrv4 I__2660 (
            .O(N__16235),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__2659 (
            .O(N__16230),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__2658 (
            .O(N__16225),
            .I(N__16222));
    LocalMux I__2657 (
            .O(N__16222),
            .I(N__16219));
    Span4Mux_h I__2656 (
            .O(N__16219),
            .I(N__16216));
    Odrv4 I__2655 (
            .O(N__16216),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__2654 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__2653 (
            .O(N__16210),
            .I(N__16207));
    Span4Mux_h I__2652 (
            .O(N__16207),
            .I(N__16204));
    Odrv4 I__2651 (
            .O(N__16204),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__2650 (
            .O(N__16201),
            .I(N__16198));
    LocalMux I__2649 (
            .O(N__16198),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__2648 (
            .O(N__16195),
            .I(N__16188));
    InMux I__2647 (
            .O(N__16194),
            .I(N__16188));
    CascadeMux I__2646 (
            .O(N__16193),
            .I(N__16185));
    LocalMux I__2645 (
            .O(N__16188),
            .I(N__16182));
    InMux I__2644 (
            .O(N__16185),
            .I(N__16179));
    Span4Mux_v I__2643 (
            .O(N__16182),
            .I(N__16176));
    LocalMux I__2642 (
            .O(N__16179),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__2641 (
            .O(N__16176),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    CascadeMux I__2640 (
            .O(N__16171),
            .I(N__16168));
    InMux I__2639 (
            .O(N__16168),
            .I(N__16165));
    LocalMux I__2638 (
            .O(N__16165),
            .I(N__16162));
    Span4Mux_h I__2637 (
            .O(N__16162),
            .I(N__16159));
    Odrv4 I__2636 (
            .O(N__16159),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__2635 (
            .O(N__16156),
            .I(N__16153));
    LocalMux I__2634 (
            .O(N__16153),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__2633 (
            .O(N__16150),
            .I(N__16145));
    InMux I__2632 (
            .O(N__16149),
            .I(N__16142));
    InMux I__2631 (
            .O(N__16148),
            .I(N__16139));
    LocalMux I__2630 (
            .O(N__16145),
            .I(N__16136));
    LocalMux I__2629 (
            .O(N__16142),
            .I(N__16133));
    LocalMux I__2628 (
            .O(N__16139),
            .I(N__16128));
    Span4Mux_h I__2627 (
            .O(N__16136),
            .I(N__16128));
    Odrv4 I__2626 (
            .O(N__16133),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    Odrv4 I__2625 (
            .O(N__16128),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__2624 (
            .O(N__16123),
            .I(N__16120));
    LocalMux I__2623 (
            .O(N__16120),
            .I(N__16117));
    Span4Mux_v I__2622 (
            .O(N__16117),
            .I(N__16114));
    Odrv4 I__2621 (
            .O(N__16114),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__2620 (
            .O(N__16111),
            .I(N__16108));
    LocalMux I__2619 (
            .O(N__16108),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__2618 (
            .O(N__16105),
            .I(N__16101));
    InMux I__2617 (
            .O(N__16104),
            .I(N__16098));
    LocalMux I__2616 (
            .O(N__16101),
            .I(N__16095));
    LocalMux I__2615 (
            .O(N__16098),
            .I(N__16092));
    Span4Mux_v I__2614 (
            .O(N__16095),
            .I(N__16089));
    Span4Mux_h I__2613 (
            .O(N__16092),
            .I(N__16086));
    Odrv4 I__2612 (
            .O(N__16089),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    Odrv4 I__2611 (
            .O(N__16086),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    CascadeMux I__2610 (
            .O(N__16081),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ));
    CascadeMux I__2609 (
            .O(N__16078),
            .I(N__16075));
    InMux I__2608 (
            .O(N__16075),
            .I(N__16072));
    LocalMux I__2607 (
            .O(N__16072),
            .I(N__16069));
    Odrv4 I__2606 (
            .O(N__16069),
            .I(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ));
    CascadeMux I__2605 (
            .O(N__16066),
            .I(N__16062));
    CascadeMux I__2604 (
            .O(N__16065),
            .I(N__16057));
    InMux I__2603 (
            .O(N__16062),
            .I(N__16047));
    InMux I__2602 (
            .O(N__16061),
            .I(N__16047));
    InMux I__2601 (
            .O(N__16060),
            .I(N__16047));
    InMux I__2600 (
            .O(N__16057),
            .I(N__16044));
    CascadeMux I__2599 (
            .O(N__16056),
            .I(N__16038));
    CascadeMux I__2598 (
            .O(N__16055),
            .I(N__16035));
    CascadeMux I__2597 (
            .O(N__16054),
            .I(N__16032));
    LocalMux I__2596 (
            .O(N__16047),
            .I(N__16028));
    LocalMux I__2595 (
            .O(N__16044),
            .I(N__16025));
    InMux I__2594 (
            .O(N__16043),
            .I(N__16020));
    InMux I__2593 (
            .O(N__16042),
            .I(N__16020));
    InMux I__2592 (
            .O(N__16041),
            .I(N__16015));
    InMux I__2591 (
            .O(N__16038),
            .I(N__16015));
    InMux I__2590 (
            .O(N__16035),
            .I(N__16012));
    InMux I__2589 (
            .O(N__16032),
            .I(N__16007));
    InMux I__2588 (
            .O(N__16031),
            .I(N__16007));
    Odrv4 I__2587 (
            .O(N__16028),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__2586 (
            .O(N__16025),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__2585 (
            .O(N__16020),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__2584 (
            .O(N__16015),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__2583 (
            .O(N__16012),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__2582 (
            .O(N__16007),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    InMux I__2581 (
            .O(N__15994),
            .I(N__15981));
    InMux I__2580 (
            .O(N__15993),
            .I(N__15981));
    InMux I__2579 (
            .O(N__15992),
            .I(N__15981));
    InMux I__2578 (
            .O(N__15991),
            .I(N__15978));
    CascadeMux I__2577 (
            .O(N__15990),
            .I(N__15974));
    CascadeMux I__2576 (
            .O(N__15989),
            .I(N__15971));
    CascadeMux I__2575 (
            .O(N__15988),
            .I(N__15966));
    LocalMux I__2574 (
            .O(N__15981),
            .I(N__15961));
    LocalMux I__2573 (
            .O(N__15978),
            .I(N__15958));
    InMux I__2572 (
            .O(N__15977),
            .I(N__15955));
    InMux I__2571 (
            .O(N__15974),
            .I(N__15950));
    InMux I__2570 (
            .O(N__15971),
            .I(N__15950));
    InMux I__2569 (
            .O(N__15970),
            .I(N__15947));
    InMux I__2568 (
            .O(N__15969),
            .I(N__15942));
    InMux I__2567 (
            .O(N__15966),
            .I(N__15942));
    InMux I__2566 (
            .O(N__15965),
            .I(N__15937));
    InMux I__2565 (
            .O(N__15964),
            .I(N__15937));
    Odrv4 I__2564 (
            .O(N__15961),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__2563 (
            .O(N__15958),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__2562 (
            .O(N__15955),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__2561 (
            .O(N__15950),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__2560 (
            .O(N__15947),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__2559 (
            .O(N__15942),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__2558 (
            .O(N__15937),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__2557 (
            .O(N__15922),
            .I(N__15919));
    LocalMux I__2556 (
            .O(N__15919),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    CascadeMux I__2555 (
            .O(N__15916),
            .I(N__15913));
    InMux I__2554 (
            .O(N__15913),
            .I(N__15910));
    LocalMux I__2553 (
            .O(N__15910),
            .I(N__15906));
    CascadeMux I__2552 (
            .O(N__15909),
            .I(N__15903));
    Span4Mux_v I__2551 (
            .O(N__15906),
            .I(N__15898));
    InMux I__2550 (
            .O(N__15903),
            .I(N__15895));
    InMux I__2549 (
            .O(N__15902),
            .I(N__15890));
    InMux I__2548 (
            .O(N__15901),
            .I(N__15890));
    Odrv4 I__2547 (
            .O(N__15898),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__2546 (
            .O(N__15895),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__2545 (
            .O(N__15890),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    CascadeMux I__2544 (
            .O(N__15883),
            .I(N__15878));
    CascadeMux I__2543 (
            .O(N__15882),
            .I(N__15875));
    CascadeMux I__2542 (
            .O(N__15881),
            .I(N__15872));
    InMux I__2541 (
            .O(N__15878),
            .I(N__15869));
    InMux I__2540 (
            .O(N__15875),
            .I(N__15866));
    InMux I__2539 (
            .O(N__15872),
            .I(N__15859));
    LocalMux I__2538 (
            .O(N__15869),
            .I(N__15856));
    LocalMux I__2537 (
            .O(N__15866),
            .I(N__15853));
    CascadeMux I__2536 (
            .O(N__15865),
            .I(N__15841));
    InMux I__2535 (
            .O(N__15864),
            .I(N__15838));
    InMux I__2534 (
            .O(N__15863),
            .I(N__15833));
    InMux I__2533 (
            .O(N__15862),
            .I(N__15833));
    LocalMux I__2532 (
            .O(N__15859),
            .I(N__15830));
    Span4Mux_h I__2531 (
            .O(N__15856),
            .I(N__15825));
    Span4Mux_v I__2530 (
            .O(N__15853),
            .I(N__15825));
    InMux I__2529 (
            .O(N__15852),
            .I(N__15818));
    InMux I__2528 (
            .O(N__15851),
            .I(N__15818));
    InMux I__2527 (
            .O(N__15850),
            .I(N__15818));
    InMux I__2526 (
            .O(N__15849),
            .I(N__15815));
    InMux I__2525 (
            .O(N__15848),
            .I(N__15812));
    InMux I__2524 (
            .O(N__15847),
            .I(N__15809));
    InMux I__2523 (
            .O(N__15846),
            .I(N__15806));
    InMux I__2522 (
            .O(N__15845),
            .I(N__15801));
    InMux I__2521 (
            .O(N__15844),
            .I(N__15801));
    InMux I__2520 (
            .O(N__15841),
            .I(N__15798));
    LocalMux I__2519 (
            .O(N__15838),
            .I(N__15793));
    LocalMux I__2518 (
            .O(N__15833),
            .I(N__15793));
    Odrv4 I__2517 (
            .O(N__15830),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__2516 (
            .O(N__15825),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2515 (
            .O(N__15818),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2514 (
            .O(N__15815),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2513 (
            .O(N__15812),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2512 (
            .O(N__15809),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2511 (
            .O(N__15806),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2510 (
            .O(N__15801),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__2509 (
            .O(N__15798),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__2508 (
            .O(N__15793),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    CascadeMux I__2507 (
            .O(N__15772),
            .I(N__15766));
    CascadeMux I__2506 (
            .O(N__15771),
            .I(N__15762));
    InMux I__2505 (
            .O(N__15770),
            .I(N__15758));
    InMux I__2504 (
            .O(N__15769),
            .I(N__15754));
    InMux I__2503 (
            .O(N__15766),
            .I(N__15747));
    InMux I__2502 (
            .O(N__15765),
            .I(N__15747));
    InMux I__2501 (
            .O(N__15762),
            .I(N__15747));
    InMux I__2500 (
            .O(N__15761),
            .I(N__15742));
    LocalMux I__2499 (
            .O(N__15758),
            .I(N__15739));
    CascadeMux I__2498 (
            .O(N__15757),
            .I(N__15736));
    LocalMux I__2497 (
            .O(N__15754),
            .I(N__15733));
    LocalMux I__2496 (
            .O(N__15747),
            .I(N__15730));
    InMux I__2495 (
            .O(N__15746),
            .I(N__15727));
    CascadeMux I__2494 (
            .O(N__15745),
            .I(N__15723));
    LocalMux I__2493 (
            .O(N__15742),
            .I(N__15720));
    Span4Mux_h I__2492 (
            .O(N__15739),
            .I(N__15717));
    InMux I__2491 (
            .O(N__15736),
            .I(N__15714));
    Span4Mux_v I__2490 (
            .O(N__15733),
            .I(N__15709));
    Span4Mux_h I__2489 (
            .O(N__15730),
            .I(N__15709));
    LocalMux I__2488 (
            .O(N__15727),
            .I(N__15706));
    InMux I__2487 (
            .O(N__15726),
            .I(N__15701));
    InMux I__2486 (
            .O(N__15723),
            .I(N__15701));
    Odrv4 I__2485 (
            .O(N__15720),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__2484 (
            .O(N__15717),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__2483 (
            .O(N__15714),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__2482 (
            .O(N__15709),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__2481 (
            .O(N__15706),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__2480 (
            .O(N__15701),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    InMux I__2479 (
            .O(N__15688),
            .I(N__15684));
    InMux I__2478 (
            .O(N__15687),
            .I(N__15681));
    LocalMux I__2477 (
            .O(N__15684),
            .I(N__15676));
    LocalMux I__2476 (
            .O(N__15681),
            .I(N__15676));
    Span4Mux_v I__2475 (
            .O(N__15676),
            .I(N__15673));
    Odrv4 I__2474 (
            .O(N__15673),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    CascadeMux I__2473 (
            .O(N__15670),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ));
    InMux I__2472 (
            .O(N__15667),
            .I(N__15664));
    LocalMux I__2471 (
            .O(N__15664),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10 ));
    CascadeMux I__2470 (
            .O(N__15661),
            .I(N__15658));
    InMux I__2469 (
            .O(N__15658),
            .I(N__15655));
    LocalMux I__2468 (
            .O(N__15655),
            .I(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ));
    InMux I__2467 (
            .O(N__15652),
            .I(N__15649));
    LocalMux I__2466 (
            .O(N__15649),
            .I(\ppm_encoder_1.N_318 ));
    CascadeMux I__2465 (
            .O(N__15646),
            .I(\ppm_encoder_1.N_300_cascade_ ));
    InMux I__2464 (
            .O(N__15643),
            .I(N__15640));
    LocalMux I__2463 (
            .O(N__15640),
            .I(N__15637));
    Span4Mux_v I__2462 (
            .O(N__15637),
            .I(N__15634));
    Odrv4 I__2461 (
            .O(N__15634),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ));
    InMux I__2460 (
            .O(N__15631),
            .I(N__15628));
    LocalMux I__2459 (
            .O(N__15628),
            .I(\ppm_encoder_1.N_139_0 ));
    CascadeMux I__2458 (
            .O(N__15625),
            .I(N__15622));
    InMux I__2457 (
            .O(N__15622),
            .I(N__15619));
    LocalMux I__2456 (
            .O(N__15619),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14 ));
    CascadeMux I__2455 (
            .O(N__15616),
            .I(N__15613));
    InMux I__2454 (
            .O(N__15613),
            .I(N__15610));
    LocalMux I__2453 (
            .O(N__15610),
            .I(N__15607));
    Odrv4 I__2452 (
            .O(N__15607),
            .I(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ));
    InMux I__2451 (
            .O(N__15604),
            .I(N__15601));
    LocalMux I__2450 (
            .O(N__15601),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    InMux I__2449 (
            .O(N__15598),
            .I(N__15593));
    InMux I__2448 (
            .O(N__15597),
            .I(N__15588));
    InMux I__2447 (
            .O(N__15596),
            .I(N__15588));
    LocalMux I__2446 (
            .O(N__15593),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__2445 (
            .O(N__15588),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__2444 (
            .O(N__15583),
            .I(N__15579));
    InMux I__2443 (
            .O(N__15582),
            .I(N__15576));
    LocalMux I__2442 (
            .O(N__15579),
            .I(N__15573));
    LocalMux I__2441 (
            .O(N__15576),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    Odrv4 I__2440 (
            .O(N__15573),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__2439 (
            .O(N__15568),
            .I(N__15563));
    InMux I__2438 (
            .O(N__15567),
            .I(N__15558));
    InMux I__2437 (
            .O(N__15566),
            .I(N__15558));
    LocalMux I__2436 (
            .O(N__15563),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__2435 (
            .O(N__15558),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__2434 (
            .O(N__15553),
            .I(N__15549));
    InMux I__2433 (
            .O(N__15552),
            .I(N__15546));
    LocalMux I__2432 (
            .O(N__15549),
            .I(N__15543));
    LocalMux I__2431 (
            .O(N__15546),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    Odrv4 I__2430 (
            .O(N__15543),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__2429 (
            .O(N__15538),
            .I(N__15535));
    LocalMux I__2428 (
            .O(N__15535),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    CascadeMux I__2427 (
            .O(N__15532),
            .I(\Commands_frame_decoder.WDT8lto13_1_cascade_ ));
    InMux I__2426 (
            .O(N__15529),
            .I(N__15526));
    LocalMux I__2425 (
            .O(N__15526),
            .I(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ));
    IoInMux I__2424 (
            .O(N__15523),
            .I(N__15520));
    LocalMux I__2423 (
            .O(N__15520),
            .I(N__15517));
    Span4Mux_s2_v I__2422 (
            .O(N__15517),
            .I(N__15514));
    Span4Mux_v I__2421 (
            .O(N__15514),
            .I(N__15511));
    Sp12to4 I__2420 (
            .O(N__15511),
            .I(N__15508));
    Span12Mux_h I__2419 (
            .O(N__15508),
            .I(N__15504));
    CascadeMux I__2418 (
            .O(N__15507),
            .I(N__15501));
    Span12Mux_v I__2417 (
            .O(N__15504),
            .I(N__15498));
    InMux I__2416 (
            .O(N__15501),
            .I(N__15495));
    Odrv12 I__2415 (
            .O(N__15498),
            .I(ppm_output_c));
    LocalMux I__2414 (
            .O(N__15495),
            .I(ppm_output_c));
    InMux I__2413 (
            .O(N__15490),
            .I(N__15487));
    LocalMux I__2412 (
            .O(N__15487),
            .I(N__15484));
    Span4Mux_s1_v I__2411 (
            .O(N__15484),
            .I(N__15480));
    InMux I__2410 (
            .O(N__15483),
            .I(N__15476));
    Span4Mux_v I__2409 (
            .O(N__15480),
            .I(N__15473));
    InMux I__2408 (
            .O(N__15479),
            .I(N__15470));
    LocalMux I__2407 (
            .O(N__15476),
            .I(N__15465));
    Span4Mux_v I__2406 (
            .O(N__15473),
            .I(N__15465));
    LocalMux I__2405 (
            .O(N__15470),
            .I(N__15462));
    Odrv4 I__2404 (
            .O(N__15465),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    Odrv4 I__2403 (
            .O(N__15462),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    InMux I__2402 (
            .O(N__15457),
            .I(N__15452));
    InMux I__2401 (
            .O(N__15456),
            .I(N__15449));
    InMux I__2400 (
            .O(N__15455),
            .I(N__15446));
    LocalMux I__2399 (
            .O(N__15452),
            .I(N__15443));
    LocalMux I__2398 (
            .O(N__15449),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    LocalMux I__2397 (
            .O(N__15446),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__2396 (
            .O(N__15443),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__2395 (
            .O(N__15436),
            .I(N__15432));
    InMux I__2394 (
            .O(N__15435),
            .I(N__15429));
    LocalMux I__2393 (
            .O(N__15432),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__2392 (
            .O(N__15429),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__2391 (
            .O(N__15424),
            .I(bfn_4_19_0_));
    CascadeMux I__2390 (
            .O(N__15421),
            .I(N__15417));
    InMux I__2389 (
            .O(N__15420),
            .I(N__15414));
    InMux I__2388 (
            .O(N__15417),
            .I(N__15411));
    LocalMux I__2387 (
            .O(N__15414),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__2386 (
            .O(N__15411),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__2385 (
            .O(N__15406),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__2384 (
            .O(N__15403),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__2383 (
            .O(N__15400),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__2382 (
            .O(N__15397),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__2381 (
            .O(N__15394),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__2380 (
            .O(N__15391),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__2379 (
            .O(N__15388),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    CascadeMux I__2378 (
            .O(N__15385),
            .I(N__15381));
    InMux I__2377 (
            .O(N__15384),
            .I(N__15378));
    InMux I__2376 (
            .O(N__15381),
            .I(N__15375));
    LocalMux I__2375 (
            .O(N__15378),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__2374 (
            .O(N__15375),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__2373 (
            .O(N__15370),
            .I(N__15366));
    InMux I__2372 (
            .O(N__15369),
            .I(N__15363));
    LocalMux I__2371 (
            .O(N__15366),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__2370 (
            .O(N__15363),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__2369 (
            .O(N__15358),
            .I(N__15355));
    LocalMux I__2368 (
            .O(N__15355),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__2367 (
            .O(N__15352),
            .I(N__15349));
    LocalMux I__2366 (
            .O(N__15349),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__2365 (
            .O(N__15346),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__2364 (
            .O(N__15343),
            .I(N__15340));
    LocalMux I__2363 (
            .O(N__15340),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__2362 (
            .O(N__15337),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__2361 (
            .O(N__15334),
            .I(N__15331));
    LocalMux I__2360 (
            .O(N__15331),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__2359 (
            .O(N__15328),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__2358 (
            .O(N__15325),
            .I(N__15321));
    InMux I__2357 (
            .O(N__15324),
            .I(N__15318));
    LocalMux I__2356 (
            .O(N__15321),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__2355 (
            .O(N__15318),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__2354 (
            .O(N__15313),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__2353 (
            .O(N__15310),
            .I(N__15306));
    InMux I__2352 (
            .O(N__15309),
            .I(N__15303));
    LocalMux I__2351 (
            .O(N__15306),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__2350 (
            .O(N__15303),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    InMux I__2349 (
            .O(N__15298),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__2348 (
            .O(N__15295),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__2347 (
            .O(N__15292),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__2346 (
            .O(N__15289),
            .I(N__15284));
    InMux I__2345 (
            .O(N__15288),
            .I(N__15278));
    InMux I__2344 (
            .O(N__15287),
            .I(N__15278));
    LocalMux I__2343 (
            .O(N__15284),
            .I(N__15275));
    InMux I__2342 (
            .O(N__15283),
            .I(N__15272));
    LocalMux I__2341 (
            .O(N__15278),
            .I(N__15269));
    Span4Mux_h I__2340 (
            .O(N__15275),
            .I(N__15264));
    LocalMux I__2339 (
            .O(N__15272),
            .I(N__15264));
    Span4Mux_h I__2338 (
            .O(N__15269),
            .I(N__15261));
    Odrv4 I__2337 (
            .O(N__15264),
            .I(uart_drone_data_2));
    Odrv4 I__2336 (
            .O(N__15261),
            .I(uart_drone_data_2));
    InMux I__2335 (
            .O(N__15256),
            .I(N__15249));
    InMux I__2334 (
            .O(N__15255),
            .I(N__15244));
    InMux I__2333 (
            .O(N__15254),
            .I(N__15244));
    InMux I__2332 (
            .O(N__15253),
            .I(N__15241));
    InMux I__2331 (
            .O(N__15252),
            .I(N__15238));
    LocalMux I__2330 (
            .O(N__15249),
            .I(N__15235));
    LocalMux I__2329 (
            .O(N__15244),
            .I(N__15230));
    LocalMux I__2328 (
            .O(N__15241),
            .I(N__15225));
    LocalMux I__2327 (
            .O(N__15238),
            .I(N__15225));
    Span4Mux_h I__2326 (
            .O(N__15235),
            .I(N__15222));
    InMux I__2325 (
            .O(N__15234),
            .I(N__15219));
    InMux I__2324 (
            .O(N__15233),
            .I(N__15216));
    Span4Mux_h I__2323 (
            .O(N__15230),
            .I(N__15213));
    Span4Mux_h I__2322 (
            .O(N__15225),
            .I(N__15210));
    Odrv4 I__2321 (
            .O(N__15222),
            .I(uart_drone_data_3));
    LocalMux I__2320 (
            .O(N__15219),
            .I(uart_drone_data_3));
    LocalMux I__2319 (
            .O(N__15216),
            .I(uart_drone_data_3));
    Odrv4 I__2318 (
            .O(N__15213),
            .I(uart_drone_data_3));
    Odrv4 I__2317 (
            .O(N__15210),
            .I(uart_drone_data_3));
    CascadeMux I__2316 (
            .O(N__15199),
            .I(N__15196));
    InMux I__2315 (
            .O(N__15196),
            .I(N__15193));
    LocalMux I__2314 (
            .O(N__15193),
            .I(N__15186));
    InMux I__2313 (
            .O(N__15192),
            .I(N__15183));
    InMux I__2312 (
            .O(N__15191),
            .I(N__15180));
    InMux I__2311 (
            .O(N__15190),
            .I(N__15175));
    InMux I__2310 (
            .O(N__15189),
            .I(N__15175));
    Span4Mux_v I__2309 (
            .O(N__15186),
            .I(N__15170));
    LocalMux I__2308 (
            .O(N__15183),
            .I(N__15170));
    LocalMux I__2307 (
            .O(N__15180),
            .I(N__15166));
    LocalMux I__2306 (
            .O(N__15175),
            .I(N__15162));
    Span4Mux_v I__2305 (
            .O(N__15170),
            .I(N__15159));
    InMux I__2304 (
            .O(N__15169),
            .I(N__15156));
    Span4Mux_h I__2303 (
            .O(N__15166),
            .I(N__15153));
    InMux I__2302 (
            .O(N__15165),
            .I(N__15150));
    Span4Mux_h I__2301 (
            .O(N__15162),
            .I(N__15147));
    Odrv4 I__2300 (
            .O(N__15159),
            .I(uart_drone_data_4));
    LocalMux I__2299 (
            .O(N__15156),
            .I(uart_drone_data_4));
    Odrv4 I__2298 (
            .O(N__15153),
            .I(uart_drone_data_4));
    LocalMux I__2297 (
            .O(N__15150),
            .I(uart_drone_data_4));
    Odrv4 I__2296 (
            .O(N__15147),
            .I(uart_drone_data_4));
    CascadeMux I__2295 (
            .O(N__15136),
            .I(N__15133));
    InMux I__2294 (
            .O(N__15133),
            .I(N__15129));
    InMux I__2293 (
            .O(N__15132),
            .I(N__15126));
    LocalMux I__2292 (
            .O(N__15129),
            .I(N__15122));
    LocalMux I__2291 (
            .O(N__15126),
            .I(N__15119));
    InMux I__2290 (
            .O(N__15125),
            .I(N__15116));
    Span4Mux_h I__2289 (
            .O(N__15122),
            .I(N__15113));
    Span4Mux_v I__2288 (
            .O(N__15119),
            .I(N__15108));
    LocalMux I__2287 (
            .O(N__15116),
            .I(N__15108));
    Span4Mux_h I__2286 (
            .O(N__15113),
            .I(N__15104));
    Span4Mux_h I__2285 (
            .O(N__15108),
            .I(N__15101));
    InMux I__2284 (
            .O(N__15107),
            .I(N__15098));
    Odrv4 I__2283 (
            .O(N__15104),
            .I(uart_drone_data_5));
    Odrv4 I__2282 (
            .O(N__15101),
            .I(uart_drone_data_5));
    LocalMux I__2281 (
            .O(N__15098),
            .I(uart_drone_data_5));
    InMux I__2280 (
            .O(N__15091),
            .I(N__15079));
    InMux I__2279 (
            .O(N__15090),
            .I(N__15070));
    InMux I__2278 (
            .O(N__15089),
            .I(N__15070));
    InMux I__2277 (
            .O(N__15088),
            .I(N__15070));
    InMux I__2276 (
            .O(N__15087),
            .I(N__15070));
    InMux I__2275 (
            .O(N__15086),
            .I(N__15067));
    InMux I__2274 (
            .O(N__15085),
            .I(N__15062));
    InMux I__2273 (
            .O(N__15084),
            .I(N__15062));
    InMux I__2272 (
            .O(N__15083),
            .I(N__15057));
    InMux I__2271 (
            .O(N__15082),
            .I(N__15057));
    LocalMux I__2270 (
            .O(N__15079),
            .I(N__15054));
    LocalMux I__2269 (
            .O(N__15070),
            .I(N__15051));
    LocalMux I__2268 (
            .O(N__15067),
            .I(N__15044));
    LocalMux I__2267 (
            .O(N__15062),
            .I(N__15044));
    LocalMux I__2266 (
            .O(N__15057),
            .I(N__15041));
    Span4Mux_h I__2265 (
            .O(N__15054),
            .I(N__15036));
    Span4Mux_h I__2264 (
            .O(N__15051),
            .I(N__15036));
    InMux I__2263 (
            .O(N__15050),
            .I(N__15033));
    InMux I__2262 (
            .O(N__15049),
            .I(N__15030));
    Span4Mux_h I__2261 (
            .O(N__15044),
            .I(N__15025));
    Span4Mux_v I__2260 (
            .O(N__15041),
            .I(N__15025));
    Odrv4 I__2259 (
            .O(N__15036),
            .I(uart_drone_data_6));
    LocalMux I__2258 (
            .O(N__15033),
            .I(uart_drone_data_6));
    LocalMux I__2257 (
            .O(N__15030),
            .I(uart_drone_data_6));
    Odrv4 I__2256 (
            .O(N__15025),
            .I(uart_drone_data_6));
    CascadeMux I__2255 (
            .O(N__15016),
            .I(N__15008));
    InMux I__2254 (
            .O(N__15015),
            .I(N__15003));
    InMux I__2253 (
            .O(N__15014),
            .I(N__15000));
    InMux I__2252 (
            .O(N__15013),
            .I(N__14993));
    InMux I__2251 (
            .O(N__15012),
            .I(N__14993));
    InMux I__2250 (
            .O(N__15011),
            .I(N__14993));
    InMux I__2249 (
            .O(N__15008),
            .I(N__14990));
    InMux I__2248 (
            .O(N__15007),
            .I(N__14985));
    InMux I__2247 (
            .O(N__15006),
            .I(N__14985));
    LocalMux I__2246 (
            .O(N__15003),
            .I(N__14980));
    LocalMux I__2245 (
            .O(N__15000),
            .I(N__14980));
    LocalMux I__2244 (
            .O(N__14993),
            .I(N__14977));
    LocalMux I__2243 (
            .O(N__14990),
            .I(N__14972));
    LocalMux I__2242 (
            .O(N__14985),
            .I(N__14972));
    Span4Mux_v I__2241 (
            .O(N__14980),
            .I(N__14968));
    Span4Mux_h I__2240 (
            .O(N__14977),
            .I(N__14965));
    Span4Mux_h I__2239 (
            .O(N__14972),
            .I(N__14962));
    InMux I__2238 (
            .O(N__14971),
            .I(N__14959));
    Odrv4 I__2237 (
            .O(N__14968),
            .I(uart_drone_data_7));
    Odrv4 I__2236 (
            .O(N__14965),
            .I(uart_drone_data_7));
    Odrv4 I__2235 (
            .O(N__14962),
            .I(uart_drone_data_7));
    LocalMux I__2234 (
            .O(N__14959),
            .I(uart_drone_data_7));
    CEMux I__2233 (
            .O(N__14950),
            .I(N__14947));
    LocalMux I__2232 (
            .O(N__14947),
            .I(\uart_drone.state_1_sqmuxa_0 ));
    SRMux I__2231 (
            .O(N__14944),
            .I(N__14941));
    LocalMux I__2230 (
            .O(N__14941),
            .I(N__14938));
    Span4Mux_v I__2229 (
            .O(N__14938),
            .I(N__14935));
    Odrv4 I__2228 (
            .O(N__14935),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    CascadeMux I__2227 (
            .O(N__14932),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ));
    InMux I__2226 (
            .O(N__14929),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__2225 (
            .O(N__14926),
            .I(N__14920));
    InMux I__2224 (
            .O(N__14925),
            .I(N__14920));
    LocalMux I__2223 (
            .O(N__14920),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__2222 (
            .O(N__14917),
            .I(N__14913));
    InMux I__2221 (
            .O(N__14916),
            .I(N__14910));
    LocalMux I__2220 (
            .O(N__14913),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__2219 (
            .O(N__14910),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__2218 (
            .O(N__14905),
            .I(N__14901));
    InMux I__2217 (
            .O(N__14904),
            .I(N__14896));
    InMux I__2216 (
            .O(N__14901),
            .I(N__14896));
    LocalMux I__2215 (
            .O(N__14896),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__2214 (
            .O(N__14893),
            .I(N__14889));
    InMux I__2213 (
            .O(N__14892),
            .I(N__14886));
    LocalMux I__2212 (
            .O(N__14889),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__2211 (
            .O(N__14886),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__2210 (
            .O(N__14881),
            .I(N__14878));
    LocalMux I__2209 (
            .O(N__14878),
            .I(N__14875));
    Odrv12 I__2208 (
            .O(N__14875),
            .I(\reset_module_System.reset6_11 ));
    CascadeMux I__2207 (
            .O(N__14872),
            .I(N__14869));
    InMux I__2206 (
            .O(N__14869),
            .I(N__14866));
    LocalMux I__2205 (
            .O(N__14866),
            .I(N__14863));
    Odrv4 I__2204 (
            .O(N__14863),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_3_0 ));
    CascadeMux I__2203 (
            .O(N__14860),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    CascadeMux I__2202 (
            .O(N__14857),
            .I(N__14854));
    InMux I__2201 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__2200 (
            .O(N__14851),
            .I(\Commands_frame_decoder.state_1_ns_0_a4_0_0_2 ));
    CascadeMux I__2199 (
            .O(N__14848),
            .I(N__14844));
    InMux I__2198 (
            .O(N__14847),
            .I(N__14841));
    InMux I__2197 (
            .O(N__14844),
            .I(N__14838));
    LocalMux I__2196 (
            .O(N__14841),
            .I(N__14835));
    LocalMux I__2195 (
            .O(N__14838),
            .I(N__14832));
    Span4Mux_h I__2194 (
            .O(N__14835),
            .I(N__14828));
    Span4Mux_v I__2193 (
            .O(N__14832),
            .I(N__14825));
    InMux I__2192 (
            .O(N__14831),
            .I(N__14822));
    Odrv4 I__2191 (
            .O(N__14828),
            .I(uart_drone_data_0));
    Odrv4 I__2190 (
            .O(N__14825),
            .I(uart_drone_data_0));
    LocalMux I__2189 (
            .O(N__14822),
            .I(uart_drone_data_0));
    CascadeMux I__2188 (
            .O(N__14815),
            .I(N__14811));
    InMux I__2187 (
            .O(N__14814),
            .I(N__14805));
    InMux I__2186 (
            .O(N__14811),
            .I(N__14800));
    InMux I__2185 (
            .O(N__14810),
            .I(N__14800));
    InMux I__2184 (
            .O(N__14809),
            .I(N__14794));
    InMux I__2183 (
            .O(N__14808),
            .I(N__14794));
    LocalMux I__2182 (
            .O(N__14805),
            .I(N__14790));
    LocalMux I__2181 (
            .O(N__14800),
            .I(N__14787));
    CascadeMux I__2180 (
            .O(N__14799),
            .I(N__14784));
    LocalMux I__2179 (
            .O(N__14794),
            .I(N__14781));
    InMux I__2178 (
            .O(N__14793),
            .I(N__14778));
    Span4Mux_v I__2177 (
            .O(N__14790),
            .I(N__14773));
    Span4Mux_v I__2176 (
            .O(N__14787),
            .I(N__14773));
    InMux I__2175 (
            .O(N__14784),
            .I(N__14770));
    Span4Mux_v I__2174 (
            .O(N__14781),
            .I(N__14765));
    LocalMux I__2173 (
            .O(N__14778),
            .I(N__14765));
    Odrv4 I__2172 (
            .O(N__14773),
            .I(uart_drone_data_1));
    LocalMux I__2171 (
            .O(N__14770),
            .I(uart_drone_data_1));
    Odrv4 I__2170 (
            .O(N__14765),
            .I(uart_drone_data_1));
    InMux I__2169 (
            .O(N__14758),
            .I(N__14755));
    LocalMux I__2168 (
            .O(N__14755),
            .I(N__14751));
    InMux I__2167 (
            .O(N__14754),
            .I(N__14748));
    Odrv12 I__2166 (
            .O(N__14751),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__2165 (
            .O(N__14748),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__2164 (
            .O(N__14743),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__2163 (
            .O(N__14740),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__2162 (
            .O(N__14737),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__2161 (
            .O(N__14734),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__2160 (
            .O(N__14731),
            .I(N__14727));
    InMux I__2159 (
            .O(N__14730),
            .I(N__14724));
    LocalMux I__2158 (
            .O(N__14727),
            .I(N__14721));
    LocalMux I__2157 (
            .O(N__14724),
            .I(\reset_module_System.countZ0Z_16 ));
    Odrv4 I__2156 (
            .O(N__14721),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__2155 (
            .O(N__14716),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__2154 (
            .O(N__14713),
            .I(bfn_4_14_0_));
    InMux I__2153 (
            .O(N__14710),
            .I(N__14706));
    InMux I__2152 (
            .O(N__14709),
            .I(N__14703));
    LocalMux I__2151 (
            .O(N__14706),
            .I(N__14700));
    LocalMux I__2150 (
            .O(N__14703),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__2149 (
            .O(N__14700),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__2148 (
            .O(N__14695),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__2147 (
            .O(N__14692),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__2146 (
            .O(N__14689),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__2145 (
            .O(N__14686),
            .I(N__14682));
    InMux I__2144 (
            .O(N__14685),
            .I(N__14679));
    LocalMux I__2143 (
            .O(N__14682),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__2142 (
            .O(N__14679),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__2141 (
            .O(N__14674),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__2140 (
            .O(N__14671),
            .I(N__14667));
    InMux I__2139 (
            .O(N__14670),
            .I(N__14664));
    LocalMux I__2138 (
            .O(N__14667),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__2137 (
            .O(N__14664),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__2136 (
            .O(N__14659),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__2135 (
            .O(N__14656),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__2134 (
            .O(N__14653),
            .I(N__14649));
    InMux I__2133 (
            .O(N__14652),
            .I(N__14646));
    LocalMux I__2132 (
            .O(N__14649),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__2131 (
            .O(N__14646),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__2130 (
            .O(N__14641),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__2129 (
            .O(N__14638),
            .I(N__14634));
    InMux I__2128 (
            .O(N__14637),
            .I(N__14631));
    LocalMux I__2127 (
            .O(N__14634),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__2126 (
            .O(N__14631),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__2125 (
            .O(N__14626),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__2124 (
            .O(N__14623),
            .I(N__14620));
    InMux I__2123 (
            .O(N__14620),
            .I(N__14616));
    InMux I__2122 (
            .O(N__14619),
            .I(N__14613));
    LocalMux I__2121 (
            .O(N__14616),
            .I(N__14610));
    LocalMux I__2120 (
            .O(N__14613),
            .I(\reset_module_System.countZ0Z_9 ));
    Odrv4 I__2119 (
            .O(N__14610),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__2118 (
            .O(N__14605),
            .I(bfn_4_13_0_));
    InMux I__2117 (
            .O(N__14602),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__2116 (
            .O(N__14599),
            .I(\reset_module_System.count_1_cry_10 ));
    CascadeMux I__2115 (
            .O(N__14596),
            .I(\reset_module_System.reset6_13_cascade_ ));
    InMux I__2114 (
            .O(N__14593),
            .I(N__14590));
    LocalMux I__2113 (
            .O(N__14590),
            .I(\reset_module_System.reset6_3 ));
    CascadeMux I__2112 (
            .O(N__14587),
            .I(\reset_module_System.reset6_17_cascade_ ));
    CascadeMux I__2111 (
            .O(N__14584),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__2110 (
            .O(N__14581),
            .I(N__14577));
    InMux I__2109 (
            .O(N__14580),
            .I(N__14573));
    LocalMux I__2108 (
            .O(N__14577),
            .I(N__14570));
    InMux I__2107 (
            .O(N__14576),
            .I(N__14567));
    LocalMux I__2106 (
            .O(N__14573),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__2105 (
            .O(N__14570),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__2104 (
            .O(N__14567),
            .I(\reset_module_System.countZ0Z_1 ));
    CascadeMux I__2103 (
            .O(N__14560),
            .I(N__14554));
    InMux I__2102 (
            .O(N__14559),
            .I(N__14551));
    InMux I__2101 (
            .O(N__14558),
            .I(N__14546));
    InMux I__2100 (
            .O(N__14557),
            .I(N__14546));
    InMux I__2099 (
            .O(N__14554),
            .I(N__14543));
    LocalMux I__2098 (
            .O(N__14551),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__2097 (
            .O(N__14546),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__2096 (
            .O(N__14543),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__2095 (
            .O(N__14536),
            .I(N__14533));
    LocalMux I__2094 (
            .O(N__14533),
            .I(\reset_module_System.count_1_2 ));
    InMux I__2093 (
            .O(N__14530),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__2092 (
            .O(N__14527),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__2091 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__2090 (
            .O(N__14521),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__2089 (
            .O(N__14518),
            .I(N__14515));
    LocalMux I__2088 (
            .O(N__14515),
            .I(N__14512));
    Span4Mux_h I__2087 (
            .O(N__14512),
            .I(N__14509));
    Odrv4 I__2086 (
            .O(N__14509),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__2085 (
            .O(N__14506),
            .I(N__14503));
    LocalMux I__2084 (
            .O(N__14503),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__2083 (
            .O(N__14500),
            .I(N__14497));
    LocalMux I__2082 (
            .O(N__14497),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ));
    InMux I__2081 (
            .O(N__14494),
            .I(N__14491));
    LocalMux I__2080 (
            .O(N__14491),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__2079 (
            .O(N__14488),
            .I(N__14485));
    LocalMux I__2078 (
            .O(N__14485),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    InMux I__2077 (
            .O(N__14482),
            .I(N__14479));
    LocalMux I__2076 (
            .O(N__14479),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ));
    CascadeMux I__2075 (
            .O(N__14476),
            .I(N__14473));
    InMux I__2074 (
            .O(N__14473),
            .I(N__14470));
    LocalMux I__2073 (
            .O(N__14470),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__2072 (
            .O(N__14467),
            .I(N__14463));
    CascadeMux I__2071 (
            .O(N__14466),
            .I(N__14459));
    LocalMux I__2070 (
            .O(N__14463),
            .I(N__14456));
    InMux I__2069 (
            .O(N__14462),
            .I(N__14453));
    InMux I__2068 (
            .O(N__14459),
            .I(N__14450));
    Span12Mux_h I__2067 (
            .O(N__14456),
            .I(N__14445));
    LocalMux I__2066 (
            .O(N__14453),
            .I(N__14445));
    LocalMux I__2065 (
            .O(N__14450),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv12 I__2064 (
            .O(N__14445),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    InMux I__2063 (
            .O(N__14440),
            .I(N__14437));
    LocalMux I__2062 (
            .O(N__14437),
            .I(N__14434));
    Odrv12 I__2061 (
            .O(N__14434),
            .I(\ppm_encoder_1.N_295 ));
    InMux I__2060 (
            .O(N__14431),
            .I(N__14428));
    LocalMux I__2059 (
            .O(N__14428),
            .I(N__14424));
    InMux I__2058 (
            .O(N__14427),
            .I(N__14421));
    Odrv12 I__2057 (
            .O(N__14424),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    LocalMux I__2056 (
            .O(N__14421),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    CascadeMux I__2055 (
            .O(N__14416),
            .I(\reset_module_System.count_1_1_cascade_ ));
    InMux I__2054 (
            .O(N__14413),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__2053 (
            .O(N__14410),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__2052 (
            .O(N__14407),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__2051 (
            .O(N__14404),
            .I(bfn_3_27_0_));
    CascadeMux I__2050 (
            .O(N__14401),
            .I(N__14398));
    InMux I__2049 (
            .O(N__14398),
            .I(N__14395));
    LocalMux I__2048 (
            .O(N__14395),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__2047 (
            .O(N__14392),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__2046 (
            .O(N__14389),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__2045 (
            .O(N__14386),
            .I(N__14383));
    LocalMux I__2044 (
            .O(N__14383),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__2043 (
            .O(N__14380),
            .I(N__14375));
    InMux I__2042 (
            .O(N__14379),
            .I(N__14370));
    InMux I__2041 (
            .O(N__14378),
            .I(N__14370));
    LocalMux I__2040 (
            .O(N__14375),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    LocalMux I__2039 (
            .O(N__14370),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    CascadeMux I__2038 (
            .O(N__14365),
            .I(N__14362));
    InMux I__2037 (
            .O(N__14362),
            .I(N__14359));
    LocalMux I__2036 (
            .O(N__14359),
            .I(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ));
    InMux I__2035 (
            .O(N__14356),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    CascadeMux I__2034 (
            .O(N__14353),
            .I(N__14350));
    InMux I__2033 (
            .O(N__14350),
            .I(N__14347));
    LocalMux I__2032 (
            .O(N__14347),
            .I(N__14344));
    Span4Mux_v I__2031 (
            .O(N__14344),
            .I(N__14341));
    Odrv4 I__2030 (
            .O(N__14341),
            .I(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ));
    InMux I__2029 (
            .O(N__14338),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__2028 (
            .O(N__14335),
            .I(N__14331));
    InMux I__2027 (
            .O(N__14334),
            .I(N__14328));
    LocalMux I__2026 (
            .O(N__14331),
            .I(N__14325));
    LocalMux I__2025 (
            .O(N__14328),
            .I(N__14322));
    Span4Mux_v I__2024 (
            .O(N__14325),
            .I(N__14319));
    Span4Mux_h I__2023 (
            .O(N__14322),
            .I(N__14316));
    Odrv4 I__2022 (
            .O(N__14319),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    Odrv4 I__2021 (
            .O(N__14316),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    CascadeMux I__2020 (
            .O(N__14311),
            .I(N__14308));
    InMux I__2019 (
            .O(N__14308),
            .I(N__14305));
    LocalMux I__2018 (
            .O(N__14305),
            .I(N__14302));
    Odrv4 I__2017 (
            .O(N__14302),
            .I(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ));
    InMux I__2016 (
            .O(N__14299),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__2015 (
            .O(N__14296),
            .I(N__14293));
    LocalMux I__2014 (
            .O(N__14293),
            .I(N__14289));
    InMux I__2013 (
            .O(N__14292),
            .I(N__14286));
    Span4Mux_v I__2012 (
            .O(N__14289),
            .I(N__14281));
    LocalMux I__2011 (
            .O(N__14286),
            .I(N__14281));
    Odrv4 I__2010 (
            .O(N__14281),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    CascadeMux I__2009 (
            .O(N__14278),
            .I(N__14275));
    InMux I__2008 (
            .O(N__14275),
            .I(N__14272));
    LocalMux I__2007 (
            .O(N__14272),
            .I(N__14269));
    Odrv12 I__2006 (
            .O(N__14269),
            .I(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ));
    InMux I__2005 (
            .O(N__14266),
            .I(N__14263));
    LocalMux I__2004 (
            .O(N__14263),
            .I(N__14260));
    Span4Mux_s2_v I__2003 (
            .O(N__14260),
            .I(N__14257));
    Odrv4 I__2002 (
            .O(N__14257),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__2001 (
            .O(N__14254),
            .I(bfn_3_26_0_));
    InMux I__2000 (
            .O(N__14251),
            .I(N__14248));
    LocalMux I__1999 (
            .O(N__14248),
            .I(N__14244));
    InMux I__1998 (
            .O(N__14247),
            .I(N__14241));
    Span4Mux_v I__1997 (
            .O(N__14244),
            .I(N__14236));
    LocalMux I__1996 (
            .O(N__14241),
            .I(N__14236));
    Odrv4 I__1995 (
            .O(N__14236),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    CascadeMux I__1994 (
            .O(N__14233),
            .I(N__14230));
    InMux I__1993 (
            .O(N__14230),
            .I(N__14227));
    LocalMux I__1992 (
            .O(N__14227),
            .I(N__14224));
    Odrv4 I__1991 (
            .O(N__14224),
            .I(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ));
    InMux I__1990 (
            .O(N__14221),
            .I(N__14218));
    LocalMux I__1989 (
            .O(N__14218),
            .I(N__14215));
    Span4Mux_s3_v I__1988 (
            .O(N__14215),
            .I(N__14212));
    Odrv4 I__1987 (
            .O(N__14212),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__1986 (
            .O(N__14209),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__1985 (
            .O(N__14206),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__1984 (
            .O(N__14203),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__1983 (
            .O(N__14200),
            .I(N__14196));
    InMux I__1982 (
            .O(N__14199),
            .I(N__14193));
    LocalMux I__1981 (
            .O(N__14196),
            .I(N__14190));
    LocalMux I__1980 (
            .O(N__14193),
            .I(N__14187));
    Span4Mux_h I__1979 (
            .O(N__14190),
            .I(N__14182));
    Span4Mux_h I__1978 (
            .O(N__14187),
            .I(N__14182));
    Odrv4 I__1977 (
            .O(N__14182),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    CascadeMux I__1976 (
            .O(N__14179),
            .I(N__14176));
    InMux I__1975 (
            .O(N__14176),
            .I(N__14173));
    LocalMux I__1974 (
            .O(N__14173),
            .I(N__14170));
    Odrv12 I__1973 (
            .O(N__14170),
            .I(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ));
    InMux I__1972 (
            .O(N__14167),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    CascadeMux I__1971 (
            .O(N__14164),
            .I(N__14161));
    InMux I__1970 (
            .O(N__14161),
            .I(N__14158));
    LocalMux I__1969 (
            .O(N__14158),
            .I(N__14155));
    Span4Mux_v I__1968 (
            .O(N__14155),
            .I(N__14152));
    Odrv4 I__1967 (
            .O(N__14152),
            .I(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ));
    CascadeMux I__1966 (
            .O(N__14149),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ));
    InMux I__1965 (
            .O(N__14146),
            .I(N__14143));
    LocalMux I__1964 (
            .O(N__14143),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5 ));
    InMux I__1963 (
            .O(N__14140),
            .I(N__14137));
    LocalMux I__1962 (
            .O(N__14137),
            .I(N__14134));
    Odrv4 I__1961 (
            .O(N__14134),
            .I(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ));
    CascadeMux I__1960 (
            .O(N__14131),
            .I(N__14128));
    InMux I__1959 (
            .O(N__14128),
            .I(N__14124));
    InMux I__1958 (
            .O(N__14127),
            .I(N__14121));
    LocalMux I__1957 (
            .O(N__14124),
            .I(N__14118));
    LocalMux I__1956 (
            .O(N__14121),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    Odrv4 I__1955 (
            .O(N__14118),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    CascadeMux I__1954 (
            .O(N__14113),
            .I(N__14110));
    InMux I__1953 (
            .O(N__14110),
            .I(N__14107));
    LocalMux I__1952 (
            .O(N__14107),
            .I(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ));
    InMux I__1951 (
            .O(N__14104),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__1950 (
            .O(N__14101),
            .I(N__14098));
    LocalMux I__1949 (
            .O(N__14098),
            .I(N__14094));
    InMux I__1948 (
            .O(N__14097),
            .I(N__14091));
    Odrv4 I__1947 (
            .O(N__14094),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    LocalMux I__1946 (
            .O(N__14091),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    CascadeMux I__1945 (
            .O(N__14086),
            .I(N__14083));
    InMux I__1944 (
            .O(N__14083),
            .I(N__14080));
    LocalMux I__1943 (
            .O(N__14080),
            .I(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ));
    InMux I__1942 (
            .O(N__14077),
            .I(N__14074));
    LocalMux I__1941 (
            .O(N__14074),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__1940 (
            .O(N__14071),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__1939 (
            .O(N__14068),
            .I(N__14065));
    LocalMux I__1938 (
            .O(N__14065),
            .I(N__14061));
    InMux I__1937 (
            .O(N__14064),
            .I(N__14058));
    Odrv4 I__1936 (
            .O(N__14061),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    LocalMux I__1935 (
            .O(N__14058),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    CascadeMux I__1934 (
            .O(N__14053),
            .I(N__14050));
    InMux I__1933 (
            .O(N__14050),
            .I(N__14047));
    LocalMux I__1932 (
            .O(N__14047),
            .I(N__14044));
    Odrv4 I__1931 (
            .O(N__14044),
            .I(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ));
    InMux I__1930 (
            .O(N__14041),
            .I(N__14038));
    LocalMux I__1929 (
            .O(N__14038),
            .I(N__14035));
    Odrv4 I__1928 (
            .O(N__14035),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__1927 (
            .O(N__14032),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    CascadeMux I__1926 (
            .O(N__14029),
            .I(N__14026));
    InMux I__1925 (
            .O(N__14026),
            .I(N__14023));
    LocalMux I__1924 (
            .O(N__14023),
            .I(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ));
    InMux I__1923 (
            .O(N__14020),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__1922 (
            .O(N__14017),
            .I(N__14014));
    LocalMux I__1921 (
            .O(N__14014),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8 ));
    CascadeMux I__1920 (
            .O(N__14011),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ));
    InMux I__1919 (
            .O(N__14008),
            .I(N__14005));
    LocalMux I__1918 (
            .O(N__14005),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9 ));
    InMux I__1917 (
            .O(N__14002),
            .I(N__13999));
    LocalMux I__1916 (
            .O(N__13999),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4 ));
    InMux I__1915 (
            .O(N__13996),
            .I(N__13991));
    InMux I__1914 (
            .O(N__13995),
            .I(N__13988));
    CascadeMux I__1913 (
            .O(N__13994),
            .I(N__13985));
    LocalMux I__1912 (
            .O(N__13991),
            .I(N__13982));
    LocalMux I__1911 (
            .O(N__13988),
            .I(N__13979));
    InMux I__1910 (
            .O(N__13985),
            .I(N__13976));
    Span4Mux_v I__1909 (
            .O(N__13982),
            .I(N__13973));
    Span4Mux_v I__1908 (
            .O(N__13979),
            .I(N__13970));
    LocalMux I__1907 (
            .O(N__13976),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__1906 (
            .O(N__13973),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__1905 (
            .O(N__13970),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__1904 (
            .O(N__13963),
            .I(N__13957));
    InMux I__1903 (
            .O(N__13962),
            .I(N__13957));
    LocalMux I__1902 (
            .O(N__13957),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__1901 (
            .O(N__13954),
            .I(N__13951));
    LocalMux I__1900 (
            .O(N__13951),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__1899 (
            .O(N__13948),
            .I(N__13945));
    LocalMux I__1898 (
            .O(N__13945),
            .I(N__13941));
    InMux I__1897 (
            .O(N__13944),
            .I(N__13938));
    Span4Mux_v I__1896 (
            .O(N__13941),
            .I(N__13935));
    LocalMux I__1895 (
            .O(N__13938),
            .I(N__13932));
    Span4Mux_v I__1894 (
            .O(N__13935),
            .I(N__13929));
    Span4Mux_v I__1893 (
            .O(N__13932),
            .I(N__13926));
    Span4Mux_v I__1892 (
            .O(N__13929),
            .I(N__13923));
    Span4Mux_v I__1891 (
            .O(N__13926),
            .I(N__13920));
    Odrv4 I__1890 (
            .O(N__13923),
            .I(throttle_command_12));
    Odrv4 I__1889 (
            .O(N__13920),
            .I(throttle_command_12));
    InMux I__1888 (
            .O(N__13915),
            .I(N__13912));
    LocalMux I__1887 (
            .O(N__13912),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    CascadeMux I__1886 (
            .O(N__13909),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    InMux I__1885 (
            .O(N__13906),
            .I(N__13903));
    LocalMux I__1884 (
            .O(N__13903),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    InMux I__1883 (
            .O(N__13900),
            .I(N__13895));
    InMux I__1882 (
            .O(N__13899),
            .I(N__13890));
    InMux I__1881 (
            .O(N__13898),
            .I(N__13890));
    LocalMux I__1880 (
            .O(N__13895),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    LocalMux I__1879 (
            .O(N__13890),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    CascadeMux I__1878 (
            .O(N__13885),
            .I(\ppm_encoder_1.N_303_cascade_ ));
    InMux I__1877 (
            .O(N__13882),
            .I(N__13873));
    InMux I__1876 (
            .O(N__13881),
            .I(N__13873));
    InMux I__1875 (
            .O(N__13880),
            .I(N__13873));
    LocalMux I__1874 (
            .O(N__13873),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    CascadeMux I__1873 (
            .O(N__13870),
            .I(N__13867));
    InMux I__1872 (
            .O(N__13867),
            .I(N__13862));
    InMux I__1871 (
            .O(N__13866),
            .I(N__13859));
    InMux I__1870 (
            .O(N__13865),
            .I(N__13856));
    LocalMux I__1869 (
            .O(N__13862),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    LocalMux I__1868 (
            .O(N__13859),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    LocalMux I__1867 (
            .O(N__13856),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    CascadeMux I__1866 (
            .O(N__13849),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ));
    IoInMux I__1865 (
            .O(N__13846),
            .I(N__13843));
    LocalMux I__1864 (
            .O(N__13843),
            .I(N__13840));
    IoSpan4Mux I__1863 (
            .O(N__13840),
            .I(N__13837));
    Span4Mux_s3_v I__1862 (
            .O(N__13837),
            .I(N__13833));
    InMux I__1861 (
            .O(N__13836),
            .I(N__13830));
    Span4Mux_v I__1860 (
            .O(N__13833),
            .I(N__13823));
    LocalMux I__1859 (
            .O(N__13830),
            .I(N__13823));
    InMux I__1858 (
            .O(N__13829),
            .I(N__13818));
    InMux I__1857 (
            .O(N__13828),
            .I(N__13818));
    Sp12to4 I__1856 (
            .O(N__13823),
            .I(N__13815));
    LocalMux I__1855 (
            .O(N__13818),
            .I(drone_frame_decoder_data_rdy_debug_c));
    Odrv12 I__1854 (
            .O(N__13815),
            .I(drone_frame_decoder_data_rdy_debug_c));
    CascadeMux I__1853 (
            .O(N__13810),
            .I(\uart_pc.N_152_cascade_ ));
    CascadeMux I__1852 (
            .O(N__13807),
            .I(\uart_pc.CO0_cascade_ ));
    InMux I__1851 (
            .O(N__13804),
            .I(N__13798));
    InMux I__1850 (
            .O(N__13803),
            .I(N__13798));
    LocalMux I__1849 (
            .O(N__13798),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__1848 (
            .O(N__13795),
            .I(N__13792));
    LocalMux I__1847 (
            .O(N__13792),
            .I(N__13788));
    InMux I__1846 (
            .O(N__13791),
            .I(N__13785));
    Span4Mux_h I__1845 (
            .O(N__13788),
            .I(N__13780));
    LocalMux I__1844 (
            .O(N__13785),
            .I(N__13780));
    Span4Mux_v I__1843 (
            .O(N__13780),
            .I(N__13777));
    Span4Mux_v I__1842 (
            .O(N__13777),
            .I(N__13774));
    Odrv4 I__1841 (
            .O(N__13774),
            .I(throttle_command_9));
    InMux I__1840 (
            .O(N__13771),
            .I(N__13768));
    LocalMux I__1839 (
            .O(N__13768),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__1838 (
            .O(N__13765),
            .I(N__13762));
    LocalMux I__1837 (
            .O(N__13762),
            .I(N__13759));
    Span4Mux_v I__1836 (
            .O(N__13759),
            .I(N__13756));
    Sp12to4 I__1835 (
            .O(N__13756),
            .I(N__13752));
    InMux I__1834 (
            .O(N__13755),
            .I(N__13749));
    Span12Mux_s2_h I__1833 (
            .O(N__13752),
            .I(N__13744));
    LocalMux I__1832 (
            .O(N__13749),
            .I(N__13744));
    Span12Mux_v I__1831 (
            .O(N__13744),
            .I(N__13741));
    Odrv12 I__1830 (
            .O(N__13741),
            .I(throttle_command_11));
    CascadeMux I__1829 (
            .O(N__13738),
            .I(N__13735));
    InMux I__1828 (
            .O(N__13735),
            .I(N__13732));
    LocalMux I__1827 (
            .O(N__13732),
            .I(N__13729));
    Odrv4 I__1826 (
            .O(N__13729),
            .I(alt_command_7));
    CEMux I__1825 (
            .O(N__13726),
            .I(N__13723));
    LocalMux I__1824 (
            .O(N__13723),
            .I(N__13718));
    CEMux I__1823 (
            .O(N__13722),
            .I(N__13715));
    CEMux I__1822 (
            .O(N__13721),
            .I(N__13712));
    Span4Mux_v I__1821 (
            .O(N__13718),
            .I(N__13707));
    LocalMux I__1820 (
            .O(N__13715),
            .I(N__13707));
    LocalMux I__1819 (
            .O(N__13712),
            .I(N__13704));
    Span4Mux_v I__1818 (
            .O(N__13707),
            .I(N__13699));
    Span4Mux_v I__1817 (
            .O(N__13704),
            .I(N__13699));
    Span4Mux_s2_h I__1816 (
            .O(N__13699),
            .I(N__13696));
    Odrv4 I__1815 (
            .O(N__13696),
            .I(\dron_frame_decoder_1.N_238_0 ));
    InMux I__1814 (
            .O(N__13693),
            .I(N__13690));
    LocalMux I__1813 (
            .O(N__13690),
            .I(N__13686));
    InMux I__1812 (
            .O(N__13689),
            .I(N__13677));
    Span4Mux_v I__1811 (
            .O(N__13686),
            .I(N__13674));
    InMux I__1810 (
            .O(N__13685),
            .I(N__13663));
    InMux I__1809 (
            .O(N__13684),
            .I(N__13663));
    InMux I__1808 (
            .O(N__13683),
            .I(N__13663));
    InMux I__1807 (
            .O(N__13682),
            .I(N__13663));
    InMux I__1806 (
            .O(N__13681),
            .I(N__13663));
    InMux I__1805 (
            .O(N__13680),
            .I(N__13660));
    LocalMux I__1804 (
            .O(N__13677),
            .I(\dron_frame_decoder_1.N_237 ));
    Odrv4 I__1803 (
            .O(N__13674),
            .I(\dron_frame_decoder_1.N_237 ));
    LocalMux I__1802 (
            .O(N__13663),
            .I(\dron_frame_decoder_1.N_237 ));
    LocalMux I__1801 (
            .O(N__13660),
            .I(\dron_frame_decoder_1.N_237 ));
    InMux I__1800 (
            .O(N__13651),
            .I(N__13647));
    CascadeMux I__1799 (
            .O(N__13650),
            .I(N__13644));
    LocalMux I__1798 (
            .O(N__13647),
            .I(N__13640));
    InMux I__1797 (
            .O(N__13644),
            .I(N__13635));
    InMux I__1796 (
            .O(N__13643),
            .I(N__13635));
    Odrv12 I__1795 (
            .O(N__13640),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__1794 (
            .O(N__13635),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    InMux I__1793 (
            .O(N__13630),
            .I(N__13627));
    LocalMux I__1792 (
            .O(N__13627),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_0_0 ));
    InMux I__1791 (
            .O(N__13624),
            .I(N__13621));
    LocalMux I__1790 (
            .O(N__13621),
            .I(N__13616));
    InMux I__1789 (
            .O(N__13620),
            .I(N__13611));
    InMux I__1788 (
            .O(N__13619),
            .I(N__13611));
    Span4Mux_v I__1787 (
            .O(N__13616),
            .I(N__13608));
    LocalMux I__1786 (
            .O(N__13611),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    Odrv4 I__1785 (
            .O(N__13608),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    CascadeMux I__1784 (
            .O(N__13603),
            .I(N__13599));
    InMux I__1783 (
            .O(N__13602),
            .I(N__13590));
    InMux I__1782 (
            .O(N__13599),
            .I(N__13590));
    InMux I__1781 (
            .O(N__13598),
            .I(N__13590));
    InMux I__1780 (
            .O(N__13597),
            .I(N__13587));
    LocalMux I__1779 (
            .O(N__13590),
            .I(N__13584));
    LocalMux I__1778 (
            .O(N__13587),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    Odrv12 I__1777 (
            .O(N__13584),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    CascadeMux I__1776 (
            .O(N__13579),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_ ));
    CascadeMux I__1775 (
            .O(N__13576),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ));
    CEMux I__1774 (
            .O(N__13573),
            .I(N__13569));
    CEMux I__1773 (
            .O(N__13572),
            .I(N__13565));
    LocalMux I__1772 (
            .O(N__13569),
            .I(N__13562));
    CEMux I__1771 (
            .O(N__13568),
            .I(N__13559));
    LocalMux I__1770 (
            .O(N__13565),
            .I(N__13556));
    Span4Mux_v I__1769 (
            .O(N__13562),
            .I(N__13553));
    LocalMux I__1768 (
            .O(N__13559),
            .I(N__13550));
    Span4Mux_v I__1767 (
            .O(N__13556),
            .I(N__13547));
    Span4Mux_s3_h I__1766 (
            .O(N__13553),
            .I(N__13544));
    Sp12to4 I__1765 (
            .O(N__13550),
            .I(N__13541));
    Odrv4 I__1764 (
            .O(N__13547),
            .I(\dron_frame_decoder_1.N_230_0 ));
    Odrv4 I__1763 (
            .O(N__13544),
            .I(\dron_frame_decoder_1.N_230_0 ));
    Odrv12 I__1762 (
            .O(N__13541),
            .I(\dron_frame_decoder_1.N_230_0 ));
    InMux I__1761 (
            .O(N__13534),
            .I(N__13527));
    InMux I__1760 (
            .O(N__13533),
            .I(N__13527));
    InMux I__1759 (
            .O(N__13532),
            .I(N__13522));
    LocalMux I__1758 (
            .O(N__13527),
            .I(N__13518));
    InMux I__1757 (
            .O(N__13526),
            .I(N__13515));
    InMux I__1756 (
            .O(N__13525),
            .I(N__13512));
    LocalMux I__1755 (
            .O(N__13522),
            .I(N__13509));
    InMux I__1754 (
            .O(N__13521),
            .I(N__13506));
    Span4Mux_v I__1753 (
            .O(N__13518),
            .I(N__13501));
    LocalMux I__1752 (
            .O(N__13515),
            .I(N__13501));
    LocalMux I__1751 (
            .O(N__13512),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv12 I__1750 (
            .O(N__13509),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__1749 (
            .O(N__13506),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__1748 (
            .O(N__13501),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    IoInMux I__1747 (
            .O(N__13492),
            .I(N__13489));
    LocalMux I__1746 (
            .O(N__13489),
            .I(N__13486));
    IoSpan4Mux I__1745 (
            .O(N__13486),
            .I(N__13479));
    CascadeMux I__1744 (
            .O(N__13485),
            .I(N__13475));
    CascadeMux I__1743 (
            .O(N__13484),
            .I(N__13472));
    CascadeMux I__1742 (
            .O(N__13483),
            .I(N__13469));
    CascadeMux I__1741 (
            .O(N__13482),
            .I(N__13465));
    Sp12to4 I__1740 (
            .O(N__13479),
            .I(N__13461));
    InMux I__1739 (
            .O(N__13478),
            .I(N__13451));
    InMux I__1738 (
            .O(N__13475),
            .I(N__13451));
    InMux I__1737 (
            .O(N__13472),
            .I(N__13451));
    InMux I__1736 (
            .O(N__13469),
            .I(N__13451));
    InMux I__1735 (
            .O(N__13468),
            .I(N__13448));
    InMux I__1734 (
            .O(N__13465),
            .I(N__13445));
    InMux I__1733 (
            .O(N__13464),
            .I(N__13442));
    Span12Mux_s9_v I__1732 (
            .O(N__13461),
            .I(N__13438));
    InMux I__1731 (
            .O(N__13460),
            .I(N__13435));
    LocalMux I__1730 (
            .O(N__13451),
            .I(N__13430));
    LocalMux I__1729 (
            .O(N__13448),
            .I(N__13430));
    LocalMux I__1728 (
            .O(N__13445),
            .I(N__13425));
    LocalMux I__1727 (
            .O(N__13442),
            .I(N__13425));
    InMux I__1726 (
            .O(N__13441),
            .I(N__13420));
    Span12Mux_h I__1725 (
            .O(N__13438),
            .I(N__13415));
    LocalMux I__1724 (
            .O(N__13435),
            .I(N__13415));
    Span4Mux_v I__1723 (
            .O(N__13430),
            .I(N__13410));
    Span4Mux_v I__1722 (
            .O(N__13425),
            .I(N__13410));
    InMux I__1721 (
            .O(N__13424),
            .I(N__13405));
    InMux I__1720 (
            .O(N__13423),
            .I(N__13405));
    LocalMux I__1719 (
            .O(N__13420),
            .I(uart_drone_data_rdy_debug_c));
    Odrv12 I__1718 (
            .O(N__13415),
            .I(uart_drone_data_rdy_debug_c));
    Odrv4 I__1717 (
            .O(N__13410),
            .I(uart_drone_data_rdy_debug_c));
    LocalMux I__1716 (
            .O(N__13405),
            .I(uart_drone_data_rdy_debug_c));
    CascadeMux I__1715 (
            .O(N__13396),
            .I(\dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_ ));
    InMux I__1714 (
            .O(N__13393),
            .I(N__13390));
    LocalMux I__1713 (
            .O(N__13390),
            .I(\dron_frame_decoder_1.N_239 ));
    InMux I__1712 (
            .O(N__13387),
            .I(N__13382));
    InMux I__1711 (
            .O(N__13386),
            .I(N__13375));
    InMux I__1710 (
            .O(N__13385),
            .I(N__13375));
    LocalMux I__1709 (
            .O(N__13382),
            .I(N__13372));
    InMux I__1708 (
            .O(N__13381),
            .I(N__13367));
    InMux I__1707 (
            .O(N__13380),
            .I(N__13367));
    LocalMux I__1706 (
            .O(N__13375),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    Odrv4 I__1705 (
            .O(N__13372),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__1704 (
            .O(N__13367),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__1703 (
            .O(N__13360),
            .I(N__13357));
    LocalMux I__1702 (
            .O(N__13357),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ));
    CascadeMux I__1701 (
            .O(N__13354),
            .I(\dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ));
    InMux I__1700 (
            .O(N__13351),
            .I(N__13348));
    LocalMux I__1699 (
            .O(N__13348),
            .I(N__13344));
    InMux I__1698 (
            .O(N__13347),
            .I(N__13341));
    Span4Mux_s3_h I__1697 (
            .O(N__13344),
            .I(N__13335));
    LocalMux I__1696 (
            .O(N__13341),
            .I(N__13335));
    InMux I__1695 (
            .O(N__13340),
            .I(N__13332));
    Odrv4 I__1694 (
            .O(N__13335),
            .I(\dron_frame_decoder_1.N_243 ));
    LocalMux I__1693 (
            .O(N__13332),
            .I(\dron_frame_decoder_1.N_243 ));
    CascadeMux I__1692 (
            .O(N__13327),
            .I(N__13324));
    InMux I__1691 (
            .O(N__13324),
            .I(N__13321));
    LocalMux I__1690 (
            .O(N__13321),
            .I(N__13318));
    Odrv4 I__1689 (
            .O(N__13318),
            .I(alt_command_4));
    CascadeMux I__1688 (
            .O(N__13315),
            .I(N__13312));
    InMux I__1687 (
            .O(N__13312),
            .I(N__13309));
    LocalMux I__1686 (
            .O(N__13309),
            .I(N__13306));
    Odrv4 I__1685 (
            .O(N__13306),
            .I(alt_command_5));
    CascadeMux I__1684 (
            .O(N__13303),
            .I(N__13300));
    InMux I__1683 (
            .O(N__13300),
            .I(N__13297));
    LocalMux I__1682 (
            .O(N__13297),
            .I(N__13294));
    Odrv4 I__1681 (
            .O(N__13294),
            .I(alt_command_6));
    InMux I__1680 (
            .O(N__13291),
            .I(N__13288));
    LocalMux I__1679 (
            .O(N__13288),
            .I(\dron_frame_decoder_1.state_ns_0_a3_0_3_3 ));
    CascadeMux I__1678 (
            .O(N__13285),
            .I(N__13281));
    CascadeMux I__1677 (
            .O(N__13284),
            .I(N__13278));
    InMux I__1676 (
            .O(N__13281),
            .I(N__13273));
    InMux I__1675 (
            .O(N__13278),
            .I(N__13273));
    LocalMux I__1674 (
            .O(N__13273),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    InMux I__1673 (
            .O(N__13270),
            .I(N__13264));
    InMux I__1672 (
            .O(N__13269),
            .I(N__13264));
    LocalMux I__1671 (
            .O(N__13264),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__1670 (
            .O(N__13261),
            .I(\dron_frame_decoder_1.N_217_cascade_ ));
    CascadeMux I__1669 (
            .O(N__13258),
            .I(N__13254));
    InMux I__1668 (
            .O(N__13257),
            .I(N__13250));
    InMux I__1667 (
            .O(N__13254),
            .I(N__13247));
    InMux I__1666 (
            .O(N__13253),
            .I(N__13244));
    LocalMux I__1665 (
            .O(N__13250),
            .I(N__13241));
    LocalMux I__1664 (
            .O(N__13247),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__1663 (
            .O(N__13244),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv4 I__1662 (
            .O(N__13241),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__1661 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__1660 (
            .O(N__13231),
            .I(\dron_frame_decoder_1.N_219 ));
    InMux I__1659 (
            .O(N__13228),
            .I(N__13225));
    LocalMux I__1658 (
            .O(N__13225),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__1657 (
            .O(N__13222),
            .I(N__13213));
    InMux I__1656 (
            .O(N__13221),
            .I(N__13213));
    InMux I__1655 (
            .O(N__13220),
            .I(N__13213));
    LocalMux I__1654 (
            .O(N__13213),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__1653 (
            .O(N__13210),
            .I(N__13207));
    LocalMux I__1652 (
            .O(N__13207),
            .I(N__13204));
    Span4Mux_s2_v I__1651 (
            .O(N__13204),
            .I(N__13201));
    Span4Mux_v I__1650 (
            .O(N__13201),
            .I(N__13198));
    Odrv4 I__1649 (
            .O(N__13198),
            .I(\ppm_encoder_1.N_299 ));
    InMux I__1648 (
            .O(N__13195),
            .I(N__13191));
    CascadeMux I__1647 (
            .O(N__13194),
            .I(N__13188));
    LocalMux I__1646 (
            .O(N__13191),
            .I(N__13185));
    InMux I__1645 (
            .O(N__13188),
            .I(N__13182));
    Span4Mux_s3_h I__1644 (
            .O(N__13185),
            .I(N__13179));
    LocalMux I__1643 (
            .O(N__13182),
            .I(alt_kp_7));
    Odrv4 I__1642 (
            .O(N__13179),
            .I(alt_kp_7));
    InMux I__1641 (
            .O(N__13174),
            .I(N__13170));
    CascadeMux I__1640 (
            .O(N__13173),
            .I(N__13167));
    LocalMux I__1639 (
            .O(N__13170),
            .I(N__13164));
    InMux I__1638 (
            .O(N__13167),
            .I(N__13161));
    Span4Mux_s3_h I__1637 (
            .O(N__13164),
            .I(N__13158));
    LocalMux I__1636 (
            .O(N__13161),
            .I(alt_kp_5));
    Odrv4 I__1635 (
            .O(N__13158),
            .I(alt_kp_5));
    CascadeMux I__1634 (
            .O(N__13153),
            .I(\dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_ ));
    CascadeMux I__1633 (
            .O(N__13150),
            .I(\dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_ ));
    InMux I__1632 (
            .O(N__13147),
            .I(N__13144));
    LocalMux I__1631 (
            .O(N__13144),
            .I(\dron_frame_decoder_1.state_ns_0_a3_0_3_1 ));
    InMux I__1630 (
            .O(N__13141),
            .I(N__13138));
    LocalMux I__1629 (
            .O(N__13138),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ));
    CascadeMux I__1628 (
            .O(N__13135),
            .I(N__13130));
    CascadeMux I__1627 (
            .O(N__13134),
            .I(N__13125));
    InMux I__1626 (
            .O(N__13133),
            .I(N__13118));
    InMux I__1625 (
            .O(N__13130),
            .I(N__13118));
    CascadeMux I__1624 (
            .O(N__13129),
            .I(N__13115));
    InMux I__1623 (
            .O(N__13128),
            .I(N__13104));
    InMux I__1622 (
            .O(N__13125),
            .I(N__13104));
    InMux I__1621 (
            .O(N__13124),
            .I(N__13104));
    InMux I__1620 (
            .O(N__13123),
            .I(N__13104));
    LocalMux I__1619 (
            .O(N__13118),
            .I(N__13101));
    InMux I__1618 (
            .O(N__13115),
            .I(N__13096));
    InMux I__1617 (
            .O(N__13114),
            .I(N__13096));
    InMux I__1616 (
            .O(N__13113),
            .I(N__13093));
    LocalMux I__1615 (
            .O(N__13104),
            .I(N__13090));
    Odrv4 I__1614 (
            .O(N__13101),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__1613 (
            .O(N__13096),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__1612 (
            .O(N__13093),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    Odrv4 I__1611 (
            .O(N__13090),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    InMux I__1610 (
            .O(N__13081),
            .I(N__13078));
    LocalMux I__1609 (
            .O(N__13078),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ));
    InMux I__1608 (
            .O(N__13075),
            .I(N__13072));
    LocalMux I__1607 (
            .O(N__13072),
            .I(N__13069));
    Odrv4 I__1606 (
            .O(N__13069),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    CascadeMux I__1605 (
            .O(N__13066),
            .I(N__13063));
    InMux I__1604 (
            .O(N__13063),
            .I(N__13060));
    LocalMux I__1603 (
            .O(N__13060),
            .I(N__13057));
    Odrv4 I__1602 (
            .O(N__13057),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__1601 (
            .O(N__13054),
            .I(N__13051));
    LocalMux I__1600 (
            .O(N__13051),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__1599 (
            .O(N__13048),
            .I(N__13045));
    LocalMux I__1598 (
            .O(N__13045),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__1597 (
            .O(N__13042),
            .I(N__13033));
    InMux I__1596 (
            .O(N__13041),
            .I(N__13033));
    InMux I__1595 (
            .O(N__13040),
            .I(N__13033));
    LocalMux I__1594 (
            .O(N__13033),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__1593 (
            .O(N__13030),
            .I(N__13027));
    LocalMux I__1592 (
            .O(N__13027),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    CascadeMux I__1591 (
            .O(N__13024),
            .I(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ));
    CascadeMux I__1590 (
            .O(N__13021),
            .I(\ppm_encoder_1.un1_init_pulses_0_cascade_ ));
    InMux I__1589 (
            .O(N__13018),
            .I(N__13015));
    LocalMux I__1588 (
            .O(N__13015),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    InMux I__1587 (
            .O(N__13012),
            .I(N__13009));
    LocalMux I__1586 (
            .O(N__13009),
            .I(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ));
    InMux I__1585 (
            .O(N__13006),
            .I(N__13003));
    LocalMux I__1584 (
            .O(N__13003),
            .I(N__13000));
    Span4Mux_v I__1583 (
            .O(N__13000),
            .I(N__12996));
    InMux I__1582 (
            .O(N__12999),
            .I(N__12993));
    Span4Mux_v I__1581 (
            .O(N__12996),
            .I(N__12988));
    LocalMux I__1580 (
            .O(N__12993),
            .I(N__12988));
    Span4Mux_v I__1579 (
            .O(N__12988),
            .I(N__12985));
    Span4Mux_v I__1578 (
            .O(N__12985),
            .I(N__12982));
    Odrv4 I__1577 (
            .O(N__12982),
            .I(throttle_command_0));
    CascadeMux I__1576 (
            .O(N__12979),
            .I(N__12976));
    InMux I__1575 (
            .O(N__12976),
            .I(N__12964));
    InMux I__1574 (
            .O(N__12975),
            .I(N__12964));
    InMux I__1573 (
            .O(N__12974),
            .I(N__12964));
    InMux I__1572 (
            .O(N__12973),
            .I(N__12964));
    LocalMux I__1571 (
            .O(N__12964),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    CascadeMux I__1570 (
            .O(N__12961),
            .I(N__12958));
    InMux I__1569 (
            .O(N__12958),
            .I(N__12955));
    LocalMux I__1568 (
            .O(N__12955),
            .I(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ));
    CascadeMux I__1567 (
            .O(N__12952),
            .I(N__12949));
    InMux I__1566 (
            .O(N__12949),
            .I(N__12946));
    LocalMux I__1565 (
            .O(N__12946),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ));
    CascadeMux I__1564 (
            .O(N__12943),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ));
    CascadeMux I__1563 (
            .O(N__12940),
            .I(N__12937));
    InMux I__1562 (
            .O(N__12937),
            .I(N__12934));
    LocalMux I__1561 (
            .O(N__12934),
            .I(N__12931));
    Odrv4 I__1560 (
            .O(N__12931),
            .I(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ));
    InMux I__1559 (
            .O(N__12928),
            .I(N__12925));
    LocalMux I__1558 (
            .O(N__12925),
            .I(N__12922));
    Odrv4 I__1557 (
            .O(N__12922),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    CascadeMux I__1556 (
            .O(N__12919),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    InMux I__1555 (
            .O(N__12916),
            .I(N__12913));
    LocalMux I__1554 (
            .O(N__12913),
            .I(N__12910));
    Odrv12 I__1553 (
            .O(N__12910),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__1552 (
            .O(N__12907),
            .I(N__12904));
    LocalMux I__1551 (
            .O(N__12904),
            .I(N__12901));
    Span4Mux_v I__1550 (
            .O(N__12901),
            .I(N__12897));
    InMux I__1549 (
            .O(N__12900),
            .I(N__12894));
    Span4Mux_v I__1548 (
            .O(N__12897),
            .I(N__12889));
    LocalMux I__1547 (
            .O(N__12894),
            .I(N__12889));
    Span4Mux_v I__1546 (
            .O(N__12889),
            .I(N__12886));
    Span4Mux_v I__1545 (
            .O(N__12886),
            .I(N__12883));
    Odrv4 I__1544 (
            .O(N__12883),
            .I(throttle_command_2));
    InMux I__1543 (
            .O(N__12880),
            .I(N__12877));
    LocalMux I__1542 (
            .O(N__12877),
            .I(N__12874));
    Odrv4 I__1541 (
            .O(N__12874),
            .I(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ));
    CascadeMux I__1540 (
            .O(N__12871),
            .I(\ppm_encoder_1.PPM_STATE_58_d_cascade_ ));
    InMux I__1539 (
            .O(N__12868),
            .I(N__12860));
    InMux I__1538 (
            .O(N__12867),
            .I(N__12860));
    InMux I__1537 (
            .O(N__12866),
            .I(N__12855));
    InMux I__1536 (
            .O(N__12865),
            .I(N__12855));
    LocalMux I__1535 (
            .O(N__12860),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__1534 (
            .O(N__12855),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__1533 (
            .O(N__12850),
            .I(N__12846));
    CascadeMux I__1532 (
            .O(N__12849),
            .I(N__12843));
    LocalMux I__1531 (
            .O(N__12846),
            .I(N__12839));
    InMux I__1530 (
            .O(N__12843),
            .I(N__12834));
    InMux I__1529 (
            .O(N__12842),
            .I(N__12834));
    Odrv4 I__1528 (
            .O(N__12839),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__1527 (
            .O(N__12834),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__1526 (
            .O(N__12829),
            .I(N__12825));
    CascadeMux I__1525 (
            .O(N__12828),
            .I(N__12822));
    InMux I__1524 (
            .O(N__12825),
            .I(N__12818));
    InMux I__1523 (
            .O(N__12822),
            .I(N__12813));
    InMux I__1522 (
            .O(N__12821),
            .I(N__12813));
    LocalMux I__1521 (
            .O(N__12818),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__1520 (
            .O(N__12813),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__1519 (
            .O(N__12808),
            .I(N__12803));
    InMux I__1518 (
            .O(N__12807),
            .I(N__12800));
    InMux I__1517 (
            .O(N__12806),
            .I(N__12797));
    LocalMux I__1516 (
            .O(N__12803),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__1515 (
            .O(N__12800),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__1514 (
            .O(N__12797),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    InMux I__1513 (
            .O(N__12790),
            .I(N__12786));
    InMux I__1512 (
            .O(N__12789),
            .I(N__12783));
    LocalMux I__1511 (
            .O(N__12786),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    LocalMux I__1510 (
            .O(N__12783),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    CascadeMux I__1509 (
            .O(N__12778),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ));
    InMux I__1508 (
            .O(N__12775),
            .I(N__12771));
    InMux I__1507 (
            .O(N__12774),
            .I(N__12768));
    LocalMux I__1506 (
            .O(N__12771),
            .I(N__12765));
    LocalMux I__1505 (
            .O(N__12768),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv4 I__1504 (
            .O(N__12765),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    CascadeMux I__1503 (
            .O(N__12760),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    CascadeMux I__1502 (
            .O(N__12757),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    InMux I__1501 (
            .O(N__12754),
            .I(N__12751));
    LocalMux I__1500 (
            .O(N__12751),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    CascadeMux I__1499 (
            .O(N__12748),
            .I(N__12745));
    InMux I__1498 (
            .O(N__12745),
            .I(N__12740));
    InMux I__1497 (
            .O(N__12744),
            .I(N__12737));
    InMux I__1496 (
            .O(N__12743),
            .I(N__12734));
    LocalMux I__1495 (
            .O(N__12740),
            .I(N__12731));
    LocalMux I__1494 (
            .O(N__12737),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    LocalMux I__1493 (
            .O(N__12734),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv4 I__1492 (
            .O(N__12731),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__1491 (
            .O(N__12724),
            .I(N__12719));
    InMux I__1490 (
            .O(N__12723),
            .I(N__12714));
    InMux I__1489 (
            .O(N__12722),
            .I(N__12714));
    LocalMux I__1488 (
            .O(N__12719),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    LocalMux I__1487 (
            .O(N__12714),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    CascadeMux I__1486 (
            .O(N__12709),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ));
    CascadeMux I__1485 (
            .O(N__12706),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    InMux I__1484 (
            .O(N__12703),
            .I(N__12700));
    LocalMux I__1483 (
            .O(N__12700),
            .I(N__12696));
    InMux I__1482 (
            .O(N__12699),
            .I(N__12693));
    Span4Mux_v I__1481 (
            .O(N__12696),
            .I(N__12688));
    LocalMux I__1480 (
            .O(N__12693),
            .I(N__12688));
    Span4Mux_v I__1479 (
            .O(N__12688),
            .I(N__12685));
    Span4Mux_v I__1478 (
            .O(N__12685),
            .I(N__12682));
    Odrv4 I__1477 (
            .O(N__12682),
            .I(throttle_command_1));
    InMux I__1476 (
            .O(N__12679),
            .I(N__12676));
    LocalMux I__1475 (
            .O(N__12676),
            .I(N__12673));
    Odrv12 I__1474 (
            .O(N__12673),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__1473 (
            .O(N__12670),
            .I(N__12667));
    LocalMux I__1472 (
            .O(N__12667),
            .I(N__12663));
    InMux I__1471 (
            .O(N__12666),
            .I(N__12660));
    Span4Mux_h I__1470 (
            .O(N__12663),
            .I(N__12657));
    LocalMux I__1469 (
            .O(N__12660),
            .I(N__12654));
    Sp12to4 I__1468 (
            .O(N__12657),
            .I(N__12649));
    Span12Mux_h I__1467 (
            .O(N__12654),
            .I(N__12649));
    Odrv12 I__1466 (
            .O(N__12649),
            .I(throttle_command_10));
    InMux I__1465 (
            .O(N__12646),
            .I(N__12643));
    LocalMux I__1464 (
            .O(N__12643),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__1463 (
            .O(N__12640),
            .I(N__12636));
    InMux I__1462 (
            .O(N__12639),
            .I(N__12633));
    LocalMux I__1461 (
            .O(N__12636),
            .I(N__12628));
    LocalMux I__1460 (
            .O(N__12633),
            .I(N__12628));
    Span4Mux_v I__1459 (
            .O(N__12628),
            .I(N__12625));
    Span4Mux_v I__1458 (
            .O(N__12625),
            .I(N__12622));
    Span4Mux_v I__1457 (
            .O(N__12622),
            .I(N__12619));
    Odrv4 I__1456 (
            .O(N__12619),
            .I(throttle_command_13));
    InMux I__1455 (
            .O(N__12616),
            .I(N__12613));
    LocalMux I__1454 (
            .O(N__12613),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__1453 (
            .O(N__12610),
            .I(N__12607));
    LocalMux I__1452 (
            .O(N__12607),
            .I(N__12603));
    InMux I__1451 (
            .O(N__12606),
            .I(N__12600));
    Span4Mux_v I__1450 (
            .O(N__12603),
            .I(N__12595));
    LocalMux I__1449 (
            .O(N__12600),
            .I(N__12595));
    Span4Mux_v I__1448 (
            .O(N__12595),
            .I(N__12592));
    Odrv4 I__1447 (
            .O(N__12592),
            .I(throttle_command_4));
    InMux I__1446 (
            .O(N__12589),
            .I(N__12586));
    LocalMux I__1445 (
            .O(N__12586),
            .I(N__12583));
    Odrv4 I__1444 (
            .O(N__12583),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__1443 (
            .O(N__12580),
            .I(N__12577));
    LocalMux I__1442 (
            .O(N__12577),
            .I(N__12574));
    Odrv4 I__1441 (
            .O(N__12574),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__1440 (
            .O(N__12571),
            .I(N__12568));
    LocalMux I__1439 (
            .O(N__12568),
            .I(N__12564));
    InMux I__1438 (
            .O(N__12567),
            .I(N__12561));
    Span4Mux_v I__1437 (
            .O(N__12564),
            .I(N__12556));
    LocalMux I__1436 (
            .O(N__12561),
            .I(N__12556));
    Span4Mux_v I__1435 (
            .O(N__12556),
            .I(N__12553));
    Span4Mux_v I__1434 (
            .O(N__12553),
            .I(N__12550));
    Odrv4 I__1433 (
            .O(N__12550),
            .I(throttle_command_5));
    InMux I__1432 (
            .O(N__12547),
            .I(N__12544));
    LocalMux I__1431 (
            .O(N__12544),
            .I(N__12540));
    InMux I__1430 (
            .O(N__12543),
            .I(N__12537));
    Span4Mux_v I__1429 (
            .O(N__12540),
            .I(N__12534));
    LocalMux I__1428 (
            .O(N__12537),
            .I(N__12531));
    Span4Mux_v I__1427 (
            .O(N__12534),
            .I(N__12526));
    Span4Mux_v I__1426 (
            .O(N__12531),
            .I(N__12526));
    Span4Mux_v I__1425 (
            .O(N__12526),
            .I(N__12523));
    Odrv4 I__1424 (
            .O(N__12523),
            .I(throttle_command_8));
    InMux I__1423 (
            .O(N__12520),
            .I(N__12517));
    LocalMux I__1422 (
            .O(N__12517),
            .I(N__12514));
    Odrv4 I__1421 (
            .O(N__12514),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__1420 (
            .O(N__12511),
            .I(N__12508));
    LocalMux I__1419 (
            .O(N__12508),
            .I(N__12505));
    Odrv4 I__1418 (
            .O(N__12505),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__1417 (
            .O(N__12502),
            .I(N__12499));
    LocalMux I__1416 (
            .O(N__12499),
            .I(N__12495));
    InMux I__1415 (
            .O(N__12498),
            .I(N__12492));
    Span4Mux_v I__1414 (
            .O(N__12495),
            .I(N__12487));
    LocalMux I__1413 (
            .O(N__12492),
            .I(N__12487));
    Span4Mux_v I__1412 (
            .O(N__12487),
            .I(N__12484));
    Span4Mux_v I__1411 (
            .O(N__12484),
            .I(N__12481));
    Odrv4 I__1410 (
            .O(N__12481),
            .I(throttle_command_7));
    InMux I__1409 (
            .O(N__12478),
            .I(N__12474));
    InMux I__1408 (
            .O(N__12477),
            .I(N__12471));
    LocalMux I__1407 (
            .O(N__12474),
            .I(N__12466));
    LocalMux I__1406 (
            .O(N__12471),
            .I(N__12466));
    Span4Mux_v I__1405 (
            .O(N__12466),
            .I(N__12463));
    Span4Mux_v I__1404 (
            .O(N__12463),
            .I(N__12460));
    Odrv4 I__1403 (
            .O(N__12460),
            .I(throttle_command_6));
    InMux I__1402 (
            .O(N__12457),
            .I(N__12454));
    LocalMux I__1401 (
            .O(N__12454),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    InMux I__1400 (
            .O(N__12451),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__1399 (
            .O(N__12448),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__1398 (
            .O(N__12445),
            .I(bfn_2_20_0_));
    InMux I__1397 (
            .O(N__12442),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__1396 (
            .O(N__12439),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__1395 (
            .O(N__12436),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__1394 (
            .O(N__12433),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__1393 (
            .O(N__12430),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__1392 (
            .O(N__12427),
            .I(N__12424));
    LocalMux I__1391 (
            .O(N__12424),
            .I(N__12421));
    Span4Mux_v I__1390 (
            .O(N__12421),
            .I(N__12418));
    Span4Mux_v I__1389 (
            .O(N__12418),
            .I(N__12415));
    Odrv4 I__1388 (
            .O(N__12415),
            .I(throttle_command_14));
    InMux I__1387 (
            .O(N__12412),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    InMux I__1386 (
            .O(N__12409),
            .I(N__12406));
    LocalMux I__1385 (
            .O(N__12406),
            .I(drone_altitude_i_9));
    InMux I__1384 (
            .O(N__12403),
            .I(N__12400));
    LocalMux I__1383 (
            .O(N__12400),
            .I(drone_altitude_14));
    InMux I__1382 (
            .O(N__12397),
            .I(N__12394));
    LocalMux I__1381 (
            .O(N__12394),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    InMux I__1380 (
            .O(N__12391),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__1379 (
            .O(N__12388),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__1378 (
            .O(N__12385),
            .I(N__12381));
    InMux I__1377 (
            .O(N__12384),
            .I(N__12378));
    LocalMux I__1376 (
            .O(N__12381),
            .I(N__12375));
    LocalMux I__1375 (
            .O(N__12378),
            .I(N__12372));
    Span12Mux_s11_v I__1374 (
            .O(N__12375),
            .I(N__12367));
    Span12Mux_h I__1373 (
            .O(N__12372),
            .I(N__12367));
    Odrv12 I__1372 (
            .O(N__12367),
            .I(throttle_command_3));
    InMux I__1371 (
            .O(N__12364),
            .I(N__12361));
    LocalMux I__1370 (
            .O(N__12361),
            .I(N__12358));
    Span4Mux_v I__1369 (
            .O(N__12358),
            .I(N__12355));
    Odrv4 I__1368 (
            .O(N__12355),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__1367 (
            .O(N__12352),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__1366 (
            .O(N__12349),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__1365 (
            .O(N__12346),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    CascadeMux I__1364 (
            .O(N__12343),
            .I(N__12339));
    CascadeMux I__1363 (
            .O(N__12342),
            .I(N__12336));
    InMux I__1362 (
            .O(N__12339),
            .I(N__12333));
    InMux I__1361 (
            .O(N__12336),
            .I(N__12330));
    LocalMux I__1360 (
            .O(N__12333),
            .I(alt_command_3));
    LocalMux I__1359 (
            .O(N__12330),
            .I(alt_command_3));
    CascadeMux I__1358 (
            .O(N__12325),
            .I(N__12321));
    InMux I__1357 (
            .O(N__12324),
            .I(N__12318));
    InMux I__1356 (
            .O(N__12321),
            .I(N__12315));
    LocalMux I__1355 (
            .O(N__12318),
            .I(alt_command_1));
    LocalMux I__1354 (
            .O(N__12315),
            .I(alt_command_1));
    CascadeMux I__1353 (
            .O(N__12310),
            .I(\Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_ ));
    CascadeMux I__1352 (
            .O(N__12307),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    CascadeMux I__1351 (
            .O(N__12304),
            .I(N__12300));
    InMux I__1350 (
            .O(N__12303),
            .I(N__12297));
    InMux I__1349 (
            .O(N__12300),
            .I(N__12294));
    LocalMux I__1348 (
            .O(N__12297),
            .I(alt_command_0));
    LocalMux I__1347 (
            .O(N__12294),
            .I(alt_command_0));
    InMux I__1346 (
            .O(N__12289),
            .I(N__12280));
    InMux I__1345 (
            .O(N__12288),
            .I(N__12280));
    InMux I__1344 (
            .O(N__12287),
            .I(N__12280));
    LocalMux I__1343 (
            .O(N__12280),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    CascadeMux I__1342 (
            .O(N__12277),
            .I(N__12274));
    InMux I__1341 (
            .O(N__12274),
            .I(N__12270));
    InMux I__1340 (
            .O(N__12273),
            .I(N__12267));
    LocalMux I__1339 (
            .O(N__12270),
            .I(N__12264));
    LocalMux I__1338 (
            .O(N__12267),
            .I(alt_command_2));
    Odrv4 I__1337 (
            .O(N__12264),
            .I(alt_command_2));
    InMux I__1336 (
            .O(N__12259),
            .I(N__12256));
    LocalMux I__1335 (
            .O(N__12256),
            .I(\Commands_frame_decoder.source_CH1data8lt7_0 ));
    InMux I__1334 (
            .O(N__12253),
            .I(N__12250));
    LocalMux I__1333 (
            .O(N__12250),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__1332 (
            .O(N__12247),
            .I(N__12244));
    LocalMux I__1331 (
            .O(N__12244),
            .I(drone_altitude_i_8));
    InMux I__1330 (
            .O(N__12241),
            .I(N__12238));
    LocalMux I__1329 (
            .O(N__12238),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__1328 (
            .O(N__12235),
            .I(N__12232));
    LocalMux I__1327 (
            .O(N__12232),
            .I(drone_altitude_i_6));
    InMux I__1326 (
            .O(N__12229),
            .I(N__12226));
    LocalMux I__1325 (
            .O(N__12226),
            .I(drone_altitude_1));
    InMux I__1324 (
            .O(N__12223),
            .I(N__12220));
    LocalMux I__1323 (
            .O(N__12220),
            .I(\pid_alt.error_axbZ0Z_1 ));
    CascadeMux I__1322 (
            .O(N__12217),
            .I(\dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_ ));
    CascadeMux I__1321 (
            .O(N__12214),
            .I(\dron_frame_decoder_1.source_Altitude8lt7_0_cascade_ ));
    InMux I__1320 (
            .O(N__12211),
            .I(N__12208));
    LocalMux I__1319 (
            .O(N__12208),
            .I(drone_altitude_2));
    InMux I__1318 (
            .O(N__12205),
            .I(N__12202));
    LocalMux I__1317 (
            .O(N__12202),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__1316 (
            .O(N__12199),
            .I(N__12188));
    InMux I__1315 (
            .O(N__12198),
            .I(N__12188));
    InMux I__1314 (
            .O(N__12197),
            .I(N__12188));
    InMux I__1313 (
            .O(N__12196),
            .I(N__12183));
    InMux I__1312 (
            .O(N__12195),
            .I(N__12183));
    LocalMux I__1311 (
            .O(N__12188),
            .I(\dron_frame_decoder_1.source_Altitude8lt7_0 ));
    LocalMux I__1310 (
            .O(N__12183),
            .I(\dron_frame_decoder_1.source_Altitude8lt7_0 ));
    InMux I__1309 (
            .O(N__12178),
            .I(N__12175));
    LocalMux I__1308 (
            .O(N__12175),
            .I(drone_altitude_3));
    InMux I__1307 (
            .O(N__12172),
            .I(N__12169));
    LocalMux I__1306 (
            .O(N__12169),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__1305 (
            .O(N__12166),
            .I(N__12163));
    LocalMux I__1304 (
            .O(N__12163),
            .I(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4 ));
    CascadeMux I__1303 (
            .O(N__12160),
            .I(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_ ));
    InMux I__1302 (
            .O(N__12157),
            .I(N__12154));
    LocalMux I__1301 (
            .O(N__12154),
            .I(\dron_frame_decoder_1.WDT10lto13_1 ));
    InMux I__1300 (
            .O(N__12151),
            .I(N__12148));
    LocalMux I__1299 (
            .O(N__12148),
            .I(\dron_frame_decoder_1.WDT10lt14_0 ));
    InMux I__1298 (
            .O(N__12145),
            .I(N__12140));
    InMux I__1297 (
            .O(N__12144),
            .I(N__12137));
    InMux I__1296 (
            .O(N__12143),
            .I(N__12134));
    LocalMux I__1295 (
            .O(N__12140),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__1294 (
            .O(N__12137),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__1293 (
            .O(N__12134),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    CascadeMux I__1292 (
            .O(N__12127),
            .I(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ));
    CascadeMux I__1291 (
            .O(N__12124),
            .I(N__12120));
    InMux I__1290 (
            .O(N__12123),
            .I(N__12116));
    InMux I__1289 (
            .O(N__12120),
            .I(N__12111));
    InMux I__1288 (
            .O(N__12119),
            .I(N__12111));
    LocalMux I__1287 (
            .O(N__12116),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__1286 (
            .O(N__12111),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    CascadeMux I__1285 (
            .O(N__12106),
            .I(N__12102));
    InMux I__1284 (
            .O(N__12105),
            .I(N__12099));
    InMux I__1283 (
            .O(N__12102),
            .I(N__12096));
    LocalMux I__1282 (
            .O(N__12099),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__1281 (
            .O(N__12096),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__1280 (
            .O(N__12091),
            .I(N__12088));
    LocalMux I__1279 (
            .O(N__12088),
            .I(N__12085));
    Span4Mux_s2_h I__1278 (
            .O(N__12085),
            .I(N__12081));
    InMux I__1277 (
            .O(N__12084),
            .I(N__12078));
    Odrv4 I__1276 (
            .O(N__12081),
            .I(drone_altitude_0));
    LocalMux I__1275 (
            .O(N__12078),
            .I(drone_altitude_0));
    InMux I__1274 (
            .O(N__12073),
            .I(N__12069));
    InMux I__1273 (
            .O(N__12072),
            .I(N__12066));
    LocalMux I__1272 (
            .O(N__12069),
            .I(\pid_alt.drone_altitude_i_0 ));
    LocalMux I__1271 (
            .O(N__12066),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__1270 (
            .O(N__12061),
            .I(N__12058));
    LocalMux I__1269 (
            .O(N__12058),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    InMux I__1268 (
            .O(N__12055),
            .I(N__12052));
    LocalMux I__1267 (
            .O(N__12052),
            .I(drone_altitude_i_4));
    InMux I__1266 (
            .O(N__12049),
            .I(N__12046));
    LocalMux I__1265 (
            .O(N__12046),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__1264 (
            .O(N__12043),
            .I(N__12040));
    LocalMux I__1263 (
            .O(N__12040),
            .I(drone_altitude_i_5));
    InMux I__1262 (
            .O(N__12037),
            .I(N__12034));
    LocalMux I__1261 (
            .O(N__12034),
            .I(N__12030));
    InMux I__1260 (
            .O(N__12033),
            .I(N__12027));
    Span4Mux_s2_h I__1259 (
            .O(N__12030),
            .I(N__12024));
    LocalMux I__1258 (
            .O(N__12027),
            .I(alt_kp_3));
    Odrv4 I__1257 (
            .O(N__12024),
            .I(alt_kp_3));
    CascadeMux I__1256 (
            .O(N__12019),
            .I(N__12015));
    InMux I__1255 (
            .O(N__12018),
            .I(N__12012));
    InMux I__1254 (
            .O(N__12015),
            .I(N__12009));
    LocalMux I__1253 (
            .O(N__12012),
            .I(N__12006));
    LocalMux I__1252 (
            .O(N__12009),
            .I(alt_kp_6));
    Odrv4 I__1251 (
            .O(N__12006),
            .I(alt_kp_6));
    SRMux I__1250 (
            .O(N__12001),
            .I(N__11997));
    SRMux I__1249 (
            .O(N__12000),
            .I(N__11994));
    LocalMux I__1248 (
            .O(N__11997),
            .I(N__11991));
    LocalMux I__1247 (
            .O(N__11994),
            .I(N__11988));
    Span4Mux_s2_h I__1246 (
            .O(N__11991),
            .I(N__11985));
    Span4Mux_s2_h I__1245 (
            .O(N__11988),
            .I(N__11982));
    Span4Mux_h I__1244 (
            .O(N__11985),
            .I(N__11979));
    Span4Mux_h I__1243 (
            .O(N__11982),
            .I(N__11976));
    Odrv4 I__1242 (
            .O(N__11979),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    Odrv4 I__1241 (
            .O(N__11976),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__1240 (
            .O(N__11971),
            .I(N__11967));
    InMux I__1239 (
            .O(N__11970),
            .I(N__11964));
    LocalMux I__1238 (
            .O(N__11967),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    LocalMux I__1237 (
            .O(N__11964),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__1236 (
            .O(N__11959),
            .I(N__11955));
    InMux I__1235 (
            .O(N__11958),
            .I(N__11952));
    LocalMux I__1234 (
            .O(N__11955),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__1233 (
            .O(N__11952),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__1232 (
            .O(N__11947),
            .I(N__11943));
    InMux I__1231 (
            .O(N__11946),
            .I(N__11940));
    LocalMux I__1230 (
            .O(N__11943),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    LocalMux I__1229 (
            .O(N__11940),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    CascadeMux I__1228 (
            .O(N__11935),
            .I(N__11931));
    InMux I__1227 (
            .O(N__11934),
            .I(N__11928));
    InMux I__1226 (
            .O(N__11931),
            .I(N__11925));
    LocalMux I__1225 (
            .O(N__11928),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__1224 (
            .O(N__11925),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__1223 (
            .O(N__11920),
            .I(N__11916));
    InMux I__1222 (
            .O(N__11919),
            .I(N__11913));
    LocalMux I__1221 (
            .O(N__11916),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    LocalMux I__1220 (
            .O(N__11913),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__1219 (
            .O(N__11908),
            .I(N__11903));
    InMux I__1218 (
            .O(N__11907),
            .I(N__11898));
    InMux I__1217 (
            .O(N__11906),
            .I(N__11898));
    LocalMux I__1216 (
            .O(N__11903),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__1215 (
            .O(N__11898),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__1214 (
            .O(N__11893),
            .I(N__11889));
    InMux I__1213 (
            .O(N__11892),
            .I(N__11886));
    LocalMux I__1212 (
            .O(N__11889),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__1211 (
            .O(N__11886),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    CascadeMux I__1210 (
            .O(N__11881),
            .I(N__11877));
    InMux I__1209 (
            .O(N__11880),
            .I(N__11874));
    InMux I__1208 (
            .O(N__11877),
            .I(N__11871));
    LocalMux I__1207 (
            .O(N__11874),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__1206 (
            .O(N__11871),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__1205 (
            .O(N__11866),
            .I(N__11861));
    InMux I__1204 (
            .O(N__11865),
            .I(N__11856));
    InMux I__1203 (
            .O(N__11864),
            .I(N__11856));
    LocalMux I__1202 (
            .O(N__11861),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__1201 (
            .O(N__11856),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__1200 (
            .O(N__11851),
            .I(N__11847));
    InMux I__1199 (
            .O(N__11850),
            .I(N__11844));
    LocalMux I__1198 (
            .O(N__11847),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    LocalMux I__1197 (
            .O(N__11844),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    InMux I__1196 (
            .O(N__11839),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__1195 (
            .O(N__11836),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__1194 (
            .O(N__11833),
            .I(bfn_1_30_0_));
    InMux I__1193 (
            .O(N__11830),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__1192 (
            .O(N__11827),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__1191 (
            .O(N__11824),
            .I(N__11821));
    LocalMux I__1190 (
            .O(N__11821),
            .I(N__11817));
    InMux I__1189 (
            .O(N__11820),
            .I(N__11814));
    Span4Mux_s2_h I__1188 (
            .O(N__11817),
            .I(N__11811));
    LocalMux I__1187 (
            .O(N__11814),
            .I(alt_kp_0));
    Odrv4 I__1186 (
            .O(N__11811),
            .I(alt_kp_0));
    InMux I__1185 (
            .O(N__11806),
            .I(N__11802));
    CascadeMux I__1184 (
            .O(N__11805),
            .I(N__11799));
    LocalMux I__1183 (
            .O(N__11802),
            .I(N__11796));
    InMux I__1182 (
            .O(N__11799),
            .I(N__11793));
    Span4Mux_s2_h I__1181 (
            .O(N__11796),
            .I(N__11790));
    LocalMux I__1180 (
            .O(N__11793),
            .I(alt_kp_2));
    Odrv4 I__1179 (
            .O(N__11790),
            .I(alt_kp_2));
    InMux I__1178 (
            .O(N__11785),
            .I(N__11782));
    LocalMux I__1177 (
            .O(N__11782),
            .I(N__11778));
    InMux I__1176 (
            .O(N__11781),
            .I(N__11775));
    Span4Mux_v I__1175 (
            .O(N__11778),
            .I(N__11772));
    LocalMux I__1174 (
            .O(N__11775),
            .I(alt_kp_1));
    Odrv4 I__1173 (
            .O(N__11772),
            .I(alt_kp_1));
    CEMux I__1172 (
            .O(N__11767),
            .I(N__11763));
    CEMux I__1171 (
            .O(N__11766),
            .I(N__11760));
    LocalMux I__1170 (
            .O(N__11763),
            .I(N__11755));
    LocalMux I__1169 (
            .O(N__11760),
            .I(N__11752));
    CEMux I__1168 (
            .O(N__11759),
            .I(N__11749));
    CEMux I__1167 (
            .O(N__11758),
            .I(N__11746));
    Span4Mux_s3_h I__1166 (
            .O(N__11755),
            .I(N__11743));
    Span4Mux_s3_h I__1165 (
            .O(N__11752),
            .I(N__11740));
    LocalMux I__1164 (
            .O(N__11749),
            .I(N__11737));
    LocalMux I__1163 (
            .O(N__11746),
            .I(N__11734));
    Odrv4 I__1162 (
            .O(N__11743),
            .I(\pid_alt.source_p_enZ0 ));
    Odrv4 I__1161 (
            .O(N__11740),
            .I(\pid_alt.source_p_enZ0 ));
    Odrv4 I__1160 (
            .O(N__11737),
            .I(\pid_alt.source_p_enZ0 ));
    Odrv12 I__1159 (
            .O(N__11734),
            .I(\pid_alt.source_p_enZ0 ));
    InMux I__1158 (
            .O(N__11725),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__1157 (
            .O(N__11722),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__1156 (
            .O(N__11719),
            .I(N__11716));
    LocalMux I__1155 (
            .O(N__11716),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__1154 (
            .O(N__11713),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__1153 (
            .O(N__11710),
            .I(bfn_1_29_0_));
    InMux I__1152 (
            .O(N__11707),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__1151 (
            .O(N__11704),
            .I(N__11701));
    LocalMux I__1150 (
            .O(N__11701),
            .I(N__11698));
    Odrv4 I__1149 (
            .O(N__11698),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__1148 (
            .O(N__11695),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__1147 (
            .O(N__11692),
            .I(N__11689));
    LocalMux I__1146 (
            .O(N__11689),
            .I(N__11686));
    Odrv12 I__1145 (
            .O(N__11686),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__1144 (
            .O(N__11683),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__1143 (
            .O(N__11680),
            .I(N__11677));
    LocalMux I__1142 (
            .O(N__11677),
            .I(N__11674));
    Span4Mux_v I__1141 (
            .O(N__11674),
            .I(N__11671));
    Odrv4 I__1140 (
            .O(N__11671),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__1139 (
            .O(N__11668),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__1138 (
            .O(N__11665),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    CascadeMux I__1137 (
            .O(N__11662),
            .I(N__11659));
    InMux I__1136 (
            .O(N__11659),
            .I(N__11656));
    LocalMux I__1135 (
            .O(N__11656),
            .I(N__11653));
    Odrv4 I__1134 (
            .O(N__11653),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ));
    InMux I__1133 (
            .O(N__11650),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__1132 (
            .O(N__11647),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    CascadeMux I__1131 (
            .O(N__11644),
            .I(N__11641));
    InMux I__1130 (
            .O(N__11641),
            .I(N__11638));
    LocalMux I__1129 (
            .O(N__11638),
            .I(N__11635));
    Odrv4 I__1128 (
            .O(N__11635),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__1127 (
            .O(N__11632),
            .I(N__11629));
    LocalMux I__1126 (
            .O(N__11629),
            .I(N__11626));
    Odrv4 I__1125 (
            .O(N__11626),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__1124 (
            .O(N__11623),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__1123 (
            .O(N__11620),
            .I(N__11617));
    LocalMux I__1122 (
            .O(N__11617),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__1121 (
            .O(N__11614),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    CascadeMux I__1120 (
            .O(N__11611),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ));
    CascadeMux I__1119 (
            .O(N__11608),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ));
    CascadeMux I__1118 (
            .O(N__11605),
            .I(N__11601));
    InMux I__1117 (
            .O(N__11604),
            .I(N__11596));
    InMux I__1116 (
            .O(N__11601),
            .I(N__11596));
    LocalMux I__1115 (
            .O(N__11596),
            .I(N__11593));
    Odrv12 I__1114 (
            .O(N__11593),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    InMux I__1113 (
            .O(N__11590),
            .I(N__11587));
    LocalMux I__1112 (
            .O(N__11587),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    InMux I__1111 (
            .O(N__11584),
            .I(N__11579));
    CascadeMux I__1110 (
            .O(N__11583),
            .I(N__11576));
    InMux I__1109 (
            .O(N__11582),
            .I(N__11573));
    LocalMux I__1108 (
            .O(N__11579),
            .I(N__11570));
    InMux I__1107 (
            .O(N__11576),
            .I(N__11567));
    LocalMux I__1106 (
            .O(N__11573),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv12 I__1105 (
            .O(N__11570),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    LocalMux I__1104 (
            .O(N__11567),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__1103 (
            .O(N__11560),
            .I(N__11557));
    LocalMux I__1102 (
            .O(N__11557),
            .I(N__11552));
    InMux I__1101 (
            .O(N__11556),
            .I(N__11547));
    InMux I__1100 (
            .O(N__11555),
            .I(N__11547));
    Odrv12 I__1099 (
            .O(N__11552),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    LocalMux I__1098 (
            .O(N__11547),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    CascadeMux I__1097 (
            .O(N__11542),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    CascadeMux I__1096 (
            .O(N__11539),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ));
    InMux I__1095 (
            .O(N__11536),
            .I(N__11533));
    LocalMux I__1094 (
            .O(N__11533),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13 ));
    CascadeMux I__1093 (
            .O(N__11530),
            .I(N__11525));
    InMux I__1092 (
            .O(N__11529),
            .I(N__11522));
    InMux I__1091 (
            .O(N__11528),
            .I(N__11519));
    InMux I__1090 (
            .O(N__11525),
            .I(N__11516));
    LocalMux I__1089 (
            .O(N__11522),
            .I(N__11511));
    LocalMux I__1088 (
            .O(N__11519),
            .I(N__11511));
    LocalMux I__1087 (
            .O(N__11516),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv12 I__1086 (
            .O(N__11511),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    CascadeMux I__1085 (
            .O(N__11506),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    InMux I__1084 (
            .O(N__11503),
            .I(N__11500));
    LocalMux I__1083 (
            .O(N__11500),
            .I(N__11497));
    Odrv12 I__1082 (
            .O(N__11497),
            .I(drone_altitude_i_7));
    InMux I__1081 (
            .O(N__11494),
            .I(N__11491));
    LocalMux I__1080 (
            .O(N__11491),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    CascadeMux I__1079 (
            .O(N__11488),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    InMux I__1078 (
            .O(N__11485),
            .I(N__11482));
    LocalMux I__1077 (
            .O(N__11482),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    InMux I__1076 (
            .O(N__11479),
            .I(N__11476));
    LocalMux I__1075 (
            .O(N__11476),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__1074 (
            .O(N__11473),
            .I(N__11470));
    LocalMux I__1073 (
            .O(N__11470),
            .I(drone_altitude_12));
    InMux I__1072 (
            .O(N__11467),
            .I(N__11464));
    LocalMux I__1071 (
            .O(N__11464),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__1070 (
            .O(N__11461),
            .I(N__11458));
    LocalMux I__1069 (
            .O(N__11458),
            .I(drone_altitude_13));
    InMux I__1068 (
            .O(N__11455),
            .I(N__11452));
    LocalMux I__1067 (
            .O(N__11452),
            .I(N__11449));
    Odrv4 I__1066 (
            .O(N__11449),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__1065 (
            .O(N__11446),
            .I(N__11443));
    LocalMux I__1064 (
            .O(N__11443),
            .I(N__11440));
    Odrv4 I__1063 (
            .O(N__11440),
            .I(drone_altitude_15));
    InMux I__1062 (
            .O(N__11437),
            .I(N__11434));
    LocalMux I__1061 (
            .O(N__11434),
            .I(N__11431));
    Span4Mux_s1_h I__1060 (
            .O(N__11431),
            .I(N__11428));
    Odrv4 I__1059 (
            .O(N__11428),
            .I(\pid_alt.error_10 ));
    InMux I__1058 (
            .O(N__11425),
            .I(\pid_alt.error_cry_9 ));
    InMux I__1057 (
            .O(N__11422),
            .I(N__11419));
    LocalMux I__1056 (
            .O(N__11419),
            .I(N__11416));
    Span4Mux_s1_h I__1055 (
            .O(N__11416),
            .I(N__11413));
    Odrv4 I__1054 (
            .O(N__11413),
            .I(\pid_alt.error_11 ));
    InMux I__1053 (
            .O(N__11410),
            .I(\pid_alt.error_cry_10 ));
    InMux I__1052 (
            .O(N__11407),
            .I(N__11404));
    LocalMux I__1051 (
            .O(N__11404),
            .I(N__11401));
    Span4Mux_s1_h I__1050 (
            .O(N__11401),
            .I(N__11398));
    Odrv4 I__1049 (
            .O(N__11398),
            .I(\pid_alt.error_12 ));
    InMux I__1048 (
            .O(N__11395),
            .I(\pid_alt.error_cry_11 ));
    InMux I__1047 (
            .O(N__11392),
            .I(N__11389));
    LocalMux I__1046 (
            .O(N__11389),
            .I(N__11386));
    Span4Mux_s1_h I__1045 (
            .O(N__11386),
            .I(N__11383));
    Odrv4 I__1044 (
            .O(N__11383),
            .I(\pid_alt.error_13 ));
    InMux I__1043 (
            .O(N__11380),
            .I(\pid_alt.error_cry_12 ));
    InMux I__1042 (
            .O(N__11377),
            .I(N__11374));
    LocalMux I__1041 (
            .O(N__11374),
            .I(N__11371));
    Span4Mux_v I__1040 (
            .O(N__11371),
            .I(N__11368));
    Odrv4 I__1039 (
            .O(N__11368),
            .I(\pid_alt.error_14 ));
    InMux I__1038 (
            .O(N__11365),
            .I(\pid_alt.error_cry_13 ));
    InMux I__1037 (
            .O(N__11362),
            .I(\pid_alt.error_cry_14 ));
    InMux I__1036 (
            .O(N__11359),
            .I(N__11356));
    LocalMux I__1035 (
            .O(N__11356),
            .I(N__11353));
    Span4Mux_v I__1034 (
            .O(N__11353),
            .I(N__11350));
    Odrv4 I__1033 (
            .O(N__11350),
            .I(\pid_alt.error_15 ));
    InMux I__1032 (
            .O(N__11347),
            .I(N__11344));
    LocalMux I__1031 (
            .O(N__11344),
            .I(drone_altitude_i_10));
    InMux I__1030 (
            .O(N__11341),
            .I(N__11338));
    LocalMux I__1029 (
            .O(N__11338),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__1028 (
            .O(N__11335),
            .I(N__11332));
    LocalMux I__1027 (
            .O(N__11332),
            .I(drone_altitude_i_11));
    InMux I__1026 (
            .O(N__11329),
            .I(N__11326));
    LocalMux I__1025 (
            .O(N__11326),
            .I(N__11323));
    Span4Mux_s1_h I__1024 (
            .O(N__11323),
            .I(N__11320));
    Odrv4 I__1023 (
            .O(N__11320),
            .I(\pid_alt.error_2 ));
    InMux I__1022 (
            .O(N__11317),
            .I(\pid_alt.error_cry_1 ));
    InMux I__1021 (
            .O(N__11314),
            .I(N__11311));
    LocalMux I__1020 (
            .O(N__11311),
            .I(N__11308));
    Span4Mux_s1_h I__1019 (
            .O(N__11308),
            .I(N__11305));
    Odrv4 I__1018 (
            .O(N__11305),
            .I(\pid_alt.error_3 ));
    InMux I__1017 (
            .O(N__11302),
            .I(\pid_alt.error_cry_2 ));
    InMux I__1016 (
            .O(N__11299),
            .I(N__11296));
    LocalMux I__1015 (
            .O(N__11296),
            .I(N__11293));
    Span4Mux_v I__1014 (
            .O(N__11293),
            .I(N__11290));
    Odrv4 I__1013 (
            .O(N__11290),
            .I(\pid_alt.error_4 ));
    InMux I__1012 (
            .O(N__11287),
            .I(\pid_alt.error_cry_3 ));
    InMux I__1011 (
            .O(N__11284),
            .I(N__11281));
    LocalMux I__1010 (
            .O(N__11281),
            .I(N__11278));
    Odrv4 I__1009 (
            .O(N__11278),
            .I(\pid_alt.error_5 ));
    InMux I__1008 (
            .O(N__11275),
            .I(\pid_alt.error_cry_4 ));
    InMux I__1007 (
            .O(N__11272),
            .I(N__11269));
    LocalMux I__1006 (
            .O(N__11269),
            .I(N__11266));
    Span4Mux_s1_h I__1005 (
            .O(N__11266),
            .I(N__11263));
    Odrv4 I__1004 (
            .O(N__11263),
            .I(\pid_alt.error_6 ));
    InMux I__1003 (
            .O(N__11260),
            .I(\pid_alt.error_cry_5 ));
    InMux I__1002 (
            .O(N__11257),
            .I(N__11254));
    LocalMux I__1001 (
            .O(N__11254),
            .I(N__11251));
    Span4Mux_s1_h I__1000 (
            .O(N__11251),
            .I(N__11248));
    Odrv4 I__999 (
            .O(N__11248),
            .I(\pid_alt.error_7 ));
    InMux I__998 (
            .O(N__11245),
            .I(\pid_alt.error_cry_6 ));
    InMux I__997 (
            .O(N__11242),
            .I(N__11239));
    LocalMux I__996 (
            .O(N__11239),
            .I(N__11236));
    Span4Mux_s2_h I__995 (
            .O(N__11236),
            .I(N__11233));
    Odrv4 I__994 (
            .O(N__11233),
            .I(\pid_alt.error_8 ));
    InMux I__993 (
            .O(N__11230),
            .I(bfn_1_16_0_));
    InMux I__992 (
            .O(N__11227),
            .I(N__11224));
    LocalMux I__991 (
            .O(N__11224),
            .I(N__11221));
    Span4Mux_v I__990 (
            .O(N__11221),
            .I(N__11218));
    Odrv4 I__989 (
            .O(N__11218),
            .I(\pid_alt.error_9 ));
    InMux I__988 (
            .O(N__11215),
            .I(\pid_alt.error_cry_8 ));
    InMux I__987 (
            .O(N__11212),
            .I(bfn_1_14_0_));
    InMux I__986 (
            .O(N__11209),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__985 (
            .O(N__11206),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__984 (
            .O(N__11203),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__983 (
            .O(N__11200),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    InMux I__982 (
            .O(N__11197),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__981 (
            .O(N__11194),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__980 (
            .O(N__11191),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    InMux I__979 (
            .O(N__11188),
            .I(N__11185));
    LocalMux I__978 (
            .O(N__11185),
            .I(N__11182));
    Span4Mux_s1_h I__977 (
            .O(N__11182),
            .I(N__11179));
    Odrv4 I__976 (
            .O(N__11179),
            .I(\pid_alt.error_1 ));
    InMux I__975 (
            .O(N__11176),
            .I(\pid_alt.error_cry_0 ));
    InMux I__974 (
            .O(N__11173),
            .I(N__11170));
    LocalMux I__973 (
            .O(N__11170),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__972 (
            .O(N__11167),
            .I(N__11164));
    LocalMux I__971 (
            .O(N__11164),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__970 (
            .O(N__11161),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__969 (
            .O(N__11158),
            .I(N__11155));
    LocalMux I__968 (
            .O(N__11155),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__967 (
            .O(N__11152),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__966 (
            .O(N__11149),
            .I(N__11146));
    LocalMux I__965 (
            .O(N__11146),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__964 (
            .O(N__11143),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__963 (
            .O(N__11140),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__962 (
            .O(N__11137),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__961 (
            .O(N__11134),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__960 (
            .O(N__11131),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__959 (
            .O(N__11128),
            .I(N__11125));
    LocalMux I__958 (
            .O(N__11125),
            .I(\pid_alt.O_11 ));
    InMux I__957 (
            .O(N__11122),
            .I(N__11119));
    LocalMux I__956 (
            .O(N__11119),
            .I(\pid_alt.O_13 ));
    InMux I__955 (
            .O(N__11116),
            .I(N__11113));
    LocalMux I__954 (
            .O(N__11113),
            .I(N__11110));
    Odrv4 I__953 (
            .O(N__11110),
            .I(\pid_alt.O_18 ));
    InMux I__952 (
            .O(N__11107),
            .I(N__11104));
    LocalMux I__951 (
            .O(N__11104),
            .I(\pid_alt.O_14 ));
    InMux I__950 (
            .O(N__11101),
            .I(N__11098));
    LocalMux I__949 (
            .O(N__11098),
            .I(\pid_alt.O_4 ));
    InMux I__948 (
            .O(N__11095),
            .I(N__11092));
    LocalMux I__947 (
            .O(N__11092),
            .I(\pid_alt.O_5 ));
    InMux I__946 (
            .O(N__11089),
            .I(N__11086));
    LocalMux I__945 (
            .O(N__11086),
            .I(\pid_alt.O_9 ));
    InMux I__944 (
            .O(N__11083),
            .I(N__11080));
    LocalMux I__943 (
            .O(N__11080),
            .I(\pid_alt.O_15 ));
    InMux I__942 (
            .O(N__11077),
            .I(N__11074));
    LocalMux I__941 (
            .O(N__11074),
            .I(\pid_alt.O_8 ));
    InMux I__940 (
            .O(N__11071),
            .I(N__11068));
    LocalMux I__939 (
            .O(N__11068),
            .I(N__11065));
    Odrv4 I__938 (
            .O(N__11065),
            .I(\pid_alt.O_17 ));
    InMux I__937 (
            .O(N__11062),
            .I(N__11059));
    LocalMux I__936 (
            .O(N__11059),
            .I(\pid_alt.O_6 ));
    InMux I__935 (
            .O(N__11056),
            .I(N__11053));
    LocalMux I__934 (
            .O(N__11053),
            .I(\pid_alt.O_7 ));
    InMux I__933 (
            .O(N__11050),
            .I(N__11047));
    LocalMux I__932 (
            .O(N__11047),
            .I(N__11044));
    Odrv4 I__931 (
            .O(N__11044),
            .I(\pid_alt.O_10 ));
    InMux I__930 (
            .O(N__11041),
            .I(N__11038));
    LocalMux I__929 (
            .O(N__11038),
            .I(N__11035));
    Odrv4 I__928 (
            .O(N__11035),
            .I(\pid_alt.O_16 ));
    InMux I__927 (
            .O(N__11032),
            .I(N__11029));
    LocalMux I__926 (
            .O(N__11029),
            .I(\pid_alt.O_12 ));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\scaler_3.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\scaler_3.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\scaler_2.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\scaler_2.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_13 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_13 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_3_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_3_27_0_));
    defparam IN_MUX_bfv_1_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_28_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_4_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_29_0_));
    defparam IN_MUX_bfv_4_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_30_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_4_30_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_7_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_29_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_7_29_0_));
    defparam IN_MUX_bfv_7_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_7_30_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_4_19_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__26679),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB pc_frame_decoder_dv_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__26833),
            .GLOBALBUFFEROUTPUT(pc_frame_decoder_dv_0_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__18883),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_168_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.source_p_ess_13_LC_1_9_0 .C_ON=1'b0;
    defparam \pid_alt.source_p_ess_13_LC_1_9_0 .SEQ_MODE=4'b1001;
    defparam \pid_alt.source_p_ess_13_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_p_ess_13_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11071),
            .lcout(throttle_command_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__11766),
            .sr(N__28714));
    defparam \pid_alt.source_p_ess_2_LC_1_9_1 .C_ON=1'b0;
    defparam \pid_alt.source_p_ess_2_LC_1_9_1 .SEQ_MODE=4'b1001;
    defparam \pid_alt.source_p_ess_2_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_p_ess_2_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11062),
            .lcout(throttle_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__11766),
            .sr(N__28714));
    defparam \pid_alt.source_p_ess_3_LC_1_9_2 .C_ON=1'b0;
    defparam \pid_alt.source_p_ess_3_LC_1_9_2 .SEQ_MODE=4'b1001;
    defparam \pid_alt.source_p_ess_3_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_p_ess_3_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11056),
            .lcout(throttle_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__11766),
            .sr(N__28714));
    defparam \pid_alt.source_p_ess_6_LC_1_9_3 .C_ON=1'b0;
    defparam \pid_alt.source_p_ess_6_LC_1_9_3 .SEQ_MODE=4'b1001;
    defparam \pid_alt.source_p_ess_6_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_p_ess_6_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11050),
            .lcout(throttle_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__11766),
            .sr(N__28714));
    defparam \pid_alt.source_p_9_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.source_p_9_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_9_LC_1_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_alt.source_p_9_LC_1_10_0  (
            .in0(N__28954),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11041),
            .lcout(throttle_command_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(N__11758),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_5_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.source_p_5_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_5_LC_1_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_5_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__28951),
            .in2(_gnd_net_),
            .in3(N__11032),
            .lcout(throttle_command_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(N__11758),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_4_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.source_p_4_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_4_LC_1_10_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_alt.source_p_4_LC_1_10_2  (
            .in0(N__28953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11128),
            .lcout(throttle_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(N__11758),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_1_6_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.source_p_1_6_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_1_6_LC_1_10_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_1_6_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__28950),
            .in2(_gnd_net_),
            .in3(N__11122),
            .lcout(throttle_command_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(N__11758),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_10_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.source_p_10_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_10_LC_1_10_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_alt.source_p_10_LC_1_10_4  (
            .in0(N__28952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11116),
            .lcout(throttle_command_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(N__11758),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_7_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.source_p_7_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_7_LC_1_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_7_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__28956),
            .in2(_gnd_net_),
            .in3(N__11107),
            .lcout(throttle_command_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(N__11759),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_0_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.source_p_0_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_0_LC_1_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_alt.source_p_0_LC_1_11_4  (
            .in0(N__28958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11101),
            .lcout(throttle_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(N__11759),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_1_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.source_p_1_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_1_LC_1_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_1_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__28955),
            .in2(_gnd_net_),
            .in3(N__11095),
            .lcout(throttle_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(N__11759),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_1_3_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.source_p_1_3_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_1_3_LC_1_11_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \pid_alt.source_p_1_3_LC_1_11_6  (
            .in0(N__28959),
            .in1(N__11089),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(throttle_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(N__11759),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_8_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.source_p_8_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_8_LC_1_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__28957),
            .in2(_gnd_net_),
            .in3(N__11083),
            .lcout(throttle_command_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(N__11759),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_1_2_LC_1_12_5 .C_ON=1'b0;
    defparam \pid_alt.source_p_1_2_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_p_1_2_LC_1_12_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.source_p_1_2_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__28963),
            .in2(_gnd_net_),
            .in3(N__11077),
            .lcout(throttle_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29381),
            .ce(N__11767),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_1_13_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_1_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__11173),
            .in2(N__12106),
            .in3(N__12105),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_1_LC_1_13_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_1_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__11167),
            .in2(_gnd_net_),
            .in3(N__11161),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_2_LC_1_13_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_1_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__11158),
            .in2(_gnd_net_),
            .in3(N__11152),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_3_LC_1_13_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_1_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__11149),
            .in2(_gnd_net_),
            .in3(N__11143),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_4_LC_1_13_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_1_13_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_1_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__11920),
            .in2(_gnd_net_),
            .in3(N__11140),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_5_LC_1_13_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_1_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__11947),
            .in2(_gnd_net_),
            .in3(N__11137),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_6_LC_1_13_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_1_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__11971),
            .in2(_gnd_net_),
            .in3(N__11134),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_7_LC_1_13_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_1_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__11851),
            .in2(_gnd_net_),
            .in3(N__11131),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__29378),
            .ce(),
            .sr(N__12000));
    defparam \dron_frame_decoder_1.WDT_8_LC_1_14_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_1_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__11959),
            .in2(_gnd_net_),
            .in3(N__11212),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_9_LC_1_14_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__11934),
            .in2(_gnd_net_),
            .in3(N__11209),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_10_LC_1_14_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_1_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__11893),
            .in2(_gnd_net_),
            .in3(N__11206),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_11_LC_1_14_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__11866),
            .in2(_gnd_net_),
            .in3(N__11203),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_12_LC_1_14_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__11908),
            .in2(_gnd_net_),
            .in3(N__11200),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_13_LC_1_14_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_1_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__11880),
            .in2(_gnd_net_),
            .in3(N__11197),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_14_LC_1_14_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_1_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__12123),
            .in2(_gnd_net_),
            .in3(N__11194),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \dron_frame_decoder_1.WDT_15_LC_1_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_1_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__12145),
            .in2(_gnd_net_),
            .in3(N__11191),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29375),
            .ce(),
            .sr(N__12001));
    defparam \pid_alt.error_cry_0_c_LC_1_15_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_1_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__12072),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_1_15_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__12223),
            .in2(_gnd_net_),
            .in3(N__11176),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_1_15_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__12205),
            .in2(_gnd_net_),
            .in3(N__11317),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_1_15_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__12172),
            .in2(_gnd_net_),
            .in3(N__11302),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_1_15_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__12055),
            .in2(N__12304),
            .in3(N__11287),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_1_15_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__12043),
            .in2(N__12325),
            .in3(N__11275),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_1_15_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_1_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__12235),
            .in2(N__12277),
            .in3(N__11260),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_1_15_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_1_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__11503),
            .in2(N__12342),
            .in3(N__11245),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_1_16_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_1_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__12247),
            .in2(N__13327),
            .in3(N__11230),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_1_16_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_1_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__12409),
            .in2(N__13315),
            .in3(N__11215),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_1_16_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_1_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__11347),
            .in2(N__13303),
            .in3(N__11425),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_1_16_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_1_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__11335),
            .in2(N__13738),
            .in3(N__11410),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_1_16_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_1_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__11479),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_1_16_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_1_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__11467),
            .in2(_gnd_net_),
            .in3(N__11380),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_1_16_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_1_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__11455),
            .in2(_gnd_net_),
            .in3(N__11365),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_1_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(N__11446),
            .in2(_gnd_net_),
            .in3(N__11362),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_1_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_1_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11341),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_1_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_1_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_1_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15289),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29363),
            .ce(N__13568),
            .sr(N__28750));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_1_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_1_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11485),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_1_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_1_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_1_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15256),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29363),
            .ce(N__13568),
            .sr(N__28750));
    defparam \pid_alt.error_axb_12_LC_1_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_1_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11473),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_1_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_1_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_1_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15192),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29363),
            .ce(N__13568),
            .sr(N__28750));
    defparam \pid_alt.error_axb_13_LC_1_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11461),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_1_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_1_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_1_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15132),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29363),
            .ce(N__13568),
            .sr(N__28750));
    defparam \pid_alt.error_axb_14_LC_1_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_1_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12403),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_1_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_1_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_1_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15015),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29357),
            .ce(N__13572),
            .sr(N__28756));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_1_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_1_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_1_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14847),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29357),
            .ce(N__13572),
            .sr(N__28756));
    defparam \ppm_encoder_1.throttle_6_LC_1_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_1_19_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_1_19_2 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_1_19_2  (
            .in0(N__12457),
            .in1(N__12478),
            .in2(N__11530),
            .in3(N__24864),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29350),
            .ce(),
            .sr(N__28763));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_1_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_1_19_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__11494),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_1_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_1_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15014),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29345),
            .ce(N__13722),
            .sr(N__28769));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_1_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_1_21_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_1_21_6  (
            .in0(N__22772),
            .in1(N__11529),
            .in2(_gnd_net_),
            .in3(N__11560),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_1_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_1_21_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(N__20959),
            .in2(N__11488),
            .in3(N__11584),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_1_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_1_22_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_1_22_0  (
            .in0(N__22761),
            .in1(N__13866),
            .in2(_gnd_net_),
            .in3(N__19801),
            .lcout(\ppm_encoder_1.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_1_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_1_22_6 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_1_22_6  (
            .in0(N__22762),
            .in1(N__28964),
            .in2(N__20980),
            .in3(N__23732),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29332),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_1_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_1_22_7 .LUT_INIT=16'b1111010011110110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_1_22_7  (
            .in0(N__23731),
            .in1(N__17818),
            .in2(N__28979),
            .in3(N__20773),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29332),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_1_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_1_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_1_23_0 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_1_23_0  (
            .in0(N__18562),
            .in1(N__28968),
            .in2(N__20979),
            .in3(N__23617),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29325),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_23_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_23_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_23_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_1_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_1_23_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_1_23_2  (
            .in0(N__18561),
            .in1(N__17801),
            .in2(N__20572),
            .in3(N__17857),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_158_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_1_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_1_23_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_1_23_4  (
            .in0(N__16150),
            .in1(N__23613),
            .in2(_gnd_net_),
            .in3(N__20782),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_1_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_1_23_5 .LUT_INIT=16'b0100000010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_1_23_5  (
            .in0(N__17858),
            .in1(N__22798),
            .in2(N__20972),
            .in3(N__20568),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_1_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_1_23_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_1_23_6  (
            .in0(N__20067),
            .in1(N__23612),
            .in2(_gnd_net_),
            .in3(N__20781),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_1_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_1_23_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_12_LC_1_23_7  (
            .in0(N__20783),
            .in1(_gnd_net_),
            .in2(N__23724),
            .in3(N__20066),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_1_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_1_24_0 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \ppm_encoder_1.elevator_RNI47DH2_13_LC_1_24_0  (
            .in0(N__15965),
            .in1(N__25006),
            .in2(N__16054),
            .in3(N__20095),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_1_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_1_24_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIKVRT5_13_LC_1_24_1  (
            .in0(N__16351),
            .in1(_gnd_net_),
            .in2(N__11539),
            .in3(N__11536),
            .lcout(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_1_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_1_24_2 .LUT_INIT=16'b1111010100110001;
    LogicCell40 \ppm_encoder_1.throttle_RNIK8JI2_13_LC_1_24_2  (
            .in0(N__15845),
            .in1(N__15726),
            .in2(N__20136),
            .in3(N__21016),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_1_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_1_24_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIO1KK2_6_LC_1_24_3  (
            .in0(N__11528),
            .in1(N__21072),
            .in2(N__15745),
            .in3(N__15844),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_1_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_1_24_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEDI96_6_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(N__18361),
            .in2(N__11506),
            .in3(N__11590),
            .lcout(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_1_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_1_24_5 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNI8GVN2_6_LC_1_24_5  (
            .in0(N__11555),
            .in1(N__15964),
            .in2(N__11583),
            .in3(N__16031),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_1_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_1_24_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_1_24_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_1_24_6  (
            .in0(N__11582),
            .in1(N__24954),
            .in2(_gnd_net_),
            .in3(N__24172),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29314),
            .ce(),
            .sr(N__28782));
    defparam \ppm_encoder_1.elevator_6_LC_1_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_1_24_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_1_24_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_1_24_7  (
            .in0(N__11556),
            .in1(N__24955),
            .in2(_gnd_net_),
            .in3(N__25996),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29314),
            .ce(),
            .sr(N__28782));
    defparam \ppm_encoder_1.init_pulses_3_LC_1_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_1_25_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_1_25_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_1_25_0  (
            .in0(N__18250),
            .in1(N__11632),
            .in2(N__18062),
            .in3(N__14041),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29306),
            .ce(),
            .sr(N__28786));
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_1_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_1_25_1 .LUT_INIT=16'b1001101001100101;
    LogicCell40 \ppm_encoder_1.throttle_RNIT9352_3_LC_1_25_1  (
            .in0(N__18461),
            .in1(N__18629),
            .in2(N__15865),
            .in3(N__16443),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_1_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_1_25_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI82223_3_LC_1_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11542),
            .in3(N__14064),
            .lcout(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_1_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_1_25_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_1_25_3  (
            .in0(N__18460),
            .in1(N__23601),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_1_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_1_25_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_1_25_4  (
            .in0(N__20686),
            .in1(_gnd_net_),
            .in2(N__23702),
            .in3(N__18462),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_3_LC_1_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_1_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_1_25_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_1_25_5  (
            .in0(N__12385),
            .in1(N__12364),
            .in2(N__24967),
            .in3(N__18630),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29306),
            .ce(),
            .sr(N__28786));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_1_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_1_26_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_1_26_0  (
            .in0(N__16149),
            .in1(N__23653),
            .in2(_gnd_net_),
            .in3(N__20702),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_1_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_1_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_1_26_1  (
            .in0(_gnd_net_),
            .in1(N__17842),
            .in2(_gnd_net_),
            .in3(N__12867),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_1_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_1_26_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_1_26_2  (
            .in0(_gnd_net_),
            .in1(N__16313),
            .in2(N__11611),
            .in3(N__12789),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_1_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_1_26_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_1_26_3  (
            .in0(N__23652),
            .in1(_gnd_net_),
            .in2(N__11608),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_1_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_1_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_1_26_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_1_26_4  (
            .in0(N__23849),
            .in1(N__13113),
            .in2(_gnd_net_),
            .in3(N__23654),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_1_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_1_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_1_26_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_1_26_5  (
            .in0(N__23655),
            .in1(N__28962),
            .in2(N__11605),
            .in3(N__17843),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29297),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_1_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_1_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_1_26_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_1_26_6  (
            .in0(N__28961),
            .in1(N__11604),
            .in2(N__12829),
            .in3(N__23657),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29297),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_1_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_1_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_1_26_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_1_26_7  (
            .in0(N__23656),
            .in1(N__26697),
            .in2(N__20593),
            .in3(N__12868),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29297),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_1_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_1_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_1_27_0 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_1_27_0  (
            .in0(N__20554),
            .in1(N__18676),
            .in2(N__20381),
            .in3(N__12774),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_4_LC_1_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_1_27_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_1_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_1_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24481),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29288),
            .ce(N__25065),
            .sr(N__28792));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_1_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_1_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_1_27_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_1_27_3  (
            .in0(N__18675),
            .in1(N__23763),
            .in2(_gnd_net_),
            .in3(N__20689),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_1_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_1_27_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_1_27_4  (
            .in0(N__20690),
            .in1(_gnd_net_),
            .in2(N__23810),
            .in3(N__20439),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_1_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_1_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_1_27_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_1_27_5  (
            .in0(N__20438),
            .in1(N__23767),
            .in2(_gnd_net_),
            .in3(N__20691),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_1_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_1_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_1_27_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_1_27_6  (
            .in0(N__20692),
            .in1(_gnd_net_),
            .in2(N__23811),
            .in3(N__16194),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_1_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_1_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_1_27_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_1_27_7  (
            .in0(N__16195),
            .in1(N__23771),
            .in2(_gnd_net_),
            .in3(N__20693),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_1_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_1_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_1_28_0  (
            .in0(_gnd_net_),
            .in1(N__13012),
            .in2(N__11662),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_28_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_1_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_1_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_1_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_1_28_1  (
            .in0(_gnd_net_),
            .in1(N__16225),
            .in2(_gnd_net_),
            .in3(N__11650),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_1_28_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_1_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_1_28_2  (
            .in0(_gnd_net_),
            .in1(N__13081),
            .in2(N__12940),
            .in3(N__11647),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_1_28_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_1_28_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_1_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11644),
            .in3(N__11623),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_1_28_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_1_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_1_28_4  (
            .in0(_gnd_net_),
            .in1(N__11620),
            .in2(_gnd_net_),
            .in3(N__11614),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_1_28_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_1_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_1_28_5  (
            .in0(_gnd_net_),
            .in1(N__17731),
            .in2(_gnd_net_),
            .in3(N__11725),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_1_28_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_1_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_1_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_1_28_6  (
            .in0(_gnd_net_),
            .in1(N__12880),
            .in2(N__12952),
            .in3(N__11722),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_1_28_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_1_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_1_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_1_28_7  (
            .in0(_gnd_net_),
            .in1(N__11719),
            .in2(_gnd_net_),
            .in3(N__11713),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_1_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_1_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_1_29_0  (
            .in0(_gnd_net_),
            .in1(N__13048),
            .in2(_gnd_net_),
            .in3(N__11710),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_1_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_1_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_1_29_1  (
            .in0(_gnd_net_),
            .in1(N__13228),
            .in2(_gnd_net_),
            .in3(N__11707),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_1_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_1_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_1_29_2  (
            .in0(_gnd_net_),
            .in1(N__11704),
            .in2(_gnd_net_),
            .in3(N__11695),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_1_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_1_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_1_29_3  (
            .in0(_gnd_net_),
            .in1(N__11692),
            .in2(_gnd_net_),
            .in3(N__11683),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_1_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_1_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_1_29_4  (
            .in0(_gnd_net_),
            .in1(N__11680),
            .in2(_gnd_net_),
            .in3(N__11668),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_1_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_1_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_1_29_5  (
            .in0(_gnd_net_),
            .in1(N__13141),
            .in2(N__12961),
            .in3(N__11665),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_1_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_1_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_1_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_1_29_6  (
            .in0(_gnd_net_),
            .in1(N__18277),
            .in2(_gnd_net_),
            .in3(N__11839),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_1_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_1_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_1_29_7  (
            .in0(_gnd_net_),
            .in1(N__16471),
            .in2(_gnd_net_),
            .in3(N__11836),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_1_30_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_1_30_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18265),
            .in3(N__11833),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_1_30_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_1_30_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_1_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13066),
            .in3(N__11830),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_1_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_1_30_2 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_1_30_2  (
            .in0(N__23780),
            .in1(N__17565),
            .in2(N__20807),
            .in3(N__11827),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_0_LC_2_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_0_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_0_LC_2_10_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Commands_frame_decoder.source_offset1data_0_LC_2_10_1  (
            .in0(N__28941),
            .in1(N__11820),
            .in2(N__16676),
            .in3(N__29846),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_2_LC_2_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_2_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_2_LC_2_10_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \Commands_frame_decoder.source_offset1data_2_LC_2_10_2  (
            .in0(N__28355),
            .in1(N__16672),
            .in2(N__11805),
            .in3(N__28944),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_1_LC_2_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_1_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_1_LC_2_10_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Commands_frame_decoder.source_offset1data_1_LC_2_10_5  (
            .in0(N__28942),
            .in1(N__11781),
            .in2(N__16677),
            .in3(N__27767),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_p_en_LC_2_10_6 .C_ON=1'b0;
    defparam \pid_alt.source_p_en_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_p_en_LC_2_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.source_p_en_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__13836),
            .in2(_gnd_net_),
            .in3(N__28940),
            .lcout(\pid_alt.source_p_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_3_LC_2_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_3_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_3_LC_2_10_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Commands_frame_decoder.source_offset1data_3_LC_2_10_7  (
            .in0(N__28943),
            .in1(N__12033),
            .in2(N__16678),
            .in3(N__28113),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_5_LC_2_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_5_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_5_LC_2_11_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \Commands_frame_decoder.source_offset1data_5_LC_2_11_1  (
            .in0(N__28230),
            .in1(N__16665),
            .in2(N__12019),
            .in3(N__28978),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29382),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_2_12_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_2_12_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_2_12_5  (
            .in0(N__13147),
            .in1(N__13680),
            .in2(N__13258),
            .in3(N__13351),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29379),
            .ce(),
            .sr(N__28720));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_2_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_2_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__13464),
            .in2(_gnd_net_),
            .in3(N__28932),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_2_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_2_13_0 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_2_13_0  (
            .in0(N__12151),
            .in1(N__12144),
            .in2(N__12124),
            .in3(N__13468),
            .lcout(\dron_frame_decoder_1.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_2_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_2_13_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_2_13_1  (
            .in0(N__11906),
            .in1(N__11864),
            .in2(_gnd_net_),
            .in3(N__11970),
            .lcout(\dron_frame_decoder_1.WDT10lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_2_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_2_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_2_13_2  (
            .in0(N__11958),
            .in1(N__11946),
            .in2(N__11935),
            .in3(N__11919),
            .lcout(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_2_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_2_13_3 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_2_13_3  (
            .in0(N__11907),
            .in1(N__11892),
            .in2(N__11881),
            .in3(N__11865),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_2_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_2_13_4 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_2_13_4  (
            .in0(N__11850),
            .in1(N__12166),
            .in2(N__12160),
            .in3(N__12157),
            .lcout(\dron_frame_decoder_1.WDT10lt14_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_2_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_2_13_5 .LUT_INIT=16'b0011001100111111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__12143),
            .in2(N__12127),
            .in3(N__12119),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_14_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_14_0  (
            .in0(N__12197),
            .in1(N__15011),
            .in2(N__14848),
            .in3(N__15088),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__13721),
            .sr(N__28730));
    defparam \pid_alt.error_cry_0_c_inv_LC_2_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_2_14_1  (
            .in0(N__12073),
            .in1(N__27273),
            .in2(_gnd_net_),
            .in3(N__12084),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_2_14_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_2_14_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_2_14_2  (
            .in0(N__12198),
            .in1(N__15087),
            .in2(N__15199),
            .in3(N__15013),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__13721),
            .sr(N__28730));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_2_14_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_2_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12061),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_2_14_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_2_14_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_2_14_4  (
            .in0(N__12199),
            .in1(N__15012),
            .in2(N__15136),
            .in3(N__15089),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__13721),
            .sr(N__28730));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_14_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12049),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_2_14_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_2_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15090),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__13721),
            .sr(N__28730));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12241),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_2_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_2_15_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_2_15_0  (
            .in0(N__12195),
            .in1(N__15006),
            .in2(N__14815),
            .in3(N__15084),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29369),
            .ce(N__13726),
            .sr(N__28734));
    defparam \pid_alt.error_axb_1_LC_2_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_2_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12229),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude8lto3_0_LC_2_15_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude8lto3_0_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude8lto3_0_LC_2_15_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude8lto3_0_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__15254),
            .in2(_gnd_net_),
            .in3(N__15287),
            .lcout(),
            .ltout(\dron_frame_decoder_1.source_Altitude8lto3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude8lto5_LC_2_15_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude8lto5_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude8lto5_LC_2_15_3 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude8lto5_LC_2_15_3  (
            .in0(N__15125),
            .in1(N__14810),
            .in2(N__12217),
            .in3(N__15191),
            .lcout(\dron_frame_decoder_1.source_Altitude8lt7_0 ),
            .ltout(\dron_frame_decoder_1.source_Altitude8lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_2_15_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_2_15_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_2_15_4  (
            .in0(N__15086),
            .in1(N__15007),
            .in2(N__12214),
            .in3(N__15288),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29369),
            .ce(N__13726),
            .sr(N__28734));
    defparam \pid_alt.error_axb_2_LC_2_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_2_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12211),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_2_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_2_15_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_2_15_6  (
            .in0(N__12196),
            .in1(N__15255),
            .in2(N__15016),
            .in3(N__15085),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29369),
            .ce(N__13726),
            .sr(N__28734));
    defparam \pid_alt.error_axb_3_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_2_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12178),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_2_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_2_16_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_2_16_0  (
            .in0(N__12289),
            .in1(N__16894),
            .in2(N__12343),
            .in3(N__28098),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29364),
            .ce(),
            .sr(N__28739));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_2_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_2_16_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_2_16_2  (
            .in0(N__12287),
            .in1(N__16892),
            .in2(N__27769),
            .in3(N__12324),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29364),
            .ce(),
            .sr(N__28739));
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_2_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_2_16_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_1_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__27812),
            .in2(_gnd_net_),
            .in3(N__27622),
            .lcout(\Commands_frame_decoder.source_CH1data8lto7Z0Z_1 ),
            .ltout(\Commands_frame_decoder.source_CH1data8lto7Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_2_16_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_2_16_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_2_16_4  (
            .in0(N__12259),
            .in1(N__28220),
            .in2(N__12310),
            .in3(N__27977),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_2_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_2_16_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_2_16_5  (
            .in0(N__16891),
            .in1(N__29845),
            .in2(N__12307),
            .in3(N__12303),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29364),
            .ce(),
            .sr(N__28739));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_2_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_2_16_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_2_16_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_2_16_6  (
            .in0(N__12288),
            .in1(N__16893),
            .in2(N__28362),
            .in3(N__12273),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29364),
            .ce(),
            .sr(N__28739));
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_2_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_2_17_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto3_LC_2_17_0  (
            .in0(N__28064),
            .in1(N__28308),
            .in2(_gnd_net_),
            .in3(N__27718),
            .lcout(\Commands_frame_decoder.source_CH1data8lt7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_2_17_3 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_2_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_2_17_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_4_LC_2_17_3  (
            .in0(N__17036),
            .in1(N__16999),
            .in2(N__17647),
            .in3(N__27825),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29358),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12253),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12397),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_2_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_2_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15091),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29351),
            .ce(N__13573),
            .sr(N__28751));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14814),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29351),
            .ce(N__13573),
            .sr(N__28751));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_2_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_2_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__12999),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_2_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_2_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__12699),
            .in2(N__27207),
            .in3(N__12391),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_2_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_2_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__12900),
            .in2(_gnd_net_),
            .in3(N__12388),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_2_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_2_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__12384),
            .in2(N__27208),
            .in3(N__12352),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_2_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_2_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__12606),
            .in2(_gnd_net_),
            .in3(N__12349),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_2_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_2_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__12567),
            .in2(_gnd_net_),
            .in3(N__12346),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_2_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_2_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__12477),
            .in2(N__27209),
            .in3(N__12451),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_2_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_2_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__12498),
            .in2(_gnd_net_),
            .in3(N__12448),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_2_20_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_2_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__12543),
            .in2(_gnd_net_),
            .in3(N__12445),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_2_20_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_2_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__13791),
            .in2(_gnd_net_),
            .in3(N__12442),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_2_20_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_2_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__12666),
            .in2(_gnd_net_),
            .in3(N__12439),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_2_20_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_2_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__13755),
            .in2(_gnd_net_),
            .in3(N__12436),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_2_20_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_2_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__13944),
            .in2(_gnd_net_),
            .in3(N__12433),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_2_20_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_2_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(N__12639),
            .in2(N__27206),
            .in3(N__12430),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_2_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_2_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(N__12427),
            .in2(_gnd_net_),
            .in3(N__12412),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29340),
            .ce(N__25066),
            .sr(N__28764));
    defparam \ppm_encoder_1.throttle_1_LC_2_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_2_21_1 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_2_21_1  (
            .in0(N__24842),
            .in1(N__12703),
            .in2(N__14466),
            .in3(N__12679),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29333),
            .ce(),
            .sr(N__28770));
    defparam \ppm_encoder_1.throttle_10_LC_2_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_2_21_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_2_21_4  (
            .in0(N__12670),
            .in1(N__12646),
            .in2(N__22712),
            .in3(N__24840),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29333),
            .ce(),
            .sr(N__28770));
    defparam \ppm_encoder_1.throttle_13_LC_2_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_2_21_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_2_21_5 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_2_21_5  (
            .in0(N__24841),
            .in1(N__12640),
            .in2(N__20129),
            .in3(N__12616),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29333),
            .ce(),
            .sr(N__28770));
    defparam \ppm_encoder_1.throttle_4_LC_2_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_2_21_7 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_2_21_7  (
            .in0(N__24843),
            .in1(N__12610),
            .in2(N__13994),
            .in3(N__12589),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29333),
            .ce(),
            .sr(N__28770));
    defparam \ppm_encoder_1.throttle_5_LC_2_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_2_22_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_2_22_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_2_22_0  (
            .in0(N__12580),
            .in1(N__12571),
            .in2(N__24911),
            .in3(N__18605),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29326),
            .ce(),
            .sr(N__28774));
    defparam \ppm_encoder_1.throttle_8_LC_2_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_2_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_2_22_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_2_22_1  (
            .in0(N__12547),
            .in1(N__12520),
            .in2(N__13870),
            .in3(N__24853),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29326),
            .ce(),
            .sr(N__28774));
    defparam \ppm_encoder_1.throttle_7_LC_2_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_2_22_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_2_22_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_2_22_2  (
            .in0(N__12511),
            .in1(N__12502),
            .in2(N__24912),
            .in3(N__12744),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29326),
            .ce(),
            .sr(N__28774));
    defparam \ppm_encoder_1.elevator_7_LC_2_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_2_22_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_2_22_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_2_22_4  (
            .in0(N__24589),
            .in1(N__25966),
            .in2(N__24910),
            .in3(N__12724),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29326),
            .ce(),
            .sr(N__28774));
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0  (
            .in0(N__20408),
            .in1(N__15746),
            .in2(N__12748),
            .in3(N__15848),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__14335),
            .in2(N__12757),
            .in3(N__12754),
            .lcout(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2  (
            .in0(N__12722),
            .in1(N__20150),
            .in2(N__16055),
            .in3(N__15970),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3  (
            .in0(N__12743),
            .in1(N__22763),
            .in2(_gnd_net_),
            .in3(N__12723),
            .lcout(\ppm_encoder_1.N_298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_2_23_5  (
            .in0(N__20151),
            .in1(N__22495),
            .in2(N__24908),
            .in3(N__24130),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29315),
            .ce(),
            .sr(N__28776));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_2_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_2_24_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_2_24_0  (
            .in0(N__12850),
            .in1(N__12807),
            .in2(N__16319),
            .in3(N__23552),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_2_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_2_24_1 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_2_24_1  (
            .in0(N__23556),
            .in1(N__12790),
            .in2(N__12709),
            .in3(N__15977),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_2_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_2_24_2 .LUT_INIT=16'b1010111100001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIALN65_1_LC_2_24_2  (
            .in0(N__14462),
            .in1(N__16264),
            .in2(N__12706),
            .in3(N__15847),
            .lcout(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_2_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_2_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_2_24_3  (
            .in0(N__18538),
            .in1(N__17809),
            .in2(N__23629),
            .in3(N__16311),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_2_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_2_24_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__17941),
            .in2(_gnd_net_),
            .in3(N__18902),
            .lcout(\ppm_encoder_1.PPM_STATE_58_d ),
            .ltout(\ppm_encoder_1.PPM_STATE_58_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_2_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_2_24_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_2_24_5  (
            .in0(N__18537),
            .in1(N__17808),
            .in2(N__12871),
            .in3(N__16312),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_2_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_2_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_2_24_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_2_24_6  (
            .in0(N__18694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18904),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29307),
            .ce(),
            .sr(N__28780));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_2_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_2_24_7 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_2_24_7  (
            .in0(N__18903),
            .in1(N__18693),
            .in2(N__17951),
            .in3(N__18976),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29307),
            .ce(),
            .sr(N__28780));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_2_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_2_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__20666),
            .in2(_gnd_net_),
            .in3(N__23557),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_2_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_2_25_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(N__12821),
            .in2(_gnd_net_),
            .in3(N__12865),
            .lcout(\ppm_encoder_1.N_226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_2_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_2_25_2 .LUT_INIT=16'b1111001011110110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_2_25_2  (
            .in0(N__12808),
            .in1(N__23560),
            .in2(N__28980),
            .in3(N__20667),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29298),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_2_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_2_25_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_2_25_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_2_25_3  (
            .in0(N__23559),
            .in1(N__20958),
            .in2(N__12849),
            .in3(N__28972),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29298),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_2_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_2_25_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_2_25_4  (
            .in0(N__12866),
            .in1(N__12842),
            .in2(N__12828),
            .in3(N__12806),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_2_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_2_25_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_2_25_5  (
            .in0(N__23558),
            .in1(_gnd_net_),
            .in2(N__12778),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_2_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_2_25_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_2_25_6  (
            .in0(N__13995),
            .in1(N__12775),
            .in2(N__12760),
            .in3(N__15846),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_2_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_2_25_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_2_25_7  (
            .in0(N__14002),
            .in1(N__18655),
            .in2(N__12943),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_2_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_2_26_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_2_26_0  (
            .in0(N__23651),
            .in1(N__15902),
            .in2(N__13135),
            .in3(N__16440),
            .lcout(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_2_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_2_26_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_2_26_1 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_2_26_1  (
            .in0(N__18227),
            .in1(N__12928),
            .in2(N__18026),
            .in3(N__14077),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29289),
            .ce(),
            .sr(N__28787));
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_2_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_2_26_2 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ppm_encoder_1.throttle_RNIR7352_2_LC_2_26_2  (
            .in0(N__14378),
            .in1(N__15864),
            .in2(N__15909),
            .in3(N__16441),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_2_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_2_26_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5V123_2_LC_2_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12919),
            .in3(N__14097),
            .lcout(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_2_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_2_26_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIANUS_2_LC_2_26_4  (
            .in0(N__23650),
            .in1(N__20687),
            .in2(_gnd_net_),
            .in3(N__15901),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_2_LC_2_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_2_26_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_2_26_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_2_26_5  (
            .in0(N__12916),
            .in1(N__12907),
            .in2(N__24966),
            .in3(N__14379),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29289),
            .ce(),
            .sr(N__28787));
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_2_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_2_26_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_2_26_7  (
            .in0(N__16442),
            .in1(N__13133),
            .in2(N__23798),
            .in3(N__21102),
            .lcout(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_2_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_2_27_0 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_2_27_0  (
            .in0(N__13114),
            .in1(N__23761),
            .in2(N__12979),
            .in3(N__16448),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_2_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_2_27_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_2_27_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_2_27_1  (
            .in0(N__13018),
            .in1(N__18010),
            .in2(N__13024),
            .in3(N__18243),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29283),
            .ce(),
            .sr(N__28789));
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_2_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_2_27_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_2_27_2  (
            .in0(N__12973),
            .in1(N__23760),
            .in2(_gnd_net_),
            .in3(N__20688),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_2_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_2_27_3 .LUT_INIT=16'b0011110000001111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_2_27_3  (
            .in0(_gnd_net_),
            .in1(N__18485),
            .in2(N__13021),
            .in3(N__15863),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_4  (
            .in0(N__12974),
            .in1(N__23762),
            .in2(N__13129),
            .in3(N__16447),
            .lcout(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_2_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_2_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_2_27_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIN3352_0_LC_2_27_5  (
            .in0(N__14127),
            .in1(N__18484),
            .in2(_gnd_net_),
            .in3(N__15862),
            .lcout(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_0_LC_2_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_2_27_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_2_27_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_2_27_6  (
            .in0(N__18486),
            .in1(N__24907),
            .in2(_gnd_net_),
            .in3(N__13006),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29283),
            .ce(),
            .sr(N__28789));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_2_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_2_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_2_27_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_2_27_7  (
            .in0(N__20361),
            .in1(N__20555),
            .in2(_gnd_net_),
            .in3(N__12975),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_2_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_2_28_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_2_28_0  (
            .in0(N__13128),
            .in1(N__21043),
            .in2(N__23809),
            .in3(N__16457),
            .lcout(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_2_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_2_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_2_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_2_28_1  (
            .in0(_gnd_net_),
            .in1(N__13124),
            .in2(_gnd_net_),
            .in3(N__23754),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_2_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_2_28_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_2_28_2  (
            .in0(N__23755),
            .in1(_gnd_net_),
            .in2(N__13134),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_2_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_2_28_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_2_28_3  (
            .in0(_gnd_net_),
            .in1(N__23753),
            .in2(_gnd_net_),
            .in3(N__13123),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_17_LC_2_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_2_28_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_2_28_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_2_28_6  (
            .in0(N__18063),
            .in1(N__18244),
            .in2(N__14401),
            .in3(N__13075),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29277),
            .ce(),
            .sr(N__28793));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_28_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_28_7  (
            .in0(N__22914),
            .in1(N__23756),
            .in2(_gnd_net_),
            .in3(N__20759),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_2_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_2_29_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_2_29_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_2_29_0  (
            .in0(N__18248),
            .in1(N__13054),
            .in2(N__18112),
            .in3(N__14266),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29270),
            .ce(),
            .sr(N__28796));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_2_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_2_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_2_29_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_2_29_1  (
            .in0(N__13040),
            .in1(_gnd_net_),
            .in2(N__23812),
            .in3(N__20792),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_2_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_2_29_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_2_29_2  (
            .in0(N__20790),
            .in1(N__23772),
            .in2(_gnd_net_),
            .in3(N__13041),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_2_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_2_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_2_29_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_2_29_3  (
            .in0(N__13042),
            .in1(N__20570),
            .in2(N__20382),
            .in3(N__19834),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_2_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_2_29_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_2_29_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_2_29_4  (
            .in0(N__18249),
            .in1(N__13030),
            .in2(N__18113),
            .in3(N__14221),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29270),
            .ce(),
            .sr(N__28796));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_2_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_2_29_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_2_29_5  (
            .in0(N__13220),
            .in1(_gnd_net_),
            .in2(N__23813),
            .in3(N__20793),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_2_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_2_29_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_2_29_6  (
            .in0(N__20791),
            .in1(N__23773),
            .in2(_gnd_net_),
            .in3(N__13221),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_2_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_2_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_2_29_7 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_2_29_7  (
            .in0(N__13222),
            .in1(N__20571),
            .in2(N__20383),
            .in3(N__19756),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_2_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_2_30_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_2_30_1  (
            .in0(N__20957),
            .in1(N__13210),
            .in2(_gnd_net_),
            .in3(N__15490),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_6_LC_3_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_6_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_6_LC_3_10_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \Commands_frame_decoder.source_offset1data_6_LC_3_10_1  (
            .in0(N__16664),
            .in1(N__27632),
            .in2(N__13194),
            .in3(N__28977),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29383),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset1data_1_4_LC_3_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_1_4_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset1data_1_4_LC_3_10_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \Commands_frame_decoder.source_offset1data_1_4_LC_3_10_3  (
            .in0(N__16663),
            .in1(N__27869),
            .in2(N__13173),
            .in3(N__28976),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29383),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_3_12_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_3_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_3_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__15252),
            .in2(_gnd_net_),
            .in3(N__15189),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_a3_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_12_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_3_12_3  (
            .in0(N__15083),
            .in1(N__13253),
            .in2(N__13153),
            .in3(N__14809),
            .lcout(\dron_frame_decoder_1.state_ns_0_a3_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_1_LC_3_12_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_1_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_1_LC_3_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_1_LC_3_12_4  (
            .in0(N__14808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15082),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_a3_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_1_LC_3_12_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_1_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_1_LC_3_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_1_LC_3_12_5  (
            .in0(N__15190),
            .in1(N__15253),
            .in2(N__13150),
            .in3(N__13387),
            .lcout(\dron_frame_decoder_1.state_ns_0_a3_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_5_LC_3_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_3_13_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_3_13_0  (
            .in0(N__13683),
            .in1(N__13270),
            .in2(N__13483),
            .in3(N__13597),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(N__28721));
    defparam \dron_frame_decoder_1.state_6_LC_3_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_3_13_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_3_13_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_3_13_2  (
            .in0(N__13684),
            .in1(N__13619),
            .in2(N__13484),
            .in3(N__13525),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(N__28721));
    defparam \dron_frame_decoder_1.state_3_LC_3_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_3_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_3_13_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_3_13_3  (
            .in0(N__13291),
            .in1(N__13682),
            .in2(N__13285),
            .in3(N__13347),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(N__28721));
    defparam \dron_frame_decoder_1.state_7_LC_3_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_3_13_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_3_13_6  (
            .in0(N__13685),
            .in1(N__13620),
            .in2(N__13485),
            .in3(N__13651),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(N__28721));
    defparam \dron_frame_decoder_1.state_2_LC_3_13_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_3_13_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_3_13_7  (
            .in0(N__13269),
            .in1(N__13681),
            .in2(N__13284),
            .in3(N__13478),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(N__28721));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_3_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_3_14_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_3_14_0  (
            .in0(N__13360),
            .in1(N__13393),
            .in2(N__14872),
            .in3(N__13340),
            .lcout(),
            .ltout(\dron_frame_decoder_1.N_217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_0_LC_3_14_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_3_14_1 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_3_14_1 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_3_14_1  (
            .in0(N__13386),
            .in1(N__13234),
            .in2(N__13261),
            .in3(N__13689),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29370),
            .ce(),
            .sr(N__28725));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_3_14_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_3_14_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_3_14_6  (
            .in0(N__13521),
            .in1(N__13385),
            .in2(N__13482),
            .in3(N__13257),
            .lcout(\dron_frame_decoder_1.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_5_0_LC_3_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_5_0_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_5_0_LC_3_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_5_0_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__15049),
            .in2(_gnd_net_),
            .in3(N__15165),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_i_a2_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_3_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_3_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_3_15_1  (
            .in0(N__14793),
            .in1(N__13380),
            .in2(N__13396),
            .in3(N__15234),
            .lcout(\dron_frame_decoder_1.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_1_2_LC_3_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_1_2_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_1_2_LC_3_15_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_1_2_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__27621),
            .in2(_gnd_net_),
            .in3(N__29831),
            .lcout(\Commands_frame_decoder.state_1_ns_0_a4_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_3_15_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_3_15_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \dron_frame_decoder_1.state_RNO_3_0_LC_3_15_3  (
            .in0(N__13526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13381),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_5  (
            .in0(N__13460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14971),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_LC_3_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_LC_3_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_2_0_LC_3_15_6  (
            .in0(N__15107),
            .in1(N__14831),
            .in2(N__13354),
            .in3(N__15283),
            .lcout(\dron_frame_decoder_1.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_1_0_LC_3_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_1_0_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_1_0_LC_3_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_ns_i_a2_3_1_0_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__27957),
            .in2(_gnd_net_),
            .in3(N__27714),
            .lcout(\Commands_frame_decoder.state_1_ns_i_a2_3_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_3_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_3_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_3_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27956),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29359),
            .ce(N__16918),
            .sr(N__28735));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_3_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_3_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27826),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29359),
            .ce(N__16918),
            .sr(N__28735));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_3_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_3_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28168),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29359),
            .ce(N__16918),
            .sr(N__28735));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_3_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_3_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27623),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29359),
            .ce(N__16918),
            .sr(N__28735));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_3_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_3_17_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_5_LC_3_17_0  (
            .in0(N__13534),
            .in1(N__13630),
            .in2(N__13603),
            .in3(N__28933),
            .lcout(\dron_frame_decoder_1.N_238_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_4_LC_3_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_3_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_3_17_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_3_17_1  (
            .in0(N__13424),
            .in1(N__13602),
            .in2(N__13650),
            .in3(N__13693),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29352),
            .ce(),
            .sr(N__28740));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_3_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_3_17_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__13643),
            .in2(_gnd_net_),
            .in3(N__13423),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_0_0 ),
            .ltout(\dron_frame_decoder_1.un1_sink_data_valid_5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_3_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_3_17_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_3_17_3  (
            .in0(N__13624),
            .in1(N__13598),
            .in2(N__13579),
            .in3(N__13533),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_3_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_3_17_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13576),
            .in3(N__26687),
            .lcout(\dron_frame_decoder_1.N_230_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_LC_3_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_3_18_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_3_18_0  (
            .in0(N__13828),
            .in1(N__13532),
            .in2(_gnd_net_),
            .in3(N__13441),
            .lcout(drone_frame_decoder_data_rdy_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29346),
            .ce(),
            .sr(N__28745));
    defparam \uart_pc.bit_Count_0_LC_3_18_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_3_18_3 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \uart_pc.bit_Count_0_LC_3_18_3  (
            .in0(N__19370),
            .in1(N__19486),
            .in2(N__17283),
            .in3(N__19558),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29346),
            .ce(),
            .sr(N__28745));
    defparam \uart_drone.data_rdy_LC_3_18_4 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_3_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.data_rdy_LC_3_18_4  (
            .in0(N__17137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21760),
            .lcout(uart_drone_data_rdy_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29346),
            .ce(),
            .sr(N__28745));
    defparam \pid_alt.source_data_valid_LC_3_18_7 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_LC_3_18_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.source_data_valid_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__13829),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29346),
            .ce(),
            .sr(N__28745));
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_3_19_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_3_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_4_LC_3_19_3  (
            .in0(N__15435),
            .in1(N__15309),
            .in2(N__15421),
            .in3(N__15324),
            .lcout(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_3_19_5 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_3_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_3_19_5  (
            .in0(N__17320),
            .in1(N__17370),
            .in2(_gnd_net_),
            .in3(N__17248),
            .lcout(\uart_pc.N_152 ),
            .ltout(\uart_pc.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_3_19_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_3_19_6 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__19482),
            .in2(N__13810),
            .in3(N__19555),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_3_19_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_3_19_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_3_19_7  (
            .in0(N__17321),
            .in1(N__17371),
            .in2(_gnd_net_),
            .in3(N__17249),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_3_20_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_3_20_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_3_20_1  (
            .in0(N__17281),
            .in1(N__19556),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_3_20_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_3_20_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_3_20_2  (
            .in0(N__13804),
            .in1(N__17386),
            .in2(N__13807),
            .in3(N__17339),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29334),
            .ce(),
            .sr(N__28757));
    defparam \uart_pc.bit_Count_1_LC_3_20_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_3_20_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_1_LC_3_20_3  (
            .in0(N__17282),
            .in1(N__19557),
            .in2(N__17348),
            .in3(N__13803),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29334),
            .ce(),
            .sr(N__28757));
    defparam \ppm_encoder_1.throttle_9_LC_3_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_3_21_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_3_21_3  (
            .in0(N__13795),
            .in1(N__13771),
            .in2(N__24870),
            .in3(N__15456),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29327),
            .ce(),
            .sr(N__28765));
    defparam \ppm_encoder_1.throttle_11_LC_3_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_3_21_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_3_21_5  (
            .in0(N__13765),
            .in1(N__13954),
            .in2(N__24868),
            .in3(N__17918),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29327),
            .ce(),
            .sr(N__28765));
    defparam \ppm_encoder_1.throttle_12_LC_3_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_3_21_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_3_21_7  (
            .in0(N__13948),
            .in1(N__13915),
            .in2(N__24869),
            .in3(N__13900),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29327),
            .ce(),
            .sr(N__28765));
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_3_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_3_22_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNII6JI2_12_LC_3_22_1  (
            .in0(N__20040),
            .in1(N__13898),
            .in2(N__15881),
            .in3(N__15769),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_3_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_3_22_2 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIFQRT5_12_LC_3_22_2  (
            .in0(N__14200),
            .in1(_gnd_net_),
            .in2(N__13909),
            .in3(N__13906),
            .lcout(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_3_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_3_22_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI25DH2_12_LC_3_22_3  (
            .in0(N__22875),
            .in1(N__13880),
            .in2(N__16065),
            .in3(N__15991),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_3_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_3_22_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_3_22_4  (
            .in0(N__13899),
            .in1(N__22876),
            .in2(_gnd_net_),
            .in3(N__22799),
            .lcout(),
            .ltout(\ppm_encoder_1.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_3_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_3_22_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_3_22_5  (
            .in0(N__20938),
            .in1(_gnd_net_),
            .in2(N__13885),
            .in3(N__13881),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_3_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_3_22_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_3_22_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_3_22_6  (
            .in0(N__13882),
            .in1(N__23926),
            .in2(N__24909),
            .in3(N__22420),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29316),
            .ce(),
            .sr(N__28771));
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_3_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_3_23_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.throttle_RNIS5KK2_8_LC_3_23_0  (
            .in0(N__13865),
            .in1(N__15765),
            .in2(N__19830),
            .in3(N__15851),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_3_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_3_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIONI96_8_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(N__14296),
            .in2(N__13849),
            .in3(N__14017),
            .lcout(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_3_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_3_23_2 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNICKVN2_8_LC_3_23_2  (
            .in0(N__19797),
            .in1(N__15479),
            .in2(N__15989),
            .in3(N__16042),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_3_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_3_23_3 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \ppm_encoder_1.throttle_RNIU7KK2_9_LC_3_23_3  (
            .in0(N__15852),
            .in1(N__15457),
            .in2(N__15772),
            .in3(N__19749),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_3_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_3_23_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNITSI96_9_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(N__14251),
            .in2(N__14011),
            .in3(N__14008),
            .lcout(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_3_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_3_23_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_3_23_5  (
            .in0(N__15850),
            .in1(N__20184),
            .in2(N__15771),
            .in3(N__19900),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_3_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_3_23_6 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNIEMVN2_9_LC_3_23_6  (
            .in0(N__19614),
            .in1(N__19875),
            .in2(N__15990),
            .in3(N__16043),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_0  (
            .in0(N__13962),
            .in1(N__14427),
            .in2(N__15988),
            .in3(N__16041),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_4_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24208),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29299),
            .ce(N__25050),
            .sr(N__28777));
    defparam \ppm_encoder_1.elevator_esr_4_LC_3_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_4_LC_3_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_4_LC_3_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_4_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24508),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29299),
            .ce(N__25050),
            .sr(N__28777));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_24_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_3_24_3  (
            .in0(N__13996),
            .in1(N__13963),
            .in2(_gnd_net_),
            .in3(N__18563),
            .lcout(\ppm_encoder_1.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_3_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_3_24_5 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_3_24_5  (
            .in0(N__17715),
            .in1(N__18612),
            .in2(N__15757),
            .in3(N__15849),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_3_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_3_24_6 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_3_24_6  (
            .in0(N__17752),
            .in1(_gnd_net_),
            .in2(N__14149),
            .in3(N__14146),
            .lcout(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_3_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_3_24_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_3_24_7  (
            .in0(N__18582),
            .in1(N__18507),
            .in2(N__16056),
            .in3(N__15969),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_3_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_3_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIVO123_0_LC_3_25_0  (
            .in0(_gnd_net_),
            .in1(N__14140),
            .in2(N__14131),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_3_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_3_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_3_25_1  (
            .in0(_gnd_net_),
            .in1(N__16260),
            .in2(N__14113),
            .in3(N__14104),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_3_25_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_3_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_3_25_2  (
            .in0(_gnd_net_),
            .in1(N__14101),
            .in2(N__14086),
            .in3(N__14071),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_3_25_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_3_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_3_25_3  (
            .in0(_gnd_net_),
            .in1(N__14068),
            .in2(N__14053),
            .in3(N__14032),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_3_25_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_3_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_3_25_4  (
            .in0(_gnd_net_),
            .in1(N__18654),
            .in2(N__14029),
            .in3(N__14020),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_3_25_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_3_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_3_25_5  (
            .in0(_gnd_net_),
            .in1(N__17745),
            .in2(N__14365),
            .in3(N__14356),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_3_25_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_3_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_3_25_6  (
            .in0(_gnd_net_),
            .in1(N__18357),
            .in2(N__14353),
            .in3(N__14338),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_3_25_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_3_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(N__14334),
            .in2(N__14311),
            .in3(N__14299),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_3_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_3_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__14292),
            .in2(N__14278),
            .in3(N__14254),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_3_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_3_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__14247),
            .in2(N__14233),
            .in3(N__14209),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_3_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_3_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__15687),
            .in2(N__15661),
            .in3(N__14206),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_3_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_3_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__16104),
            .in2(N__16078),
            .in3(N__14203),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_3_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_3_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(N__14199),
            .in2(N__14179),
            .in3(N__14167),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_3_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_3_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_3_26_5  (
            .in0(_gnd_net_),
            .in1(N__16344),
            .in2(N__14164),
            .in3(N__14413),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_3_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_3_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_3_26_6  (
            .in0(_gnd_net_),
            .in1(N__18294),
            .in2(N__15616),
            .in3(N__14410),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_3_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_3_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_3_26_7  (
            .in0(_gnd_net_),
            .in1(N__16504),
            .in2(N__16381),
            .in3(N__14407),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_3_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_3_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_3_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__14524),
            .in2(_gnd_net_),
            .in3(N__14404),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_3_27_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_3_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_3_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_3_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_3_27_1  (
            .in0(_gnd_net_),
            .in1(N__14386),
            .in2(_gnd_net_),
            .in3(N__14392),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_3_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_3_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_3_27_2  (
            .in0(_gnd_net_),
            .in1(N__16405),
            .in2(_gnd_net_),
            .in3(N__14389),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_3_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_3_27_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_3_27_3  (
            .in0(N__22913),
            .in1(N__23795),
            .in2(_gnd_net_),
            .in3(N__20798),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_27_4 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_27_4  (
            .in0(_gnd_net_),
            .in1(N__22856),
            .in2(N__16333),
            .in3(N__20885),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_3_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_3_27_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_3_27_5 .LUT_INIT=16'b1011101010111110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_3_27_5  (
            .in0(N__28960),
            .in1(N__23796),
            .in2(N__20931),
            .in3(N__20799),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29278),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_3_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_3_27_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_3_27_6  (
            .in0(N__20921),
            .in1(N__22855),
            .in2(_gnd_net_),
            .in3(N__14380),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_3_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_3_27_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_3_27_7  (
            .in0(N__22955),
            .in1(N__23794),
            .in2(_gnd_net_),
            .in3(N__20797),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_3_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_3_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_3_28_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_3_28_2  (
            .in0(N__18231),
            .in1(N__14518),
            .in2(N__18094),
            .in3(N__14506),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29271),
            .ce(),
            .sr(N__28790));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_3_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_3_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_3_29_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_3_29_0  (
            .in0(N__21147),
            .in1(N__14488),
            .in2(N__14476),
            .in3(N__22591),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_3_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_3_29_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_3_29_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_3_29_1  (
            .in0(N__23106),
            .in1(N__14500),
            .in2(_gnd_net_),
            .in3(N__14494),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29267),
            .ce(N__23061),
            .sr(N__28794));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_3_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_3_29_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_3_29_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_3_29_5  (
            .in0(N__23107),
            .in1(N__15643),
            .in2(_gnd_net_),
            .in3(N__14482),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29267),
            .ce(N__23061),
            .sr(N__28794));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_3_30_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_3_30_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_3_30_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_3_30_4  (
            .in0(N__20932),
            .in1(N__22857),
            .in2(_gnd_net_),
            .in3(N__14467),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_30_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_30_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_30_5  (
            .in0(N__20933),
            .in1(N__14440),
            .in2(_gnd_net_),
            .in3(N__14431),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_4_10_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__14559),
            .in2(_gnd_net_),
            .in3(N__14580),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_4_10_5 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_4_10_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_4_10_5  (
            .in0(N__16782),
            .in1(N__16702),
            .in2(N__14416),
            .in3(N__16597),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_4_11_2 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_4_11_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \reset_module_System.count_2_LC_4_11_2  (
            .in0(N__16701),
            .in1(N__14536),
            .in2(N__16783),
            .in3(N__16596),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29376),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_4_11_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_4_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_4_11_3  (
            .in0(N__14685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14576),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_4_11_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_4_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_4_11_4  (
            .in0(N__14637),
            .in1(N__14652),
            .in2(N__14623),
            .in3(N__14670),
            .lcout(),
            .ltout(\reset_module_System.reset6_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_4_11_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_4_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_4_11_5  (
            .in0(N__14710),
            .in1(N__14731),
            .in2(N__14596),
            .in3(N__14593),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_4_11_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_4_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_4_11_6  (
            .in0(N__14758),
            .in1(N__14557),
            .in2(N__14587),
            .in3(N__14881),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_4_11_7 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_4_11_7 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_4_11_7  (
            .in0(N__14558),
            .in1(N__16777),
            .in2(N__14584),
            .in3(N__16700),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29376),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_4_12_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__14581),
            .in2(N__14560),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_4_12_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_4_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__16794),
            .in2(_gnd_net_),
            .in3(N__14530),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_4_12_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_4_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__16824),
            .in2(_gnd_net_),
            .in3(N__14527),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_4_12_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_4_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__14686),
            .in2(_gnd_net_),
            .in3(N__14674),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_4_12_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_4_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__14671),
            .in2(_gnd_net_),
            .in3(N__14659),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_4_12_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_4_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__16836),
            .in2(_gnd_net_),
            .in3(N__14656),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_4_12_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_4_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__14653),
            .in2(_gnd_net_),
            .in3(N__14641),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_4_12_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_4_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__14638),
            .in2(_gnd_net_),
            .in3(N__14626),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__29374),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_4_13_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_4_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__14619),
            .in2(_gnd_net_),
            .in3(N__14605),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_4_13_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_4_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__16740),
            .in2(_gnd_net_),
            .in3(N__14602),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_4_13_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_4_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__16713),
            .in2(_gnd_net_),
            .in3(N__14599),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_4_13_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_4_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__14754),
            .in2(_gnd_net_),
            .in3(N__14743),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_4_13_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_4_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__14893),
            .in2(_gnd_net_),
            .in3(N__14740),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_4_13_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_4_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__16752),
            .in2(_gnd_net_),
            .in3(N__14737),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_4_13_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_4_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__14917),
            .in2(_gnd_net_),
            .in3(N__14734),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_4_13_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_4_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__14730),
            .in2(_gnd_net_),
            .in3(N__14716),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_4_14_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_4_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__16725),
            .in2(_gnd_net_),
            .in3(N__14713),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__29365),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_4_14_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_4_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__14709),
            .in2(_gnd_net_),
            .in3(N__14695),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__29365),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_4_14_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_4_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__14926),
            .in2(_gnd_net_),
            .in3(N__14692),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__29365),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_4_14_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_4_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__16809),
            .in2(_gnd_net_),
            .in3(N__14689),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__29365),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_4_14_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_4_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__14904),
            .in2(_gnd_net_),
            .in3(N__14929),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29365),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_4_14_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_4_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_4_14_7  (
            .in0(N__14925),
            .in1(N__14916),
            .in2(N__14905),
            .in3(N__14892),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_4_0_LC_4_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_4_0_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_4_0_LC_4_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_RNO_4_0_LC_4_15_0  (
            .in0(N__15233),
            .in1(N__15050),
            .in2(N__14799),
            .in3(N__15169),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_4_15_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_4_15_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_4_15_1  (
            .in0(N__21756),
            .in1(N__17135),
            .in2(_gnd_net_),
            .in3(N__26647),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_4_15_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_4_15_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_4_15_2  (
            .in0(N__17136),
            .in1(_gnd_net_),
            .in2(N__14860),
            .in3(_gnd_net_),
            .lcout(\uart_drone.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_4_15_4 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_4_15_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \uart_pc.data_5_LC_4_15_4  (
            .in0(N__28203),
            .in1(N__17037),
            .in2(N__17593),
            .in3(N__16987),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29360),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_0_2_LC_4_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_0_2_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_0_2_LC_4_15_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_0_2_LC_4_15_7  (
            .in0(N__28312),
            .in1(N__27857),
            .in2(N__14857),
            .in3(N__24361),
            .lcout(\Commands_frame_decoder.state_1_ns_0_a4_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_0_LC_4_16_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_4_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21505),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_1_LC_4_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_4_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21487),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_2_LC_4_16_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_4_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21841),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_3_LC_4_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_4_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone.data_esr_3_LC_4_16_3  (
            .in0(N__21814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_4_LC_4_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_4_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21655),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_5_LC_4_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_4_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17088),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_6_LC_4_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17073),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_drone.data_esr_7_LC_4_16_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_4_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17058),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29353),
            .ce(N__14950),
            .sr(N__14944));
    defparam \uart_pc.data_3_LC_4_17_0 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_4_17_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \uart_pc.data_3_LC_4_17_0  (
            .in0(N__16993),
            .in1(N__28063),
            .in2(N__17698),
            .in3(N__17024),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29347),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_17_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_17_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_17_2  (
            .in0(N__26646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19327),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_4_17_3 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_4_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_4_17_3 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \uart_pc.data_1_LC_4_17_3  (
            .in0(N__17188),
            .in1(N__16992),
            .in2(N__14932),
            .in3(N__27713),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29347),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_4_17_5 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_4_17_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \uart_pc.data_4_LC_4_17_5  (
            .in0(N__19328),
            .in1(N__16991),
            .in2(N__27976),
            .in3(N__17671),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29347),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_4_18_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_4_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_4_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__15358),
            .in2(N__17415),
            .in3(N__17416),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_1_LC_4_18_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_4_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_4_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__15352),
            .in2(_gnd_net_),
            .in3(N__15346),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_2_LC_4_18_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_4_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_4_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__15343),
            .in2(_gnd_net_),
            .in3(N__15337),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_3_LC_4_18_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_4_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_4_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__15334),
            .in2(_gnd_net_),
            .in3(N__15328),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_4_LC_4_18_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_4_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_4_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__15325),
            .in2(_gnd_net_),
            .in3(N__15313),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_5_LC_4_18_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_4_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_4_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__15310),
            .in2(_gnd_net_),
            .in3(N__15298),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_6_LC_4_18_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_4_18_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_4_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__15582),
            .in2(_gnd_net_),
            .in3(N__15295),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_7_LC_4_18_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_4_18_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_4_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__15552),
            .in2(_gnd_net_),
            .in3(N__15292),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__29341),
            .ce(),
            .sr(N__17112));
    defparam \Commands_frame_decoder.WDT_8_LC_4_19_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_4_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_4_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__15436),
            .in2(_gnd_net_),
            .in3(N__15424),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_9_LC_4_19_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_4_19_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_4_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__15420),
            .in2(_gnd_net_),
            .in3(N__15406),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_10_LC_4_19_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_4_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_4_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__15370),
            .in2(_gnd_net_),
            .in3(N__15403),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_11_LC_4_19_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_4_19_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_4_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__15598),
            .in2(_gnd_net_),
            .in3(N__15400),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_12_LC_4_19_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_4_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__15568),
            .in2(_gnd_net_),
            .in3(N__15397),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_13_LC_4_19_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_4_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_4_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(N__15384),
            .in2(_gnd_net_),
            .in3(N__15394),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_14_LC_4_19_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_4_19_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_4_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__22337),
            .in2(_gnd_net_),
            .in3(N__15391),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_15_LC_4_19_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_4_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(N__17438),
            .in2(_gnd_net_),
            .in3(N__15388),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29335),
            .ce(),
            .sr(N__17116));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_4_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_4_20_0 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_4_20_0  (
            .in0(N__15566),
            .in1(N__15596),
            .in2(N__15385),
            .in3(N__15369),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_4_20_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_4_20_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_4_20_1  (
            .in0(N__17387),
            .in1(N__17322),
            .in2(_gnd_net_),
            .in3(N__17277),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_4_20_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_4_20_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_4_20_2  (
            .in0(N__17278),
            .in1(_gnd_net_),
            .in2(N__17340),
            .in3(N__17388),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_4_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_4_20_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Commands_frame_decoder.WDT_RNID7P31_6_LC_4_20_3  (
            .in0(N__15597),
            .in1(N__15583),
            .in2(_gnd_net_),
            .in3(N__15567),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_4_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_4_20_4 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_4_20_4  (
            .in0(N__15553),
            .in1(N__15538),
            .in2(N__15532),
            .in3(N__15529),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_4_20_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_4_20_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_4_20_5  (
            .in0(N__17389),
            .in1(N__17326),
            .in2(_gnd_net_),
            .in3(N__17279),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_4_20_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_4_20_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_4_20_6  (
            .in0(N__17280),
            .in1(_gnd_net_),
            .in2(N__17341),
            .in3(N__17390),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_4_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_4_21_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_4_21_2 .LUT_INIT=16'b1110010011110100;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_4_21_2  (
            .in0(N__22510),
            .in1(N__15631),
            .in2(N__15507),
            .in3(N__17956),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29317),
            .ce(),
            .sr(N__28758));
    defparam \ppm_encoder_1.aileron_8_LC_4_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_4_21_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_4_21_7  (
            .in0(N__22477),
            .in1(N__24091),
            .in2(N__24798),
            .in3(N__15483),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29317),
            .ce(),
            .sr(N__28758));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_4_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_4_22_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_4_22_1  (
            .in0(N__22828),
            .in1(N__15455),
            .in2(_gnd_net_),
            .in3(N__19615),
            .lcout(),
            .ltout(\ppm_encoder_1.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2  (
            .in0(_gnd_net_),
            .in1(N__20934),
            .in2(N__15646),
            .in3(N__19876),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_4_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_4_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__18969),
            .in2(_gnd_net_),
            .in3(N__18935),
            .lcout(\ppm_encoder_1.N_139_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_5_LC_4_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_5_LC_4_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_5_LC_4_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_5_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24265),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29300),
            .ce(N__25042),
            .sr(N__28772));
    defparam \ppm_encoder_1.elevator_esr_5_LC_4_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_5_LC_4_23_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_5_LC_4_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_5_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24250),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29300),
            .ce(N__25042),
            .sr(N__28772));
    defparam \ppm_encoder_1.rudder_esr_5_LC_4_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_4_23_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_4_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24232),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29300),
            .ce(N__25042),
            .sr(N__28772));
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_4_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_4_24_0 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_4_24_0  (
            .in0(N__18295),
            .in1(_gnd_net_),
            .in2(N__15625),
            .in3(N__15604),
            .lcout(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_4_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_4_24_1 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNIU0DH2_10_LC_4_24_1  (
            .in0(N__22683),
            .in1(N__16061),
            .in2(N__19963),
            .in3(N__15993),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_4_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_4_24_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_4_24_2  (
            .in0(N__15994),
            .in1(N__25099),
            .in2(N__16066),
            .in3(N__22387),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_4_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_4_24_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNIG4JI2_11_LC_4_24_3  (
            .in0(N__17919),
            .in1(N__19710),
            .in2(N__15883),
            .in3(N__15770),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_4_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_4_24_4 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIALRT5_11_LC_4_24_4  (
            .in0(N__16105),
            .in1(_gnd_net_),
            .in2(N__16081),
            .in3(N__15922),
            .lcout(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_4_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_4_24_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI03DH2_11_LC_4_24_5  (
            .in0(N__24675),
            .in1(N__16060),
            .in2(N__17898),
            .in3(N__15992),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_4_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_4_24_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_4_24_7  (
            .in0(N__16148),
            .in1(N__20559),
            .in2(_gnd_net_),
            .in3(N__19711),
            .lcout(\ppm_encoder_1.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_25_0 .LUT_INIT=16'b1111010111000101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_25_0  (
            .in0(N__20004),
            .in1(N__20551),
            .in2(N__20351),
            .in3(N__16243),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_25_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_4_25_1  (
            .in0(N__20553),
            .in1(N__20322),
            .in2(N__15916),
            .in3(N__20005),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_4_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_4_25_2 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_4_25_2  (
            .in0(N__20323),
            .in1(N__20552),
            .in2(N__16193),
            .in3(N__19639),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_4_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_4_25_4 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIE2JI2_10_LC_4_25_4  (
            .in0(N__22713),
            .in1(N__19638),
            .in2(N__15882),
            .in3(N__15761),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_4_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_4_25_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI5GRT5_10_LC_4_25_5  (
            .in0(N__15688),
            .in1(_gnd_net_),
            .in2(N__15670),
            .in3(N__15667),
            .lcout(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_4_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_4_25_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_4_25_6  (
            .in0(N__20327),
            .in1(_gnd_net_),
            .in2(N__20010),
            .in3(N__15652),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_4_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_4_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_4_25_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_4_25_7  (
            .in0(_gnd_net_),
            .in1(N__24797),
            .in2(_gnd_net_),
            .in3(N__28925),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_4_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_4_26_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_4_26_0  (
            .in0(N__17823),
            .in1(N__16326),
            .in2(N__18570),
            .in3(N__18937),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_4_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_4_26_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_4_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16288),
            .in3(N__18968),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_4_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_4_26_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_4_26_2 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_4_26_2  (
            .in0(N__16285),
            .in1(N__18049),
            .in2(N__16279),
            .in3(N__16276),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29279),
            .ce(),
            .sr(N__28781));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_4_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_4_26_3 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_4_26_3  (
            .in0(N__16239),
            .in1(_gnd_net_),
            .in2(N__23799),
            .in3(N__20714),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_4_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_4_26_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_4_26_4  (
            .in0(N__20713),
            .in1(N__23733),
            .in2(_gnd_net_),
            .in3(N__16238),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_4_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_4_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_4_26_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_4_26_5  (
            .in0(N__18198),
            .in1(N__16213),
            .in2(N__18079),
            .in3(N__16201),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29279),
            .ce(),
            .sr(N__28781));
    defparam \ppm_encoder_1.init_pulses_11_LC_4_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_4_26_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_4_26_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_4_26_6  (
            .in0(N__18200),
            .in1(N__18045),
            .in2(N__16171),
            .in3(N__16156),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29279),
            .ce(),
            .sr(N__28781));
    defparam \ppm_encoder_1.init_pulses_12_LC_4_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_4_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_4_26_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_4_26_7  (
            .in0(N__18199),
            .in1(N__16123),
            .in2(N__18080),
            .in3(N__16111),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29279),
            .ce(),
            .sr(N__28781));
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_4_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_4_27_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_4_27_0  (
            .in0(N__23788),
            .in1(N__23885),
            .in2(N__20809),
            .in3(N__16458),
            .lcout(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_4_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_4_27_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_4_27_1  (
            .in0(N__18205),
            .in1(N__18090),
            .in2(N__16492),
            .in3(N__16477),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29272),
            .ce(),
            .sr(N__28783));
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_4_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_4_27_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_4_27_2  (
            .in0(N__23784),
            .in1(N__23886),
            .in2(_gnd_net_),
            .in3(N__20784),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_4_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_4_27_3 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_4_27_3  (
            .in0(N__16459),
            .in1(N__17552),
            .in2(N__20806),
            .in3(N__23787),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_4_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_4_27_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_4_27_4  (
            .in0(N__18202),
            .in1(N__16399),
            .in2(N__18111),
            .in3(N__16387),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29272),
            .ce(),
            .sr(N__28783));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_4_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_4_27_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_4_27_5  (
            .in0(N__20786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23786),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_4_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_4_27_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_4_27_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_4_27_6  (
            .in0(N__18201),
            .in1(N__16369),
            .in2(N__18110),
            .in3(N__16357),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29272),
            .ce(),
            .sr(N__28783));
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_4_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_4_27_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISFRP_13_LC_4_27_7  (
            .in0(N__20785),
            .in1(N__21032),
            .in2(_gnd_net_),
            .in3(N__23785),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_28_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_28_0  (
            .in0(N__16555),
            .in1(N__22633),
            .in2(N__16549),
            .in3(N__22612),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_28_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_4_28_1  (
            .in0(N__23096),
            .in1(_gnd_net_),
            .in2(N__16579),
            .in3(N__16567),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29268),
            .ce(N__23052),
            .sr(N__28788));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_28_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_4_28_2  (
            .in0(N__18394),
            .in1(N__18496),
            .in2(_gnd_net_),
            .in3(N__23097),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29268),
            .ce(N__23052),
            .sr(N__28788));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_4_28_3  (
            .in0(N__23093),
            .in1(N__19933),
            .in2(_gnd_net_),
            .in3(N__16540),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29268),
            .ce(N__23052),
            .sr(N__28788));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_28_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_28_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_4_28_5  (
            .in0(N__23094),
            .in1(N__17872),
            .in2(_gnd_net_),
            .in3(N__16531),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29268),
            .ce(N__23052),
            .sr(N__28788));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_4_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_4_28_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_4_28_6  (
            .in0(N__16522),
            .in1(N__23095),
            .in2(_gnd_net_),
            .in3(N__19975),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29268),
            .ce(N__23052),
            .sr(N__28788));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_4_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_4_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_4_29_0  (
            .in0(_gnd_net_),
            .in1(N__18778),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_29_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_4_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_4_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_4_29_1  (
            .in0(_gnd_net_),
            .in1(N__18445),
            .in2(N__27272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_4_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_4_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_4_29_2  (
            .in0(_gnd_net_),
            .in1(N__16510),
            .in2(N__27266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_4_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_4_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_4_29_3  (
            .in0(_gnd_net_),
            .in1(N__23236),
            .in2(N__27269),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_4_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_4_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_4_29_4  (
            .in0(_gnd_net_),
            .in1(N__16609),
            .in2(N__27267),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_4_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_4_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_4_29_5  (
            .in0(_gnd_net_),
            .in1(N__18724),
            .in2(N__27270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_4_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_4_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_4_29_6  (
            .in0(_gnd_net_),
            .in1(N__18712),
            .in2(N__27268),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_4_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_4_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_4_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_4_29_7  (
            .in0(_gnd_net_),
            .in1(N__22978),
            .in2(N__27271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_4_30_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_4_30_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_4_30_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_4_30_0  (
            .in0(_gnd_net_),
            .in1(N__18847),
            .in2(N__27274),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_30_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_4_30_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_4_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_4_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_4_30_1  (
            .in0(_gnd_net_),
            .in1(N__18853),
            .in2(N__27275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_4_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_4_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_4_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16600),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_5_10_1 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_5_10_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_5_10_1  (
            .in0(N__16781),
            .in1(N__16699),
            .in2(_gnd_net_),
            .in3(N__16595),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29377),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI08RE_4_LC_5_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI08RE_4_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI08RE_4_LC_5_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI08RE_4_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__16852),
            .in2(_gnd_net_),
            .in3(N__29618),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_5_12_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_5_12_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_5_12_3  (
            .in0(N__16837),
            .in1(N__16825),
            .in2(N__16813),
            .in3(N__16795),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_5_12_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_5_12_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_5_12_6  (
            .in0(N__19092),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__26608),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_5_13_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_5_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_5_13_2  (
            .in0(N__16756),
            .in1(N__16741),
            .in2(N__16729),
            .in3(N__16714),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_5_13_3 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_5_13_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \uart_pc.data_0_LC_5_13_3  (
            .in0(N__16971),
            .in1(N__17041),
            .in2(N__29826),
            .in3(N__17212),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29366),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNIVM1O_6_LC_5_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIVM1O_6_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIVM1O_6_LC_5_13_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_1_RNIVM1O_6_LC_5_13_5  (
            .in0(N__25616),
            .in1(N__29600),
            .in2(_gnd_net_),
            .in3(N__28926),
            .lcout(\Commands_frame_decoder.state_1_RNIVM1OZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI19RE_5_LC_5_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI19RE_5_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI19RE_5_LC_5_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI19RE_5_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__16944),
            .in2(_gnd_net_),
            .in3(N__29587),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_6_LC_5_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_6_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_6_LC_5_14_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_1_6_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__25612),
            .in2(N__16633),
            .in3(N__29459),
            .lcout(\Commands_frame_decoder.state_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29361),
            .ce(),
            .sr(N__28717));
    defparam \Commands_frame_decoder.source_offset1data_4_LC_5_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset1data_4_LC_5_14_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset1data_4_LC_5_14_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_offset1data_4_LC_5_14_2  (
            .in0(N__16623),
            .in1(N__29588),
            .in2(N__25617),
            .in3(N__27972),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29361),
            .ce(),
            .sr(N__28717));
    defparam \Commands_frame_decoder.state_1_5_LC_5_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_5_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_5_LC_5_14_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_1_5_LC_5_14_3  (
            .in0(N__16945),
            .in1(N__24652),
            .in2(_gnd_net_),
            .in3(N__29458),
            .lcout(\Commands_frame_decoder.state_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29361),
            .ce(),
            .sr(N__28717));
    defparam \uart_pc.data_rdy_LC_5_14_5 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_5_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.data_rdy_LC_5_14_5  (
            .in0(N__19132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19338),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29361),
            .ce(),
            .sr(N__28717));
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_0_LC_5_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_0_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_ns_i_a2_3_0_LC_5_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_1_ns_i_a2_3_0_LC_5_15_0  (
            .in0(N__29591),
            .in1(N__28076),
            .in2(N__28175),
            .in3(N__16936),
            .lcout(\Commands_frame_decoder.N_323 ),
            .ltout(\Commands_frame_decoder.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_2_LC_5_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_2_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_2_LC_5_15_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_1_2_LC_5_15_1  (
            .in0(N__16906),
            .in1(N__16927),
            .in2(N__16921),
            .in3(N__29455),
            .lcout(\Commands_frame_decoder.state_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29354),
            .ce(),
            .sr(N__28722));
    defparam \Commands_frame_decoder.state_1_RNIRI1O_2_LC_5_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIRI1O_2_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIRI1O_2_LC_5_15_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_1_RNIRI1O_2_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__16878),
            .in2(_gnd_net_),
            .in3(N__28938),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNIU5RE_2_LC_5_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIU5RE_2_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIU5RE_2_LC_5_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNIU5RE_2_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__16905),
            .in2(_gnd_net_),
            .in3(N__29589),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_3_LC_5_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_3_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_3_LC_5_15_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \Commands_frame_decoder.state_1_3_LC_5_15_4  (
            .in0(N__29456),
            .in1(_gnd_net_),
            .in2(N__16867),
            .in3(N__16864),
            .lcout(\Commands_frame_decoder.state_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29354),
            .ce(),
            .sr(N__28722));
    defparam \Commands_frame_decoder.state_1_RNIV6RE_3_LC_5_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIV6RE_3_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIV6RE_3_LC_5_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNIV6RE_3_LC_5_15_6  (
            .in0(N__29590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16863),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_4_LC_5_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_4_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_4_LC_5_15_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_1_4_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__16851),
            .in2(N__16855),
            .in3(N__29457),
            .lcout(\Commands_frame_decoder.state_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29354),
            .ce(),
            .sr(N__28722));
    defparam \uart_drone.data_Aux_5_LC_5_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_5_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_5_16_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_5_LC_5_16_1  (
            .in0(N__19165),
            .in1(N__21746),
            .in2(N__17089),
            .in3(N__21775),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29348),
            .ce(),
            .sr(N__21586));
    defparam \uart_drone.data_Aux_6_LC_5_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_5_16_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_5_16_3  (
            .in0(N__19228),
            .in1(N__21747),
            .in2(N__17074),
            .in3(N__21776),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29348),
            .ce(),
            .sr(N__21586));
    defparam \uart_drone.data_Aux_7_LC_5_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_5_16_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_5_16_4  (
            .in0(N__21777),
            .in1(N__21748),
            .in2(N__17059),
            .in3(N__25525),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29348),
            .ce(),
            .sr(N__21586));
    defparam \uart_pc.data_2_LC_5_17_0 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_5_17_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_2_LC_5_17_0  (
            .in0(N__17025),
            .in1(N__16994),
            .in2(N__17158),
            .in3(N__28307),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29342),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_5_17_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_5_17_1 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \uart_drone.timer_Count_0_LC_5_17_1  (
            .in0(N__21552),
            .in1(N__17516),
            .in2(N__19278),
            .in3(N__26625),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29342),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_5_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_5_17_2 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_5_17_2  (
            .in0(N__29614),
            .in1(N__22338),
            .in2(N__17443),
            .in3(N__22305),
            .lcout(\Commands_frame_decoder.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_17_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__17515),
            .in2(_gnd_net_),
            .in3(N__17535),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_5_17_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_5_17_4 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_drone.timer_Count_1_LC_5_17_4  (
            .in0(N__26624),
            .in1(N__19274),
            .in2(N__17044),
            .in3(N__21553),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29342),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_5_17_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_5_17_5 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_5_17_5  (
            .in0(N__19191),
            .in1(N__25582),
            .in2(N__17497),
            .in3(N__21887),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_5_17_6 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_5_17_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_6_LC_5_17_6  (
            .in0(N__17026),
            .in1(N__16995),
            .in2(N__17626),
            .in3(N__27577),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29342),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_4_0_LC_5_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_4_0_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_4_0_LC_5_17_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_4_0_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__17439),
            .in2(_gnd_net_),
            .in3(N__29613),
            .lcout(\Commands_frame_decoder.state_1_RNO_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_5_18_0 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_5_18_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_drone.timer_Count_2_LC_5_18_0  (
            .in0(N__26622),
            .in1(N__17470),
            .in2(N__19291),
            .in3(N__21557),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29336),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_18_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_18_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_5_18_1  (
            .in0(N__17273),
            .in1(N__17398),
            .in2(_gnd_net_),
            .in3(N__17350),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_5_18_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_5_18_2 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_5_18_2  (
            .in0(N__21917),
            .in1(N__17483),
            .in2(N__21999),
            .in3(N__21888),
            .lcout(\uart_drone.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state49_i_LC_5_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state49_i_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state49_i_LC_5_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state49_i_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__29640),
            .in2(_gnd_net_),
            .in3(N__28929),
            .lcout(\Commands_frame_decoder.un1_state49_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_5_18_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_5_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_5_18_4  (
            .in0(N__21918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17484),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_5_18_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_5_18_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_5_18_5  (
            .in0(N__21889),
            .in1(N__21985),
            .in2(N__17095),
            .in3(N__26621),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_5_18_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_5_18_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_5_18_6  (
            .in0(N__19289),
            .in1(N__26626),
            .in2(N__17092),
            .in3(N__17461),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29336),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_5_18_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_5_18_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_4_LC_5_18_7  (
            .in0(N__17449),
            .in1(N__19290),
            .in2(N__21564),
            .in3(N__26623),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29336),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_19_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_19_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_5_19_0  (
            .in0(N__17520),
            .in1(N__17536),
            .in2(N__17521),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_19_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__17485),
            .in2(_gnd_net_),
            .in3(N__17464),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_19_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__21922),
            .in2(_gnd_net_),
            .in3(N__17455),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_19_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(N__21991),
            .in2(_gnd_net_),
            .in3(N__17452),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_5_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_5_19_4 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \Commands_frame_decoder.preinit_RNIF92K5_LC_5_19_4  (
            .in0(N__22330),
            .in1(N__17432),
            .in2(N__27388),
            .in3(N__22298),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_19_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_19_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_5_19_6  (
            .in0(N__17397),
            .in1(N__17349),
            .in2(_gnd_net_),
            .in3(N__17284),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_5_20_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_5_20_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_5_20_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_5_20_0  (
            .in0(N__17221),
            .in1(N__19133),
            .in2(N__17211),
            .in3(N__19428),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_1_LC_5_20_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_5_20_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_1_LC_5_20_1  (
            .in0(N__19429),
            .in1(N__17181),
            .in2(N__19152),
            .in3(N__17194),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_2_LC_5_20_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_5_20_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_5_20_2  (
            .in0(N__17170),
            .in1(N__19137),
            .in2(N__17154),
            .in3(N__19430),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_3_LC_5_20_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_5_20_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_5_20_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_3_LC_5_20_3  (
            .in0(N__19431),
            .in1(N__17688),
            .in2(N__19153),
            .in3(N__17704),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_4_LC_5_20_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_5_20_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_5_20_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_5_20_4  (
            .in0(N__17677),
            .in1(N__19141),
            .in2(N__17670),
            .in3(N__19432),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_5_LC_5_20_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_5_20_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_5_20_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_5_LC_5_20_5  (
            .in0(N__19433),
            .in1(N__17637),
            .in2(N__19154),
            .in3(N__17653),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_7_LC_5_20_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_5_20_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_5_20_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_7_LC_5_20_7  (
            .in0(N__19434),
            .in1(N__17616),
            .in2(N__19155),
            .in3(N__19378),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29318),
            .ce(),
            .sr(N__19581));
    defparam \uart_pc.data_Aux_6_LC_5_21_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_5_21_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_pc.data_Aux_6_LC_5_21_0  (
            .in0(N__19156),
            .in1(N__17605),
            .in2(N__17586),
            .in3(N__19435),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29308),
            .ce(),
            .sr(N__19585));
    defparam \ppm_encoder_1.pulses2count_18_LC_5_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_5_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_5_23_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_5_23_0  (
            .in0(N__23808),
            .in1(N__23850),
            .in2(N__17569),
            .in3(N__18867),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29290),
            .ce(),
            .sr(N__28766));
    defparam \ppm_encoder_1.rudder_7_LC_5_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_5_23_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_5_23_1 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_5_23_1  (
            .in0(N__19393),
            .in1(N__24867),
            .in2(N__20412),
            .in3(N__25468),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29290),
            .ce(),
            .sr(N__28766));
    defparam \ppm_encoder_1.rudder_6_LC_5_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_5_23_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_5_23_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_5_23_2  (
            .in0(N__24865),
            .in1(N__25132),
            .in2(_gnd_net_),
            .in3(N__21065),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29290),
            .ce(),
            .sr(N__28766));
    defparam \ppm_encoder_1.aileron_11_LC_5_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_5_23_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_5_23_3 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_5_23_3  (
            .in0(N__23965),
            .in1(N__24866),
            .in2(N__17899),
            .in3(N__22435),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29290),
            .ce(),
            .sr(N__28766));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_24_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_24_1  (
            .in0(N__21235),
            .in1(N__20224),
            .in2(N__21202),
            .in3(N__17952),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_5_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_5_24_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_5_24_2  (
            .in0(N__17923),
            .in1(_gnd_net_),
            .in2(N__22846),
            .in3(N__24676),
            .lcout(),
            .ltout(\ppm_encoder_1.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_5_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_5_24_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_5_24_3  (
            .in0(N__17894),
            .in1(_gnd_net_),
            .in2(N__17875),
            .in3(N__20948),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_24_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_24_6  (
            .in0(N__22815),
            .in1(N__17819),
            .in2(_gnd_net_),
            .in3(N__17859),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_5_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_5_24_7 .LUT_INIT=16'b0000010101010101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_5_24_7  (
            .in0(N__17860),
            .in1(_gnd_net_),
            .in2(N__17824),
            .in3(N__22816),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_5_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_5_25_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_5_25_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_5_25_0  (
            .in0(N__18209),
            .in1(N__17773),
            .in2(N__18114),
            .in3(N__17761),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29280),
            .ce(),
            .sr(N__28775));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_5_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_5_25_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_5_25_1  (
            .in0(N__18405),
            .in1(_gnd_net_),
            .in2(N__23823),
            .in3(N__20775),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_5_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_5_25_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_5_25_2  (
            .in0(N__20774),
            .in1(N__18404),
            .in2(_gnd_net_),
            .in3(N__23800),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_5_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_5_25_3 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_5_25_3  (
            .in0(N__17719),
            .in1(N__20321),
            .in2(N__18409),
            .in3(N__20569),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_6_LC_5_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_5_25_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_5_25_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_5_25_4  (
            .in0(N__18210),
            .in1(N__18385),
            .in2(N__18115),
            .in3(N__18370),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29280),
            .ce(),
            .sr(N__28775));
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_5_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_5_25_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIERUS_6_LC_5_25_5  (
            .in0(N__21089),
            .in1(_gnd_net_),
            .in2(N__23824),
            .in3(N__20776),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_5_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_5_25_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_5_25_7 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_5_25_7  (
            .in0(N__18340),
            .in1(N__18107),
            .in2(N__18328),
            .in3(N__18211),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29280),
            .ce(),
            .sr(N__28775));
    defparam \ppm_encoder_1.init_pulses_14_LC_5_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_5_26_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_5_26_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_5_26_0  (
            .in0(N__18203),
            .in1(N__18316),
            .in2(N__18108),
            .in3(N__18304),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29273),
            .ce(),
            .sr(N__28778));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_5_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_5_26_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_14_LC_5_26_1  (
            .in0(N__19913),
            .in1(N__23749),
            .in2(_gnd_net_),
            .in3(N__20780),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_5_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_5_26_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_5_26_2  (
            .in0(N__20778),
            .in1(_gnd_net_),
            .in2(N__23807),
            .in3(N__19914),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_5_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_5_26_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_5_26_5  (
            .in0(N__22968),
            .in1(N__23748),
            .in2(_gnd_net_),
            .in3(N__20779),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_5_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_5_26_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_5_26_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_5_26_6  (
            .in0(N__18204),
            .in1(N__18130),
            .in2(N__18109),
            .in3(N__17968),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29273),
            .ce(),
            .sr(N__28778));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_5_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_5_26_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_4_LC_5_26_7  (
            .in0(N__18666),
            .in1(N__23744),
            .in2(_gnd_net_),
            .in3(N__20777),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_5_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_5_27_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_5_27_0  (
            .in0(N__22849),
            .in1(N__20922),
            .in2(_gnd_net_),
            .in3(N__18637),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_5_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_5_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_5_27_2  (
            .in0(N__18616),
            .in1(N__18589),
            .in2(_gnd_net_),
            .in3(N__18571),
            .lcout(),
            .ltout(\ppm_encoder_1.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_5_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_5_27_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_5_27_3  (
            .in0(N__20923),
            .in1(_gnd_net_),
            .in2(N__18517),
            .in3(N__18514),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_27_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_27_5  (
            .in0(N__20924),
            .in1(N__22848),
            .in2(_gnd_net_),
            .in3(N__18490),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_27_7 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_27_7  (
            .in0(N__20360),
            .in1(N__20537),
            .in2(N__20017),
            .in3(N__18469),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_28_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_28_1  (
            .in0(N__21231),
            .in1(N__18928),
            .in2(N__21198),
            .in3(N__20220),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_28_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_28_2  (
            .in0(N__18415),
            .in1(N__21191),
            .in2(N__18814),
            .in3(N__21230),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_5_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_5_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_5_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_5_28_3  (
            .in0(N__23125),
            .in1(N__18439),
            .in2(_gnd_net_),
            .in3(N__18427),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29265),
            .ce(N__23060),
            .sr(N__28784));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_5_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_5_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_5_28_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_5_28_4  (
            .in0(N__18829),
            .in1(N__23126),
            .in2(_gnd_net_),
            .in3(N__18820),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29265),
            .ce(N__23060),
            .sr(N__28784));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_5_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_5_28_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_5_28_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_5_28_5  (
            .in0(N__23123),
            .in1(_gnd_net_),
            .in2(N__18805),
            .in3(N__18796),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29265),
            .ce(N__23060),
            .sr(N__28784));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_28_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_28_6  (
            .in0(N__20219),
            .in1(N__18784),
            .in2(N__18748),
            .in3(N__20244),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_5_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_5_28_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_5_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_5_28_7  (
            .in0(N__23124),
            .in1(N__18772),
            .in2(_gnd_net_),
            .in3(N__18760),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29265),
            .ce(N__23060),
            .sr(N__28784));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_5_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_5_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_5_29_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_5_29_0  (
            .in0(N__18739),
            .in1(N__21297),
            .in2(N__18733),
            .in3(N__21123),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_5_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_5_29_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_5_29_2  (
            .in0(N__23314),
            .in1(N__18718),
            .in2(N__23170),
            .in3(N__22570),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_29_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_5_29_5  (
            .in0(N__21124),
            .in1(N__21148),
            .in2(N__21301),
            .in3(N__20248),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_5_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_5_29_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_5_29_6  (
            .in0(N__23386),
            .in1(N__18706),
            .in2(N__18697),
            .in3(N__22546),
            .lcout(\ppm_encoder_1.N_237 ),
            .ltout(\ppm_encoder_1.N_237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_29_7 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_29_7  (
            .in0(N__26642),
            .in1(N__18958),
            .in2(N__18940),
            .in3(N__18936),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_5_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_5_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_5_30_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_5_30_1  (
            .in0(_gnd_net_),
            .in1(N__18868),
            .in2(_gnd_net_),
            .in3(N__23427),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_30_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_30_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_30_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_30_6  (
            .in0(N__22939),
            .in1(N__23470),
            .in2(N__22897),
            .in3(N__23449),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_7_1_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_7_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_7_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_7_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23353),
            .lcout(\uart_pc_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29392),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_7_2_2 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_7_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18835),
            .lcout(uart_commands_input_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29390),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_7_2_4 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_7_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18841),
            .lcout(\uart_pc_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29390),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_7_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_7_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(frame_decoder_CH2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29367),
            .ce(N__21339),
            .sr(N__28711));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_7_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_7_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27871),
            .lcout(frame_decoder_CH2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_7_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_7_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28221),
            .lcout(frame_decoder_CH2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_7_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_7_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27989),
            .lcout(frame_decoder_CH2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_7_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_7_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27736),
            .lcout(frame_decoder_CH2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_7_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_7_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28105),
            .lcout(frame_decoder_CH2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_7_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_7_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28354),
            .lcout(frame_decoder_CH2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29355),
            .ce(N__21338),
            .sr(N__28715));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_7_14_1 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_7_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_7_14_1  (
            .in0(N__26348),
            .in1(N__26271),
            .in2(_gnd_net_),
            .in3(N__26109),
            .lcout(\uart_drone.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNIUL1O_5_LC_7_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIUL1O_5_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIUL1O_5_LC_7_14_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_1_RNIUL1O_5_LC_7_14_3  (
            .in0(N__19018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28935),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNISJ1O_3_LC_7_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNISJ1O_3_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNISJ1O_3_LC_7_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_1_RNISJ1O_3_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__19009),
            .in2(_gnd_net_),
            .in3(N__28936),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_7_15_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_7_15_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_7_15_0  (
            .in0(N__21619),
            .in1(N__21754),
            .in2(N__18994),
            .in3(N__28948),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_7_15_1 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_7_15_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_7_15_1  (
            .in0(N__18993),
            .in1(N__22020),
            .in2(N__18997),
            .in3(N__21944),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29343),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_7_15_2 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_7_15_2 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \uart_drone.state_1_LC_7_15_2  (
            .in0(N__18992),
            .in1(N__19177),
            .in2(N__28981),
            .in3(N__21755),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29343),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_7_15_3 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_7_15_3 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.state_1_LC_7_15_3  (
            .in0(N__28949),
            .in1(N__19038),
            .in2(N__19213),
            .in3(N__19104),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29343),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_7_15_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_7_15_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_7_15_7  (
            .in0(N__26353),
            .in1(N__26273),
            .in2(_gnd_net_),
            .in3(N__26111),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_7_16_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_7_16_0 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_7_16_0  (
            .in0(N__19209),
            .in1(N__19094),
            .in2(_gnd_net_),
            .in3(N__28946),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_7_16_1 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_7_16_1 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_pc.state_0_LC_7_16_1  (
            .in0(N__22242),
            .in1(N__19528),
            .in2(N__19216),
            .in3(N__19513),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29337),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_7_16_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_7_16_2 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_7_16_2  (
            .in0(N__21750),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__28945),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_7_16_3 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_7_16_3 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_7_16_3  (
            .in0(N__19198),
            .in1(N__22019),
            .in2(N__19180),
            .in3(N__21881),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29337),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_7_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_7_16_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_7_16_4  (
            .in0(N__26341),
            .in1(N__26272),
            .in2(_gnd_net_),
            .in3(N__26110),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_2_LC_7_16_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_7_16_6 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_7_16_6  (
            .in0(N__19250),
            .in1(N__19093),
            .in2(N__19039),
            .in3(N__28947),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_7_16_7 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_7_16_7 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_pc.state_2_LC_7_16_7  (
            .in0(N__22243),
            .in1(N__19037),
            .in2(N__19021),
            .in3(N__22060),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29337),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_7_17_0 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_7_17_0 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_pc.state_3_LC_7_17_0  (
            .in0(N__19249),
            .in1(N__19348),
            .in2(N__19300),
            .in3(N__26694),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29328),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_17_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_17_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_7_17_1  (
            .in0(N__22053),
            .in1(_gnd_net_),
            .in2(N__22240),
            .in3(N__19377),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(\uart_pc.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_7_17_2 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_7_17_2 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \uart_pc.state_4_LC_7_17_2  (
            .in0(N__22118),
            .in1(N__19475),
            .in2(N__19342),
            .in3(N__26695),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29328),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_17_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_17_3 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_7_17_3  (
            .in0(N__22052),
            .in1(N__22271),
            .in2(N__22239),
            .in3(N__19508),
            .lcout(\uart_pc.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_7_17_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_7_17_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_7_17_4  (
            .in0(N__22230),
            .in1(N__22054),
            .in2(N__19251),
            .in3(N__19474),
            .lcout(\uart_pc.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_7_17_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_7_17_5 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_7_17_5  (
            .in0(N__25567),
            .in1(N__22014),
            .in2(N__21630),
            .in3(N__21946),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_17_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_17_6 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_7_17_6  (
            .in0(N__22231),
            .in1(N__22055),
            .in2(N__19252),
            .in3(N__19473),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_7_17_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_7_17_7 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_7_17_7  (
            .in0(N__25566),
            .in1(N__22015),
            .in2(N__21629),
            .in3(N__21945),
            .lcout(\uart_drone.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_7_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_7_18_0  (
            .in0(N__19524),
            .in1(N__19510),
            .in2(N__22238),
            .in3(N__26683),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_7_18_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_7_18_1 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_2_LC_7_18_1  (
            .in0(N__26685),
            .in1(N__22083),
            .in2(N__19588),
            .in3(N__22255),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29319),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_7_18_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_18_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_7_18_2  (
            .in0(N__19472),
            .in1(N__19512),
            .in2(_gnd_net_),
            .in3(N__28928),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_7_18_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_7_18_3 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_pc.timer_Count_4_LC_7_18_3  (
            .in0(N__26686),
            .in1(N__22180),
            .in2(N__22092),
            .in3(N__22117),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29319),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_7_18_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_18_4 .LUT_INIT=16'b0000000010110011;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_7_18_4  (
            .in0(N__22050),
            .in1(N__19465),
            .in2(N__22237),
            .in3(N__19509),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_7_18_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_7_18_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \uart_pc.timer_Count_0_LC_7_18_5  (
            .in0(N__26684),
            .in1(N__22084),
            .in2(N__22174),
            .in3(N__22116),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29319),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_7_18_6  (
            .in0(N__22051),
            .in1(N__22272),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_18_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_18_7 .LUT_INIT=16'b1010111011101110;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_7_18_7  (
            .in0(N__19511),
            .in1(N__19471),
            .in2(N__19438),
            .in3(N__22282),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__25131),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__25461),
            .in2(_gnd_net_),
            .in3(N__19381),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__25437),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__25413),
            .in2(_gnd_net_),
            .in3(N__19666),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__25389),
            .in2(_gnd_net_),
            .in3(N__19663),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__25365),
            .in2(_gnd_net_),
            .in3(N__19660),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__25341),
            .in2(_gnd_net_),
            .in3(N__19657),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__25314),
            .in2(N__27276),
            .in3(N__19654),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_7_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__25291),
            .in2(_gnd_net_),
            .in3(N__19651),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29301),
            .ce(N__25076),
            .sr(N__28746));
    defparam \ppm_encoder_1.rudder_10_LC_7_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_7_21_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_7_21_0  (
            .in0(N__19648),
            .in1(N__25393),
            .in2(N__19637),
            .in3(N__24950),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.elevator_9_LC_7_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_7_21_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_7_21_2  (
            .in0(N__24553),
            .in1(N__25915),
            .in2(N__19613),
            .in3(N__24949),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.aileron_10_LC_7_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_7_21_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_7_21_3  (
            .in0(N__24010),
            .in1(N__22450),
            .in2(N__24964),
            .in3(N__19952),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.aileron_9_LC_7_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_7_21_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_7_21_4  (
            .in0(N__22462),
            .in1(N__24052),
            .in2(N__19874),
            .in3(N__24947),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.rudder_8_LC_7_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_7_21_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_7_21_5  (
            .in0(N__19843),
            .in1(N__25441),
            .in2(N__24965),
            .in3(N__19817),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.elevator_8_LC_7_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_7_21_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_7_21_6  (
            .in0(N__24568),
            .in1(N__25939),
            .in2(N__19796),
            .in3(N__24948),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29291),
            .ce(),
            .sr(N__28752));
    defparam \ppm_encoder_1.rudder_9_LC_7_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_7_22_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_7_22_0  (
            .in0(N__19765),
            .in1(N__25417),
            .in2(N__19748),
            .in3(N__24940),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29284),
            .ce(),
            .sr(N__28759));
    defparam \ppm_encoder_1.rudder_11_LC_7_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_7_22_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_7_22_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_7_22_2  (
            .in0(N__25369),
            .in1(N__19720),
            .in2(N__19709),
            .in3(N__24938),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29284),
            .ce(),
            .sr(N__28759));
    defparam \ppm_encoder_1.rudder_12_LC_7_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_7_22_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_7_22_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_7_22_3  (
            .in0(N__25345),
            .in1(N__19687),
            .in2(N__24963),
            .in3(N__20039),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29284),
            .ce(),
            .sr(N__28759));
    defparam \ppm_encoder_1.rudder_13_LC_7_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_7_22_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_7_22_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_7_22_4  (
            .in0(N__25321),
            .in1(N__19678),
            .in2(N__21015),
            .in3(N__24939),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29284),
            .ce(),
            .sr(N__28759));
    defparam \ppm_encoder_1.aileron_13_LC_7_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_7_22_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_7_22_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_7_22_7  (
            .in0(N__22402),
            .in1(N__24307),
            .in2(N__24962),
            .in3(N__20087),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29284),
            .ce(),
            .sr(N__28759));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_7_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_7_23_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_7_23_3  (
            .in0(N__25098),
            .in1(N__22850),
            .in2(_gnd_net_),
            .in3(N__20191),
            .lcout(),
            .ltout(\ppm_encoder_1.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_7_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_7_23_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__20960),
            .in2(N__20170),
            .in3(N__22386),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_7_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_7_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_7_23_5  (
            .in0(N__20961),
            .in1(N__20167),
            .in2(_gnd_net_),
            .in3(N__20155),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_7_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_7_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_7_24_0  (
            .in0(N__22851),
            .in1(N__20137),
            .in2(_gnd_net_),
            .in3(N__25005),
            .lcout(),
            .ltout(\ppm_encoder_1.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_7_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_7_24_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_7_24_1  (
            .in0(N__20962),
            .in1(_gnd_net_),
            .in2(N__20098),
            .in3(N__20091),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_24_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_24_4  (
            .in0(N__20544),
            .in1(N__20068),
            .in2(_gnd_net_),
            .in3(N__20041),
            .lcout(),
            .ltout(\ppm_encoder_1.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_7_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_7_24_5 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__20009),
            .in2(N__19978),
            .in3(N__20345),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_25_1  (
            .in0(N__20947),
            .in1(N__22657),
            .in2(_gnd_net_),
            .in3(N__19962),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_7_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_7_26_2 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_7_26_2  (
            .in0(N__20514),
            .in1(N__19918),
            .in2(N__20379),
            .in3(N__19896),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_26_7 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_26_7  (
            .in0(N__20517),
            .in1(N__21103),
            .in2(N__21076),
            .in3(N__20365),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_27_0 .LUT_INIT=16'b1110111101001111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_7_27_0  (
            .in0(N__20515),
            .in1(N__21042),
            .in2(N__20380),
            .in3(N__21014),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_7_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_7_27_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23821),
            .lcout(\ppm_encoder_1.N_590_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_27_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_27_5  (
            .in0(N__22858),
            .in1(N__20920),
            .in2(N__20545),
            .in3(N__20808),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_7_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_7_27_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_7_27_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_7_27_6  (
            .in0(N__20516),
            .in1(N__26707),
            .in2(N__20575),
            .in3(N__23822),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29264),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_7_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_7_27_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_7_27_7  (
            .in0(N__20513),
            .in1(N__20440),
            .in2(N__20416),
            .in3(N__20369),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_0_LC_7_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_7_28_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_7_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__20243),
            .in2(N__20265),
            .in3(N__20266),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_1_LC_7_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_7_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_7_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__20218),
            .in2(_gnd_net_),
            .in3(N__20194),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_2_LC_7_28_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_7_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_7_28_2  (
            .in0(_gnd_net_),
            .in1(N__21229),
            .in2(_gnd_net_),
            .in3(N__21205),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_3_LC_7_28_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_7_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_7_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_7_28_3  (
            .in0(_gnd_net_),
            .in1(N__21190),
            .in2(_gnd_net_),
            .in3(N__21166),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_4_LC_7_28_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_7_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_7_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_7_28_4  (
            .in0(_gnd_net_),
            .in1(N__22611),
            .in2(_gnd_net_),
            .in3(N__21163),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_5_LC_7_28_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_7_28_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_7_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_7_28_5  (
            .in0(_gnd_net_),
            .in1(N__22632),
            .in2(_gnd_net_),
            .in3(N__21160),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_6_LC_7_28_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_7_28_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_7_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_7_28_6  (
            .in0(_gnd_net_),
            .in1(N__23254),
            .in2(_gnd_net_),
            .in3(N__21157),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_7_LC_7_28_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_7_28_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_7_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_7_28_7  (
            .in0(_gnd_net_),
            .in1(N__23286),
            .in2(_gnd_net_),
            .in3(N__21154),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__29262),
            .ce(),
            .sr(N__21256));
    defparam \ppm_encoder_1.counter_8_LC_7_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_7_29_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_7_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_7_29_0  (
            .in0(_gnd_net_),
            .in1(N__22590),
            .in2(_gnd_net_),
            .in3(N__21151),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_29_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_9_LC_7_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_7_29_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_7_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_7_29_1  (
            .in0(_gnd_net_),
            .in1(N__21146),
            .in2(_gnd_net_),
            .in3(N__21127),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_10_LC_7_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_7_29_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_7_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_7_29_2  (
            .in0(_gnd_net_),
            .in1(N__21122),
            .in2(_gnd_net_),
            .in3(N__21106),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_11_LC_7_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_7_29_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_7_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_7_29_3  (
            .in0(_gnd_net_),
            .in1(N__21296),
            .in2(_gnd_net_),
            .in3(N__21280),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_12_LC_7_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_7_29_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_7_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_7_29_4  (
            .in0(_gnd_net_),
            .in1(N__22569),
            .in2(_gnd_net_),
            .in3(N__21277),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_13_LC_7_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_7_29_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_7_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_7_29_5  (
            .in0(_gnd_net_),
            .in1(N__23313),
            .in2(_gnd_net_),
            .in3(N__21274),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_14_LC_7_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_7_29_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_7_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_7_29_6  (
            .in0(_gnd_net_),
            .in1(N__22996),
            .in2(_gnd_net_),
            .in3(N__21271),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_15_LC_7_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_7_29_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_7_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_7_29_7  (
            .in0(_gnd_net_),
            .in1(N__23404),
            .in2(_gnd_net_),
            .in3(N__21268),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__29261),
            .ce(),
            .sr(N__21255));
    defparam \ppm_encoder_1.counter_16_LC_7_30_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_7_30_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_7_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_7_30_0  (
            .in0(_gnd_net_),
            .in1(N__23448),
            .in2(_gnd_net_),
            .in3(N__21265),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_30_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__29259),
            .ce(),
            .sr(N__21254));
    defparam \ppm_encoder_1.counter_17_LC_7_30_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_7_30_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_7_30_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_7_30_1  (
            .in0(_gnd_net_),
            .in1(N__23469),
            .in2(_gnd_net_),
            .in3(N__21262),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__29259),
            .ce(),
            .sr(N__21254));
    defparam \ppm_encoder_1.counter_18_LC_7_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_7_30_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_7_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_7_30_2  (
            .in0(_gnd_net_),
            .in1(N__23426),
            .in2(_gnd_net_),
            .in3(N__21259),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29259),
            .ce(),
            .sr(N__21254));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_0 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21241),
            .lcout(\uart_drone_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29391),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_8_1_1 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21358),
            .lcout(\uart_drone_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29391),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_6 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21364),
            .lcout(\uart_drone_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29391),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21352),
            .lcout(\uart_drone_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29388),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_8_2_7 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_8_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21346),
            .lcout(uart_drone_input_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29388),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_10_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27647),
            .lcout(frame_decoder_CH2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29368),
            .ce(N__21340),
            .sr(N__28712));
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_8_11_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_8_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__23340),
            .in2(_gnd_net_),
            .in3(N__21309),
            .lcout(\scaler_2.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.N_521_i_l_ofx_LC_8_11_2 .C_ON=1'b0;
    defparam \scaler_2.N_521_i_l_ofx_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.N_521_i_l_ofx_LC_8_11_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \scaler_2.N_521_i_l_ofx_LC_8_11_2  (
            .in0(N__21310),
            .in1(_gnd_net_),
            .in2(N__23344),
            .in3(_gnd_net_),
            .lcout(\scaler_2.N_521_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_8_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_8_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_6_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28213),
            .lcout(frame_decoder_OFF2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29356),
            .ce(N__24625),
            .sr(N__28716));
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_8_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_8_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_3_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28114),
            .lcout(frame_decoder_OFF2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29356),
            .ce(N__24625),
            .sr(N__28716));
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_8_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_8_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_5_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27883),
            .lcout(frame_decoder_OFF2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29356),
            .ce(N__24625),
            .sr(N__28716));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_8_13_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_8_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__25198),
            .in2(N__25241),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_8_13_1 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__21466),
            .in2(N__23332),
            .in3(N__21457),
            .lcout(\scaler_2.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_0 ),
            .carryout(\scaler_2.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_8_13_2 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__21454),
            .in2(N__24181),
            .in3(N__21448),
            .lcout(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_1 ),
            .carryout(\scaler_2.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_8_13_3 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__21445),
            .in2(N__21439),
            .in3(N__21430),
            .lcout(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_2 ),
            .carryout(\scaler_2.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_8_13_4 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__21427),
            .in2(N__23323),
            .in3(N__21418),
            .lcout(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_3 ),
            .carryout(\scaler_2.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_8_13_5 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__21415),
            .in2(N__21409),
            .in3(N__21400),
            .lcout(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_4 ),
            .carryout(\scaler_2.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_8_13_6 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__21397),
            .in2(N__21391),
            .in3(N__21379),
            .lcout(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_5 ),
            .carryout(\scaler_2.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_8_13_7 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__21376),
            .in2(_gnd_net_),
            .in3(N__21367),
            .lcout(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_6 ),
            .carryout(\scaler_2.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_8_14_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_8_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__21520),
            .in2(N__27265),
            .in3(N__21511),
            .lcout(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_8_14_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_8_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21508),
            .lcout(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_8_14_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_8_14_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_8_14_4  (
            .in0(N__26349),
            .in1(N__26278),
            .in2(_gnd_net_),
            .in3(N__26113),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_ns_0_a4_0_0_1_LC_8_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_ns_0_a4_0_0_1_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_ns_0_a4_0_0_1_LC_8_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_ns_0_a4_0_0_1_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__27617),
            .in2(_gnd_net_),
            .in3(N__29827),
            .lcout(\Commands_frame_decoder.state_1_ns_0_a4_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_8_15_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_8_15_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_8_15_1  (
            .in0(N__25522),
            .in1(N__22021),
            .in2(_gnd_net_),
            .in3(N__21943),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_8_15_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_8_15_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_8_15_3  (
            .in0(N__26112),
            .in1(N__26340),
            .in2(_gnd_net_),
            .in3(N__26274),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_15_4 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_15_4  (
            .in0(N__25819),
            .in1(N__25861),
            .in2(_gnd_net_),
            .in3(N__26810),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_0_LC_8_16_0  (
            .in0(N__24214),
            .in1(N__21738),
            .in2(N__21504),
            .in3(N__21792),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29329),
            .ce(),
            .sr(N__21576));
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_8_16_1  (
            .in0(N__21793),
            .in1(N__26206),
            .in2(N__21483),
            .in3(N__21740),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29329),
            .ce(),
            .sr(N__21576));
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_8_16_2  (
            .in0(N__21847),
            .in1(N__21739),
            .in2(N__21840),
            .in3(N__21794),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29329),
            .ce(),
            .sr(N__21576));
    defparam \uart_drone.data_Aux_3_LC_8_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_8_16_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_8_16_5  (
            .in0(N__21795),
            .in1(N__21823),
            .in2(N__21813),
            .in3(N__21741),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29329),
            .ce(),
            .sr(N__21576));
    defparam \uart_drone.data_Aux_4_LC_8_16_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_8_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_8_16_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_4_LC_8_16_7  (
            .in0(N__21796),
            .in1(N__21637),
            .in2(N__21654),
            .in3(N__21742),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29329),
            .ce(),
            .sr(N__21576));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_8_17_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_8_17_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_8_17_0  (
            .in0(N__26243),
            .in1(N__26313),
            .in2(_gnd_net_),
            .in3(N__26095),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_0_1_LC_8_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_0_1_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_0_1_LC_8_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_0_1_LC_8_17_2  (
            .in0(N__28310),
            .in1(N__27853),
            .in2(N__24394),
            .in3(N__24448),
            .lcout(\Commands_frame_decoder.state_1_ns_0_a4_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_8_17_3 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_8_17_3 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \uart_drone.state_3_LC_8_17_3  (
            .in0(N__21531),
            .in1(N__21631),
            .in2(N__21598),
            .in3(N__26692),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29320),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_8_17_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_8_17_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_8_17_4  (
            .in0(N__25571),
            .in1(N__21880),
            .in2(_gnd_net_),
            .in3(N__28931),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_8_17_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_8_17_5 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_pc.timer_Count_1_LC_8_17_5  (
            .in0(N__22120),
            .in1(N__22091),
            .in2(N__22138),
            .in3(N__26693),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29320),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_8_17_6 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_8_17_6 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \uart_drone.state_4_LC_8_17_6  (
            .in0(N__26691),
            .in1(N__21565),
            .in2(N__25583),
            .in3(N__21532),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29320),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_1_0_LC_8_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_1_0_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_1_0_LC_8_17_7 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_1_0_LC_8_17_7  (
            .in0(N__22360),
            .in1(N__24393),
            .in2(N__22348),
            .in3(N__22309),
            .lcout(\Commands_frame_decoder.state_1_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_8_18_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_8_18_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_8_18_0  (
            .in0(N__22165),
            .in1(N__22149),
            .in2(N__22173),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_8_18_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_8_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__22273),
            .in2(_gnd_net_),
            .in3(N__22249),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_8_18_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_8_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__22056),
            .in2(_gnd_net_),
            .in3(N__22246),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_8_18_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_8_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__22241),
            .in2(_gnd_net_),
            .in3(N__22183),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_8_18_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_8_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_8_18_4  (
            .in0(N__22169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22150),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_8_18_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_8_18_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_3_LC_8_18_5  (
            .in0(N__22126),
            .in1(N__22119),
            .in2(N__22093),
            .in3(N__26696),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29309),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_8_18_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_8_18_7 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_8_18_7  (
            .in0(N__21998),
            .in1(N__21931),
            .in2(N__25578),
            .in3(N__21876),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_8_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_8_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_c_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__24162),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_8_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_8_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__24129),
            .in2(_gnd_net_),
            .in3(N__22480),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_8_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_8_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__24084),
            .in2(_gnd_net_),
            .in3(N__22465),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_8_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_8_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__24048),
            .in2(_gnd_net_),
            .in3(N__22453),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_8_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_8_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__24003),
            .in2(_gnd_net_),
            .in3(N__22438),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_8_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_8_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__23958),
            .in2(_gnd_net_),
            .in3(N__22423),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_8_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_8_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__23919),
            .in2(_gnd_net_),
            .in3(N__22405),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_8_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_8_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__24306),
            .in2(N__27296),
            .in3(N__22393),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_8_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_8_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_8_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__24277),
            .in2(_gnd_net_),
            .in3(N__22390),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29292),
            .ce(N__25078),
            .sr(N__28753));
    defparam \ppm_encoder_1.elevator_10_LC_8_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_8_21_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_8_21_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_8_21_6  (
            .in0(N__25888),
            .in1(N__24535),
            .in2(N__24960),
            .in3(N__22676),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29285),
            .ce(),
            .sr(N__28760));
    defparam \ppm_encoder_1.elevator_12_LC_8_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_8_22_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_8_22_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_8_22_1  (
            .in0(N__24520),
            .in1(N__26452),
            .in2(N__24959),
            .in3(N__22874),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29281),
            .ce(),
            .sr(N__28767));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_8_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_8_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_8_25_2  (
            .in0(N__22847),
            .in1(N__22717),
            .in2(_gnd_net_),
            .in3(N__22684),
            .lcout(\ppm_encoder_1.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_8_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_8_27_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_8_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_8_27_3  (
            .in0(N__23127),
            .in1(N__22651),
            .in2(_gnd_net_),
            .in3(N__22639),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29263),
            .ce(N__23062),
            .sr(N__28785));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_8_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_8_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_8_28_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_8_28_1  (
            .in0(N__23253),
            .in1(N__22631),
            .in2(N__23287),
            .in3(N__22610),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_8_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_8_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_8_28_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_8_28_2  (
            .in0(N__22589),
            .in1(N__22568),
            .in2(N__22549),
            .in3(N__23293),
            .lcout(\ppm_encoder_1.N_144_17 ),
            .ltout(\ppm_encoder_1.N_144_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_8_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_8_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_8_28_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_8_28_3  (
            .in0(N__22534),
            .in1(N__22525),
            .in2(N__22513),
            .in3(N__23385),
            .lcout(\ppm_encoder_1.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_8_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_8_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_8_28_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_8_28_4  (
            .in0(_gnd_net_),
            .in1(N__28930),
            .in2(_gnd_net_),
            .in3(N__23797),
            .lcout(\ppm_encoder_1.N_590_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_8_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_8_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_8_28_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_8_28_5  (
            .in0(_gnd_net_),
            .in1(N__22995),
            .in2(_gnd_net_),
            .in3(N__23312),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_8_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_8_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_8_29_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_8_29_0  (
            .in0(N__23200),
            .in1(N__23282),
            .in2(N__23266),
            .in3(N__23252),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_8_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_8_29_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_8_29_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_8_29_1  (
            .in0(N__23227),
            .in1(N__23137),
            .in2(_gnd_net_),
            .in3(N__23209),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29260),
            .ce(N__23056),
            .sr(N__28791));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_8_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_8_29_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_8_29_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_8_29_3  (
            .in0(N__23194),
            .in1(N__23135),
            .in2(_gnd_net_),
            .in3(N__23179),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29260),
            .ce(N__23056),
            .sr(N__28791));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_8_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_8_29_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_8_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_8_29_5  (
            .in0(N__23158),
            .in1(N__23146),
            .in2(_gnd_net_),
            .in3(N__23136),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29260),
            .ce(N__23056),
            .sr(N__28791));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_29_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_29_6  (
            .in0(N__23002),
            .in1(N__23402),
            .in2(N__23485),
            .in3(N__22994),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_16_LC_8_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_8_30_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_8_30_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_8_30_1  (
            .in0(N__22969),
            .in1(N__22938),
            .in2(N__23872),
            .in3(N__23827),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29258),
            .ce(),
            .sr(N__28795));
    defparam \ppm_encoder_1.pulses2count_17_LC_8_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_8_30_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_8_30_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_8_30_2  (
            .in0(N__23825),
            .in1(N__22924),
            .in2(N__22896),
            .in3(N__23870),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29258),
            .ce(),
            .sr(N__28795));
    defparam \ppm_encoder_1.pulses2count_15_LC_8_30_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_8_30_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_8_30_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_8_30_3  (
            .in0(N__23893),
            .in1(N__23484),
            .in2(N__23871),
            .in3(N__23826),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29258),
            .ce(),
            .sr(N__28795));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_30_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_30_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_30_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_8_30_6  (
            .in0(N__23468),
            .in1(N__23447),
            .in2(N__23428),
            .in3(N__23403),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_1 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23365),
            .lcout(\uart_pc_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29389),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23359),
            .lcout(\uart_pc_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29389),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_9_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_9_10_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_9_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset2data_ess_7_LC_9_10_7  (
            .in0(N__27649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29362),
            .ce(N__24617),
            .sr(N__28713));
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_9_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29860),
            .lcout(frame_decoder_OFF2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29349),
            .ce(N__24624),
            .sr(N__28718));
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_9_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_1_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27774),
            .lcout(frame_decoder_OFF2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29349),
            .ce(N__24624),
            .sr(N__28718));
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_9_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_4_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27993),
            .lcout(frame_decoder_OFF2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29349),
            .ce(N__24624),
            .sr(N__28718));
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_9_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_9_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_2_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28361),
            .lcout(frame_decoder_OFF2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29349),
            .ce(N__24624),
            .sr(N__28718));
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_9_13_0 .C_ON=1'b1;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__25261),
            .in2(N__25165),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_6_LC_9_13_1 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_6_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_6_LC_9_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_6_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__24138),
            .in2(N__25271),
            .in3(N__24145),
            .lcout(scaler_2_data_6),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_1 ),
            .carryout(\scaler_2.un2_source_data_0_cry_2 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_7_LC_9_13_2 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_7_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_7_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_7_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(N__24142),
            .in3(N__24106),
            .lcout(scaler_2_data_7),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_2 ),
            .carryout(\scaler_2.un2_source_data_0_cry_3 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_8_LC_9_13_3 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_8_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_8_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_8_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__24060),
            .in2(N__24103),
            .in3(N__24067),
            .lcout(scaler_2_data_8),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_3 ),
            .carryout(\scaler_2.un2_source_data_0_cry_4 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_9_LC_9_13_4 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_9_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_9_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_9_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__24018),
            .in2(N__24064),
            .in3(N__24025),
            .lcout(scaler_2_data_9),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_4 ),
            .carryout(\scaler_2.un2_source_data_0_cry_5 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_10_LC_9_13_5 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_10_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_10_LC_9_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_10_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__23973),
            .in2(N__24022),
            .in3(N__23980),
            .lcout(scaler_2_data_10),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_5 ),
            .carryout(\scaler_2.un2_source_data_0_cry_6 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_11_LC_9_13_6 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_11_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_11_LC_9_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_11_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__23934),
            .in2(N__23977),
            .in3(N__23941),
            .lcout(scaler_2_data_11),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_6 ),
            .carryout(\scaler_2.un2_source_data_0_cry_7 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_12_LC_9_13_7 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_12_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_12_LC_9_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_12_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__24327),
            .in2(N__23938),
            .in3(N__23896),
            .lcout(scaler_2_data_12),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_7 ),
            .carryout(\scaler_2.un2_source_data_0_cry_8 ),
            .clk(N__29344),
            .ce(N__26374),
            .sr(N__28723));
    defparam \scaler_2.source_data_1_esr_13_LC_9_14_0 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_13_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_13_LC_9_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_13_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__24328),
            .in2(N__24316),
            .in3(N__24283),
            .lcout(scaler_2_data_13),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_9 ),
            .clk(N__29338),
            .ce(N__26377),
            .sr(N__28726));
    defparam \scaler_2.source_data_1_esr_14_LC_9_14_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_14_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_14_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_2.source_data_1_esr_14_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24280),
            .lcout(scaler_2_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29338),
            .ce(N__26377),
            .sr(N__28726));
    defparam \scaler_2.source_data_1_esr_5_LC_9_15_0 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_5_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_5_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.source_data_1_esr_5_LC_9_15_0  (
            .in0(N__25242),
            .in1(N__25276),
            .in2(_gnd_net_),
            .in3(N__25210),
            .lcout(scaler_2_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29330),
            .ce(N__26380),
            .sr(N__28731));
    defparam \scaler_3.source_data_1_esr_5_LC_9_15_2 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_5_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_5_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.source_data_1_esr_5_LC_9_15_2  (
            .in0(N__27517),
            .in1(N__29734),
            .in2(_gnd_net_),
            .in3(N__27490),
            .lcout(scaler_3_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29330),
            .ce(N__26380),
            .sr(N__28731));
    defparam \scaler_4.source_data_1_esr_5_LC_9_15_4 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_9_15_4  (
            .in0(N__25818),
            .in1(N__25852),
            .in2(_gnd_net_),
            .in3(N__26812),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29330),
            .ce(N__26380),
            .sr(N__28731));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_15_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_15_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_9_15_6  (
            .in0(N__26264),
            .in1(N__26335),
            .in2(_gnd_net_),
            .in3(N__26094),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_9_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_9_16_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_9_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_9_16_2  (
            .in0(N__29657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27374),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29321),
            .ce(),
            .sr(N__28736));
    defparam \scaler_2.source_data_1_4_LC_9_16_4 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_4_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_4_LC_9_16_4 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_2.source_data_1_4_LC_9_16_4  (
            .in0(N__27347),
            .in1(N__25243),
            .in2(N__24198),
            .in3(N__25209),
            .lcout(scaler_2_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29321),
            .ce(),
            .sr(N__28736));
    defparam \scaler_3.source_data_1_4_LC_9_16_5 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_4_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_4_LC_9_16_5 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_3.source_data_1_4_LC_9_16_5  (
            .in0(N__27349),
            .in1(N__29730),
            .in2(N__24498),
            .in3(N__27489),
            .lcout(scaler_3_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29321),
            .ce(),
            .sr(N__28736));
    defparam \scaler_4.source_data_1_4_LC_9_16_6 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_9_16_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_9_16_6  (
            .in0(N__27348),
            .in1(N__25860),
            .in2(N__24468),
            .in3(N__26811),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29321),
            .ce(),
            .sr(N__28736));
    defparam \Commands_frame_decoder.state_1_RNI2D06_1_LC_9_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI2D06_1_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI2D06_1_LC_9_17_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_1_RNI2D06_1_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__26183),
            .in2(_gnd_net_),
            .in3(N__24343),
            .lcout(\Commands_frame_decoder.N_282_0 ),
            .ltout(\Commands_frame_decoder.N_282_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_2_0_LC_9_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_2_0_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_2_0_LC_9_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_2_0_LC_9_17_1  (
            .in0(N__28309),
            .in1(N__27852),
            .in2(N__24451),
            .in3(N__24447),
            .lcout(\Commands_frame_decoder.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_3_0_LC_9_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_3_0_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_3_0_LC_9_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_3_0_LC_9_17_3  (
            .in0(N__29847),
            .in1(N__28311),
            .in2(N__24353),
            .in3(N__24433),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNO_0_0_LC_9_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNO_0_0_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNO_0_0_LC_9_17_4 .LUT_INIT=16'b0001000100010101;
    LogicCell40 \Commands_frame_decoder.state_1_RNO_0_0_LC_9_17_4  (
            .in0(N__26163),
            .in1(N__24381),
            .in2(N__24418),
            .in3(N__24415),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_1_ns_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_0_LC_9_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_0_LC_9_17_5 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_1_0_LC_9_17_5 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \Commands_frame_decoder.state_1_0_LC_9_17_5  (
            .in0(N__24409),
            .in1(N__24403),
            .in2(N__24397),
            .in3(N__29461),
            .lcout(\Commands_frame_decoder.state_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29310),
            .ce(),
            .sr(N__28741));
    defparam \Commands_frame_decoder.state_1_10_LC_9_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_10_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_10_LC_9_17_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Commands_frame_decoder.state_1_10_LC_9_17_6  (
            .in0(N__29462),
            .in1(N__29698),
            .in2(N__26167),
            .in3(N__26184),
            .lcout(\Commands_frame_decoder.state_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29310),
            .ce(),
            .sr(N__28741));
    defparam \Commands_frame_decoder.state_1_1_LC_9_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_1_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_1_LC_9_17_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_1_1_LC_9_17_7  (
            .in0(N__24382),
            .in1(N__24367),
            .in2(N__24354),
            .in3(N__29460),
            .lcout(\Commands_frame_decoder.state_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29310),
            .ce(),
            .sr(N__28741));
    defparam \uart_drone.bit_Count_2_LC_9_18_3 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_9_18_3 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uart_drone.bit_Count_2_LC_9_18_3  (
            .in0(N__25489),
            .in1(N__26737),
            .in2(N__26336),
            .in3(N__26253),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29302),
            .ce(),
            .sr(N__28747));
    defparam \uart_drone.bit_Count_1_LC_9_18_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_9_18_6 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uart_drone.bit_Count_1_LC_9_18_6  (
            .in0(N__26252),
            .in1(N__25488),
            .in2(N__26149),
            .in3(N__26090),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29302),
            .ce(),
            .sr(N__28747));
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_9_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__25986),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_9_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25959),
            .in2(_gnd_net_),
            .in3(N__24571),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_9_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_9_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__25935),
            .in2(_gnd_net_),
            .in3(N__24556),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_9_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25911),
            .in2(_gnd_net_),
            .in3(N__24538),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_9_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_9_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__25887),
            .in2(_gnd_net_),
            .in3(N__24526),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_9_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_9_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__26478),
            .in2(_gnd_net_),
            .in3(N__24523),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_9_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_9_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__26451),
            .in2(_gnd_net_),
            .in3(N__24511),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_9_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_9_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__26421),
            .in2(N__27297),
            .in3(N__25105),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_9_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_9_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__26392),
            .in2(_gnd_net_),
            .in3(N__25102),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29286),
            .ce(N__25077),
            .sr(N__28761));
    defparam \ppm_encoder_1.elevator_13_LC_9_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_9_22_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_9_22_1 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_9_22_1  (
            .in0(N__26425),
            .in1(N__25015),
            .in2(N__25001),
            .in3(N__24913),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29274),
            .ce(),
            .sr(N__28773));
    defparam \ppm_encoder_1.elevator_11_LC_9_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_9_24_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_9_24_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_9_24_0  (
            .in0(N__26479),
            .in1(N__24976),
            .in2(N__24961),
            .in3(N__24674),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29266),
            .ce(),
            .sr(N__28779));
    defparam \Commands_frame_decoder.state_1_RNITK1O_4_LC_10_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNITK1O_4_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNITK1O_4_LC_10_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_1_RNITK1O_4_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__24651),
            .in2(_gnd_net_),
            .in3(N__28934),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_12_1 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27648),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29339),
            .ce(N__26773),
            .sr(N__28719));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_10_13_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_10_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__25155),
            .in2(_gnd_net_),
            .in3(N__24633),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_545_i_l_ofx_LC_10_13_3 .C_ON=1'b0;
    defparam \scaler_4.N_545_i_l_ofx_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_545_i_l_ofx_LC_10_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_545_i_l_ofx_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__25156),
            .in2(_gnd_net_),
            .in3(N__24634),
            .lcout(\scaler_4.N_545_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI0O1O_7_LC_10_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI0O1O_7_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI0O1O_7_LC_10_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_1_RNI0O1O_7_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__29505),
            .in2(_gnd_net_),
            .in3(N__28927),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_10_13_7 .C_ON=1'b0;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_10_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_10_13_7  (
            .in0(N__25275),
            .in1(N__25234),
            .in2(_gnd_net_),
            .in3(N__25208),
            .lcout(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_10_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28356),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28001),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_10_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_10_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29856),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_10_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27870),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_10_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27768),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_14_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_10_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27639),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29323),
            .ce(N__29683),
            .sr(N__28727));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_10_15_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_10_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__25802),
            .in2(N__25147),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_10_15_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__25767),
            .in2(N__25811),
            .in3(N__25108),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_7_LC_10_15_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__25746),
            .in2(N__25771),
            .in3(N__25444),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_8_LC_10_15_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__25713),
            .in2(N__25750),
            .in3(N__25420),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_9_LC_10_15_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__25683),
            .in2(N__25717),
            .in3(N__25396),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_10_LC_10_15_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__25659),
            .in2(N__25687),
            .in3(N__25372),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_11_LC_10_15_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__25638),
            .in2(N__25663),
            .in3(N__25348),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_12_LC_10_15_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__26022),
            .in2(N__25642),
            .in3(N__25324),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__29312),
            .ce(N__26375),
            .sr(N__28732));
    defparam \scaler_4.source_data_1_esr_13_LC_10_16_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__26023),
            .in2(N__26005),
            .in3(N__25297),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__29304),
            .ce(N__26378),
            .sr(N__28737));
    defparam \scaler_4.source_data_1_esr_14_LC_10_16_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25294),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29304),
            .ce(N__26378),
            .sr(N__28737));
    defparam \uart_drone.bit_Count_0_LC_10_17_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_10_17_2 .LUT_INIT=16'b0100010001100100;
    LogicCell40 \uart_drone.bit_Count_0_LC_10_17_2  (
            .in0(N__26148),
            .in1(N__26108),
            .in2(N__25588),
            .in3(N__25524),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29293),
            .ce(),
            .sr(N__28742));
    defparam \Commands_frame_decoder.state_1_7_LC_10_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_7_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_7_LC_10_17_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_1_7_LC_10_17_6  (
            .in0(N__25480),
            .in1(N__29649),
            .in2(N__25627),
            .in3(N__29463),
            .lcout(\Commands_frame_decoder.state_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29293),
            .ce(),
            .sr(N__28742));
    defparam \uart_drone.state_RNI63LK2_3_LC_10_18_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_18_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_10_18_6  (
            .in0(N__25587),
            .in1(N__26137),
            .in2(_gnd_net_),
            .in3(N__25523),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI3BRE_7_LC_10_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI3BRE_7_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI3BRE_7_LC_10_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI3BRE_7_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__25479),
            .in2(_gnd_net_),
            .in3(N__29648),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_11_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29849),
            .lcout(frame_decoder_CH3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29331),
            .ce(N__27404),
            .sr(N__28724));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_11_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28353),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29324),
            .ce(N__26774),
            .sr(N__28728));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_11_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28115),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29324),
            .ce(N__26774),
            .sr(N__28728));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_11_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29324),
            .ce(N__26774),
            .sr(N__28728));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_11_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27890),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29324),
            .ce(N__26774),
            .sr(N__28728));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_11_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28231),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29324),
            .ce(N__26774),
            .sr(N__28728));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_14_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__26793),
            .in2(N__25856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_14_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__25825),
            .in2(N__26824),
            .in3(N__25789),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_14_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__25786),
            .in2(N__25780),
            .in3(N__25759),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_14_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__25756),
            .in2(N__28387),
            .in3(N__25738),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_14_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__25735),
            .in2(N__25729),
            .in3(N__25705),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_14_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__25702),
            .in2(N__25696),
            .in3(N__25675),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_14_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__25672),
            .in2(N__28375),
            .in3(N__25651),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_14_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__25648),
            .in2(_gnd_net_),
            .in3(N__25630),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_15_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__26032),
            .in2(N__27307),
            .in3(N__26011),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_15_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26008),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_16_0 .C_ON=1'b1;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__27508),
            .in2(N__27454),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.source_data_1_esr_6_LC_11_16_1 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_6_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_6_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_6_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__26973),
            .in2(N__27516),
            .in3(N__25969),
            .lcout(scaler_3_data_6),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_1 ),
            .carryout(\scaler_3.un2_source_data_0_cry_2 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_7_LC_11_16_2 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_7_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_7_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_7_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__26952),
            .in2(N__26977),
            .in3(N__25942),
            .lcout(scaler_3_data_7),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_2 ),
            .carryout(\scaler_3.un2_source_data_0_cry_3 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_8_LC_11_16_3 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_8_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_8_LC_11_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_8_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__26931),
            .in2(N__26956),
            .in3(N__25918),
            .lcout(scaler_3_data_8),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_3 ),
            .carryout(\scaler_3.un2_source_data_0_cry_4 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_9_LC_11_16_4 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_9_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_9_LC_11_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_9_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__26907),
            .in2(N__26935),
            .in3(N__25891),
            .lcout(scaler_3_data_9),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_4 ),
            .carryout(\scaler_3.un2_source_data_0_cry_5 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_10_LC_11_16_5 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_10_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_10_LC_11_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_10_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__26886),
            .in2(N__26911),
            .in3(N__25864),
            .lcout(scaler_3_data_10),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_5 ),
            .carryout(\scaler_3.un2_source_data_0_cry_6 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_11_LC_11_16_6 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_11_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_11_LC_11_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_11_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__26871),
            .in2(N__26890),
            .in3(N__26455),
            .lcout(scaler_3_data_11),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_6 ),
            .carryout(\scaler_3.un2_source_data_0_cry_7 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_12_LC_11_16_7 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_12_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_12_LC_11_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_12_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__26859),
            .in2(N__26875),
            .in3(N__26428),
            .lcout(scaler_3_data_12),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_7 ),
            .carryout(\scaler_3.un2_source_data_0_cry_8 ),
            .clk(N__29294),
            .ce(N__26376),
            .sr(N__28743));
    defparam \scaler_3.source_data_1_esr_13_LC_11_17_0 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_13_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_13_LC_11_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_13_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__26860),
            .in2(N__26842),
            .in3(N__26398),
            .lcout(scaler_3_data_13),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_9 ),
            .clk(N__29287),
            .ce(N__26379),
            .sr(N__28748));
    defparam \scaler_3.source_data_1_esr_14_LC_11_17_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_14_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_14_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_3.source_data_1_esr_14_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26395),
            .lcout(scaler_3_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29287),
            .ce(N__26379),
            .sr(N__28748));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_18_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_18_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_11_18_0  (
            .in0(N__26073),
            .in1(N__26334),
            .in2(_gnd_net_),
            .in3(N__26263),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_11_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_11_18_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_11_18_2  (
            .in0(N__26194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26713),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNIDIPF_10_LC_11_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNIDIPF_10_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNIDIPF_10_LC_11_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNIDIPF_10_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__29647),
            .in2(_gnd_net_),
            .in3(N__26193),
            .lcout(\Commands_frame_decoder.state_1_ns_i_a4_2_0_0 ),
            .ltout(\Commands_frame_decoder.state_1_ns_i_a4_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNI0PVH1_2_LC_11_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNI0PVH1_2_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNI0PVH1_2_LC_11_18_4 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Commands_frame_decoder.count_RNI0PVH1_2_LC_11_18_4  (
            .in0(N__26521),
            .in1(N__26497),
            .in2(N__26170),
            .in3(N__27003),
            .lcout(\Commands_frame_decoder.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_11_18_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_11_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__26147),
            .in2(_gnd_net_),
            .in3(N__26072),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count8_cry_0_c_LC_11_19_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.count8_cry_0_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_cry_0_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Commands_frame_decoder.count8_cry_0_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__27042),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\Commands_frame_decoder.count8_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count8_cry_1_c_inv_LC_11_19_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.count8_cry_1_c_inv_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_cry_1_c_inv_LC_11_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Commands_frame_decoder.count8_cry_1_c_inv_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__26728),
            .in2(_gnd_net_),
            .in3(N__26494),
            .lcout(\Commands_frame_decoder.count8_axb_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.count8_cry_0 ),
            .carryout(\Commands_frame_decoder.count8_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count8_cry_2_c_inv_LC_11_19_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.count8_cry_2_c_inv_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_cry_2_c_inv_LC_11_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Commands_frame_decoder.count8_cry_2_c_inv_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__26722),
            .in2(N__27299),
            .in3(N__26519),
            .lcout(\Commands_frame_decoder.count_i_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.count8_cry_1 ),
            .carryout(\Commands_frame_decoder.count8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count8_THRU_LUT4_0_LC_11_19_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count8_THRU_LUT4_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_THRU_LUT4_0_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.count8_THRU_LUT4_0_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26716),
            .lcout(\Commands_frame_decoder.count8_THRU_CO ),
            .ltout(\Commands_frame_decoder.count8_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count8_cry_2_c_RNIARGV_LC_11_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count8_cry_2_c_RNIARGV_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_cry_2_c_RNIARGV_LC_11_19_4 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \Commands_frame_decoder.count8_cry_2_c_RNIARGV_LC_11_19_4  (
            .in0(N__26657),
            .in1(_gnd_net_),
            .in2(N__26527),
            .in3(N__27018),
            .lcout(\Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0 ),
            .ltout(\Commands_frame_decoder.count8_cry_2_c_RNIARGVZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_2_LC_11_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_2_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_2_LC_11_19_5 .LUT_INIT=16'b0110000010100000;
    LogicCell40 \Commands_frame_decoder.count_2_LC_11_19_5  (
            .in0(N__26520),
            .in1(N__26506),
            .in2(N__26524),
            .in3(N__26496),
            .lcout(\Commands_frame_decoder.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29276),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIT86R_0_LC_11_19_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIT86R_0_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIT86R_0_LC_11_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.count_RNIT86R_0_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__27017),
            .in2(_gnd_net_),
            .in3(N__27004),
            .lcout(\Commands_frame_decoder.CO0 ),
            .ltout(\Commands_frame_decoder.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_1_LC_11_19_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_1_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_1_LC_11_19_7 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \Commands_frame_decoder.count_1_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__27030),
            .in2(N__26500),
            .in3(N__26495),
            .lcout(\Commands_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29276),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_12_3_3 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_12_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_2.source_data_1_esr_ctle_14_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__27346),
            .in2(_gnd_net_),
            .in3(N__28924),
            .lcout(pc_frame_decoder_dv_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_12_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27775),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29322),
            .ce(N__26782),
            .sr(N__28729));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_12_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29848),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29311),
            .ce(N__26781),
            .sr(N__28733));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28002),
            .lcout(frame_decoder_CH3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29303),
            .ce(N__27417),
            .sr(N__28738));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28360),
            .lcout(frame_decoder_CH3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29303),
            .ce(N__27417),
            .sr(N__28738));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28106),
            .lcout(frame_decoder_CH3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29303),
            .ce(N__27417),
            .sr(N__28738));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27891),
            .lcout(frame_decoder_CH3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29303),
            .ce(N__27417),
            .sr(N__28738));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28228),
            .lcout(frame_decoder_CH3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29303),
            .ce(N__27417),
            .sr(N__28738));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_12_15_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__27487),
            .in2(N__29729),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_12_15_1 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__27439),
            .in2(N__27658),
            .in3(N__26740),
            .lcout(\scaler_3.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_0 ),
            .carryout(\scaler_3.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_12_15_2 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__26983),
            .in2(N__28240),
            .in3(N__26965),
            .lcout(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_1 ),
            .carryout(\scaler_3.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_12_15_3 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__26962),
            .in2(N__28012),
            .in3(N__26944),
            .lcout(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_2 ),
            .carryout(\scaler_3.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_12_15_4 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__26941),
            .in2(N__27901),
            .in3(N__26923),
            .lcout(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_3 ),
            .carryout(\scaler_3.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_12_15_5 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__27781),
            .in2(N__26920),
            .in3(N__26899),
            .lcout(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_4 ),
            .carryout(\scaler_3.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_12_15_6 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__26896),
            .in2(N__28126),
            .in3(N__26878),
            .lcout(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_5 ),
            .carryout(\scaler_3.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_12_15_7 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_12_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__27445),
            .in2(_gnd_net_),
            .in3(N__26863),
            .lcout(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_6 ),
            .carryout(\scaler_3.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_12_16_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__27523),
            .in2(N__27306),
            .in3(N__26848),
            .lcout(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_12_16_1 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26845),
            .lcout(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.N_533_i_l_ofx_LC_12_16_2 .C_ON=1'b0;
    defparam \scaler_3.N_533_i_l_ofx_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.N_533_i_l_ofx_LC_12_16_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \scaler_3.N_533_i_l_ofx_LC_12_16_2  (
            .in0(N__27430),
            .in1(_gnd_net_),
            .in2(N__27535),
            .in3(_gnd_net_),
            .lcout(\scaler_3.N_533_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_12_16_3 .C_ON=1'b0;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_12_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_12_16_3  (
            .in0(N__27515),
            .in1(N__29722),
            .in2(_gnd_net_),
            .in3(N__27488),
            .lcout(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_12_16_5 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_12_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__27531),
            .in2(_gnd_net_),
            .in3(N__27429),
            .lcout(\scaler_3.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27763),
            .lcout(frame_decoder_CH3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29282),
            .ce(N__27421),
            .sr(N__28754));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_17_3 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27605),
            .lcout(frame_decoder_CH3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29282),
            .ce(N__27421),
            .sr(N__28754));
    defparam \Commands_frame_decoder.source_data_valid_LC_12_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_12_18_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_12_18_7  (
            .in0(N__27387),
            .in1(N__29658),
            .in2(N__27337),
            .in3(N__27355),
            .lcout(pc_frame_decoder_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29275),
            .ce(),
            .sr(N__28762));
    defparam \Commands_frame_decoder.count8_cry_0_c_inv_LC_12_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count8_cry_0_c_inv_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count8_cry_0_c_inv_LC_12_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Commands_frame_decoder.count8_cry_0_c_inv_LC_12_19_0  (
            .in0(N__27043),
            .in1(N__27298),
            .in2(_gnd_net_),
            .in3(N__27001),
            .lcout(\Commands_frame_decoder.count8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_12_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_12_19_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_12_19_4  (
            .in0(N__27031),
            .in1(N__27019),
            .in2(_gnd_net_),
            .in3(N__27002),
            .lcout(\Commands_frame_decoder.count8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29269),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_13_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_13_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_13_14_1  (
            .in0(N__28117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29313),
            .ce(N__29682),
            .sr(N__28744));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_13_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_13_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_13_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28229),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29313),
            .ce(N__29682),
            .sr(N__28744));
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_13_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_13_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_2_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28363),
            .lcout(frame_decoder_OFF3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_13_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_13_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_6_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28194),
            .lcout(frame_decoder_OFF3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_13_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_13_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_3_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28116),
            .lcout(frame_decoder_OFF3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_13_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_13_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_4_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28003),
            .lcout(frame_decoder_OFF3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_13_15_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_13_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_5_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27892),
            .lcout(frame_decoder_OFF3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_13_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_1_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27770),
            .lcout(frame_decoder_OFF3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29305),
            .ce(N__29527),
            .sr(N__28749));
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_13_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_13_16_5 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_13_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_ess_7_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27646),
            .lcout(frame_decoder_OFF3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29295),
            .ce(N__29523),
            .sr(N__28755));
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_13_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_13_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_0_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29839),
            .lcout(frame_decoder_OFF3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29295),
            .ce(N__29523),
            .sr(N__28755));
    defparam \Commands_frame_decoder.state_1_RNI5DRE_9_LC_13_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI5DRE_9_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI5DRE_9_LC_13_17_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI5DRE_9_LC_13_17_4  (
            .in0(N__29403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29656),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI2Q1O_9_LC_13_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI2Q1O_9_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI2Q1O_9_LC_13_17_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI2Q1O_9_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29686),
            .in3(N__28937),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI4CRE_8_LC_14_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI4CRE_8_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI4CRE_8_LC_14_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI4CRE_8_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__29481),
            .in2(_gnd_net_),
            .in3(N__29659),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_RNI1P1O_8_LC_14_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_RNI1P1O_8_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_1_RNI1P1O_8_LC_14_16_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_1_RNI1P1O_8_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29530),
            .in3(N__28939),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_8_LC_14_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_8_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_8_LC_14_17_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_1_8_LC_14_17_3  (
            .in0(N__29482),
            .in1(N__29506),
            .in2(_gnd_net_),
            .in3(N__29469),
            .lcout(\Commands_frame_decoder.state_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29296),
            .ce(),
            .sr(N__28768));
    defparam \Commands_frame_decoder.state_1_9_LC_14_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_9_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_9_LC_14_17_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_1_9_LC_14_17_6  (
            .in0(N__29470),
            .in1(N__29410),
            .in2(_gnd_net_),
            .in3(N__29404),
            .lcout(\Commands_frame_decoder.state_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29296),
            .ce(),
            .sr(N__28768));
endmodule // Pc2drone
