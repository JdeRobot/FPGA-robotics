// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Apr 14 2019 14:18:13

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__37457;
    wire N__37456;
    wire N__37455;
    wire N__37446;
    wire N__37445;
    wire N__37444;
    wire N__37437;
    wire N__37436;
    wire N__37435;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37410;
    wire N__37409;
    wire N__37408;
    wire N__37401;
    wire N__37400;
    wire N__37399;
    wire N__37392;
    wire N__37391;
    wire N__37390;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37374;
    wire N__37373;
    wire N__37372;
    wire N__37365;
    wire N__37364;
    wire N__37363;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37327;
    wire N__37326;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37299;
    wire N__37296;
    wire N__37289;
    wire N__37288;
    wire N__37287;
    wire N__37286;
    wire N__37283;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37251;
    wire N__37248;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37236;
    wire N__37233;
    wire N__37228;
    wire N__37227;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37212;
    wire N__37209;
    wire N__37204;
    wire N__37193;
    wire N__37192;
    wire N__37191;
    wire N__37190;
    wire N__37189;
    wire N__37186;
    wire N__37185;
    wire N__37176;
    wire N__37175;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37161;
    wire N__37158;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37133;
    wire N__37132;
    wire N__37131;
    wire N__37128;
    wire N__37127;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37119;
    wire N__37118;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37108;
    wire N__37107;
    wire N__37106;
    wire N__37097;
    wire N__37094;
    wire N__37087;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37064;
    wire N__37063;
    wire N__37062;
    wire N__37061;
    wire N__37052;
    wire N__37051;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37041;
    wire N__37038;
    wire N__37033;
    wire N__37030;
    wire N__37029;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36969;
    wire N__36966;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36929;
    wire N__36926;
    wire N__36921;
    wire N__36914;
    wire N__36913;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36901;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36894;
    wire N__36893;
    wire N__36892;
    wire N__36891;
    wire N__36890;
    wire N__36889;
    wire N__36888;
    wire N__36887;
    wire N__36886;
    wire N__36885;
    wire N__36884;
    wire N__36883;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36851;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36774;
    wire N__36773;
    wire N__36772;
    wire N__36771;
    wire N__36770;
    wire N__36769;
    wire N__36768;
    wire N__36767;
    wire N__36766;
    wire N__36765;
    wire N__36764;
    wire N__36763;
    wire N__36762;
    wire N__36761;
    wire N__36760;
    wire N__36759;
    wire N__36758;
    wire N__36757;
    wire N__36756;
    wire N__36755;
    wire N__36754;
    wire N__36753;
    wire N__36752;
    wire N__36751;
    wire N__36750;
    wire N__36749;
    wire N__36748;
    wire N__36747;
    wire N__36746;
    wire N__36745;
    wire N__36744;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36740;
    wire N__36739;
    wire N__36738;
    wire N__36737;
    wire N__36736;
    wire N__36735;
    wire N__36734;
    wire N__36733;
    wire N__36732;
    wire N__36731;
    wire N__36730;
    wire N__36729;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36717;
    wire N__36716;
    wire N__36715;
    wire N__36714;
    wire N__36713;
    wire N__36712;
    wire N__36711;
    wire N__36710;
    wire N__36709;
    wire N__36708;
    wire N__36707;
    wire N__36706;
    wire N__36705;
    wire N__36704;
    wire N__36703;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36352;
    wire N__36351;
    wire N__36346;
    wire N__36345;
    wire N__36344;
    wire N__36343;
    wire N__36340;
    wire N__36339;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36328;
    wire N__36327;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36303;
    wire N__36294;
    wire N__36291;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36270;
    wire N__36263;
    wire N__36260;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36218;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36208;
    wire N__36201;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36167;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36163;
    wire N__36162;
    wire N__36161;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36157;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36153;
    wire N__36152;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36142;
    wire N__36141;
    wire N__36140;
    wire N__36139;
    wire N__36138;
    wire N__36137;
    wire N__36136;
    wire N__36135;
    wire N__36134;
    wire N__36133;
    wire N__36132;
    wire N__36131;
    wire N__36130;
    wire N__36129;
    wire N__36128;
    wire N__36127;
    wire N__36126;
    wire N__36125;
    wire N__36124;
    wire N__36123;
    wire N__36122;
    wire N__36121;
    wire N__36120;
    wire N__36119;
    wire N__36118;
    wire N__36117;
    wire N__36116;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36112;
    wire N__36111;
    wire N__36110;
    wire N__36109;
    wire N__36108;
    wire N__36107;
    wire N__36106;
    wire N__36105;
    wire N__36104;
    wire N__36103;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36098;
    wire N__36097;
    wire N__36096;
    wire N__36095;
    wire N__36094;
    wire N__36093;
    wire N__36092;
    wire N__36091;
    wire N__36090;
    wire N__36089;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36081;
    wire N__36080;
    wire N__36079;
    wire N__36078;
    wire N__36077;
    wire N__36076;
    wire N__36075;
    wire N__36074;
    wire N__36073;
    wire N__36072;
    wire N__36071;
    wire N__36070;
    wire N__36069;
    wire N__36068;
    wire N__36067;
    wire N__36066;
    wire N__36065;
    wire N__36064;
    wire N__36063;
    wire N__36062;
    wire N__36061;
    wire N__36060;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36056;
    wire N__36055;
    wire N__36054;
    wire N__36053;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36048;
    wire N__36047;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36043;
    wire N__36042;
    wire N__36041;
    wire N__36040;
    wire N__36039;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36035;
    wire N__36034;
    wire N__36033;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36027;
    wire N__36026;
    wire N__36025;
    wire N__36024;
    wire N__36023;
    wire N__36022;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35683;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35652;
    wire N__35645;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35630;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35582;
    wire N__35575;
    wire N__35572;
    wire N__35567;
    wire N__35566;
    wire N__35565;
    wire N__35560;
    wire N__35557;
    wire N__35552;
    wire N__35549;
    wire N__35548;
    wire N__35547;
    wire N__35544;
    wire N__35539;
    wire N__35534;
    wire N__35533;
    wire N__35532;
    wire N__35529;
    wire N__35524;
    wire N__35519;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35507;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35495;
    wire N__35492;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35480;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35468;
    wire N__35465;
    wire N__35464;
    wire N__35463;
    wire N__35462;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35441;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35429;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35417;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35337;
    wire N__35332;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35319;
    wire N__35314;
    wire N__35309;
    wire N__35306;
    wire N__35297;
    wire N__35294;
    wire N__35293;
    wire N__35292;
    wire N__35289;
    wire N__35284;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35269;
    wire N__35268;
    wire N__35265;
    wire N__35264;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35246;
    wire N__35241;
    wire N__35240;
    wire N__35237;
    wire N__35236;
    wire N__35233;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35217;
    wire N__35214;
    wire N__35209;
    wire N__35206;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35179;
    wire N__35176;
    wire N__35171;
    wire N__35168;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35156;
    wire N__35155;
    wire N__35154;
    wire N__35153;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35145;
    wire N__35140;
    wire N__35135;
    wire N__35130;
    wire N__35127;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35115;
    wire N__35114;
    wire N__35109;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35091;
    wire N__35084;
    wire N__35081;
    wire N__35080;
    wire N__35079;
    wire N__35078;
    wire N__35077;
    wire N__35076;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35064;
    wire N__35063;
    wire N__35060;
    wire N__35059;
    wire N__35058;
    wire N__35057;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35035;
    wire N__35034;
    wire N__35033;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35025;
    wire N__35024;
    wire N__35023;
    wire N__35022;
    wire N__35021;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__34999;
    wire N__34994;
    wire N__34991;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34902;
    wire N__34899;
    wire N__34894;
    wire N__34887;
    wire N__34884;
    wire N__34879;
    wire N__34874;
    wire N__34869;
    wire N__34866;
    wire N__34861;
    wire N__34850;
    wire N__34849;
    wire N__34848;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34833;
    wire N__34826;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34814;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34802;
    wire N__34799;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34784;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34760;
    wire N__34757;
    wire N__34756;
    wire N__34753;
    wire N__34752;
    wire N__34751;
    wire N__34748;
    wire N__34747;
    wire N__34746;
    wire N__34743;
    wire N__34738;
    wire N__34733;
    wire N__34730;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34625;
    wire N__34622;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34533;
    wire N__34530;
    wire N__34525;
    wire N__34518;
    wire N__34505;
    wire N__34504;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34481;
    wire N__34480;
    wire N__34475;
    wire N__34472;
    wire N__34471;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34449;
    wire N__34448;
    wire N__34443;
    wire N__34440;
    wire N__34435;
    wire N__34430;
    wire N__34427;
    wire N__34422;
    wire N__34409;
    wire N__34406;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34379;
    wire N__34378;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34364;
    wire N__34363;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34352;
    wire N__34339;
    wire N__34336;
    wire N__34335;
    wire N__34332;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34324;
    wire N__34323;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34287;
    wire N__34274;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34268;
    wire N__34267;
    wire N__34266;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34245;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34202;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34166;
    wire N__34165;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34161;
    wire N__34160;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34144;
    wire N__34137;
    wire N__34134;
    wire N__34133;
    wire N__34132;
    wire N__34131;
    wire N__34130;
    wire N__34129;
    wire N__34124;
    wire N__34121;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34091;
    wire N__34088;
    wire N__34083;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34042;
    wire N__34041;
    wire N__34040;
    wire N__34037;
    wire N__34032;
    wire N__34029;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34015;
    wire N__34012;
    wire N__34011;
    wire N__34010;
    wire N__34007;
    wire N__34000;
    wire N__33995;
    wire N__33992;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33956;
    wire N__33955;
    wire N__33954;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33918;
    wire N__33911;
    wire N__33908;
    wire N__33907;
    wire N__33906;
    wire N__33905;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33898;
    wire N__33893;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33874;
    wire N__33871;
    wire N__33860;
    wire N__33859;
    wire N__33858;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33836;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33826;
    wire N__33825;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33813;
    wire N__33812;
    wire N__33811;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33799;
    wire N__33792;
    wire N__33787;
    wire N__33776;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33764;
    wire N__33761;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33749;
    wire N__33746;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33734;
    wire N__33731;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33701;
    wire N__33698;
    wire N__33697;
    wire N__33696;
    wire N__33693;
    wire N__33688;
    wire N__33683;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33670;
    wire N__33665;
    wire N__33662;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33647;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33641;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33631;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33625;
    wire N__33624;
    wire N__33623;
    wire N__33622;
    wire N__33621;
    wire N__33618;
    wire N__33617;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33592;
    wire N__33589;
    wire N__33580;
    wire N__33577;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33563;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33538;
    wire N__33535;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33519;
    wire N__33514;
    wire N__33507;
    wire N__33494;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33485;
    wire N__33482;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33449;
    wire N__33448;
    wire N__33447;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33433;
    wire N__33428;
    wire N__33425;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33419;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33392;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33332;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33317;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33309;
    wire N__33304;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33288;
    wire N__33283;
    wire N__33278;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33254;
    wire N__33251;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33227;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33210;
    wire N__33203;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33175;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33149;
    wire N__33144;
    wire N__33139;
    wire N__33134;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33119;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33104;
    wire N__33101;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33089;
    wire N__33086;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33071;
    wire N__33068;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33056;
    wire N__33053;
    wire N__33052;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33035;
    wire N__33032;
    wire N__33031;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33014;
    wire N__33011;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32924;
    wire N__32921;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32890;
    wire N__32885;
    wire N__32882;
    wire N__32881;
    wire N__32876;
    wire N__32875;
    wire N__32874;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32869;
    wire N__32868;
    wire N__32867;
    wire N__32864;
    wire N__32857;
    wire N__32852;
    wire N__32849;
    wire N__32842;
    wire N__32837;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32806;
    wire N__32805;
    wire N__32802;
    wire N__32797;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32711;
    wire N__32710;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32696;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32637;
    wire N__32634;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32614;
    wire N__32609;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32568;
    wire N__32565;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32535;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32517;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32500;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32492;
    wire N__32491;
    wire N__32488;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32422;
    wire N__32421;
    wire N__32418;
    wire N__32417;
    wire N__32416;
    wire N__32415;
    wire N__32414;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32390;
    wire N__32389;
    wire N__32384;
    wire N__32381;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32357;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32345;
    wire N__32342;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32326;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32279;
    wire N__32278;
    wire N__32275;
    wire N__32274;
    wire N__32271;
    wire N__32266;
    wire N__32261;
    wire N__32260;
    wire N__32259;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32243;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32189;
    wire N__32188;
    wire N__32187;
    wire N__32186;
    wire N__32179;
    wire N__32178;
    wire N__32175;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32107;
    wire N__32104;
    wire N__32101;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32071;
    wire N__32068;
    wire N__32063;
    wire N__32060;
    wire N__32059;
    wire N__32056;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32045;
    wire N__32038;
    wire N__32035;
    wire N__32030;
    wire N__32027;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32009;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31991;
    wire N__31988;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31879;
    wire N__31878;
    wire N__31877;
    wire N__31876;
    wire N__31875;
    wire N__31870;
    wire N__31867;
    wire N__31866;
    wire N__31859;
    wire N__31856;
    wire N__31851;
    wire N__31848;
    wire N__31841;
    wire N__31840;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31830;
    wire N__31829;
    wire N__31828;
    wire N__31827;
    wire N__31824;
    wire N__31823;
    wire N__31822;
    wire N__31819;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31747;
    wire N__31736;
    wire N__31727;
    wire N__31726;
    wire N__31725;
    wire N__31724;
    wire N__31723;
    wire N__31722;
    wire N__31721;
    wire N__31716;
    wire N__31711;
    wire N__31704;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31690;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31670;
    wire N__31667;
    wire N__31660;
    wire N__31655;
    wire N__31654;
    wire N__31653;
    wire N__31652;
    wire N__31651;
    wire N__31648;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31602;
    wire N__31595;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31544;
    wire N__31541;
    wire N__31540;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31499;
    wire N__31498;
    wire N__31495;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31490;
    wire N__31487;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31477;
    wire N__31476;
    wire N__31475;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31449;
    wire N__31446;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31432;
    wire N__31427;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31415;
    wire N__31410;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31380;
    wire N__31373;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31362;
    wire N__31361;
    wire N__31360;
    wire N__31359;
    wire N__31358;
    wire N__31357;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31323;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31311;
    wire N__31308;
    wire N__31307;
    wire N__31304;
    wire N__31299;
    wire N__31296;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31272;
    wire N__31265;
    wire N__31256;
    wire N__31255;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31243;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31158;
    wire N__31149;
    wire N__31144;
    wire N__31143;
    wire N__31138;
    wire N__31135;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31093;
    wire N__31088;
    wire N__31085;
    wire N__31084;
    wire N__31083;
    wire N__31080;
    wire N__31079;
    wire N__31078;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30988;
    wire N__30987;
    wire N__30984;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30974;
    wire N__30973;
    wire N__30970;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30959;
    wire N__30958;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30921;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30905;
    wire N__30902;
    wire N__30897;
    wire N__30892;
    wire N__30889;
    wire N__30880;
    wire N__30869;
    wire N__30868;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30857;
    wire N__30856;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30852;
    wire N__30847;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30834;
    wire N__30829;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30821;
    wire N__30818;
    wire N__30813;
    wire N__30810;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30788;
    wire N__30785;
    wire N__30780;
    wire N__30777;
    wire N__30768;
    wire N__30759;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30738;
    wire N__30737;
    wire N__30736;
    wire N__30731;
    wire N__30730;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30717;
    wire N__30716;
    wire N__30715;
    wire N__30712;
    wire N__30711;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30642;
    wire N__30629;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30608;
    wire N__30607;
    wire N__30602;
    wire N__30599;
    wire N__30594;
    wire N__30591;
    wire N__30584;
    wire N__30583;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30575;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30567;
    wire N__30564;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30546;
    wire N__30545;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30533;
    wire N__30532;
    wire N__30531;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30506;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30490;
    wire N__30487;
    wire N__30482;
    wire N__30479;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30433;
    wire N__30430;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30394;
    wire N__30391;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30343;
    wire N__30342;
    wire N__30339;
    wire N__30334;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30308;
    wire N__30305;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30275;
    wire N__30272;
    wire N__30271;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30249;
    wire N__30246;
    wire N__30241;
    wire N__30236;
    wire N__30235;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30215;
    wire N__30214;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30186;
    wire N__30181;
    wire N__30176;
    wire N__30175;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30145;
    wire N__30140;
    wire N__30139;
    wire N__30138;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30121;
    wire N__30118;
    wire N__30113;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30101;
    wire N__30100;
    wire N__30099;
    wire N__30098;
    wire N__30097;
    wire N__30096;
    wire N__30093;
    wire N__30092;
    wire N__30091;
    wire N__30090;
    wire N__30089;
    wire N__30088;
    wire N__30087;
    wire N__30086;
    wire N__30085;
    wire N__30084;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30076;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30065;
    wire N__30056;
    wire N__30053;
    wire N__30052;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30048;
    wire N__30047;
    wire N__30046;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30041;
    wire N__30040;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30036;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30028;
    wire N__30027;
    wire N__30026;
    wire N__30025;
    wire N__30024;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__29994;
    wire N__29991;
    wire N__29982;
    wire N__29973;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29963;
    wire N__29962;
    wire N__29959;
    wire N__29952;
    wire N__29945;
    wire N__29940;
    wire N__29929;
    wire N__29928;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29914;
    wire N__29913;
    wire N__29912;
    wire N__29911;
    wire N__29910;
    wire N__29909;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29889;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29883;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29879;
    wire N__29866;
    wire N__29855;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29832;
    wire N__29823;
    wire N__29816;
    wire N__29803;
    wire N__29794;
    wire N__29785;
    wire N__29768;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29753;
    wire N__29750;
    wire N__29749;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29716;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29610;
    wire N__29609;
    wire N__29606;
    wire N__29601;
    wire N__29598;
    wire N__29593;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29568;
    wire N__29567;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29509;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29494;
    wire N__29491;
    wire N__29490;
    wire N__29489;
    wire N__29486;
    wire N__29485;
    wire N__29484;
    wire N__29483;
    wire N__29482;
    wire N__29481;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29467;
    wire N__29466;
    wire N__29463;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29449;
    wire N__29446;
    wire N__29441;
    wire N__29436;
    wire N__29431;
    wire N__29428;
    wire N__29427;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29392;
    wire N__29389;
    wire N__29388;
    wire N__29385;
    wire N__29374;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29344;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29308;
    wire N__29303;
    wire N__29302;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29279;
    wire N__29276;
    wire N__29275;
    wire N__29274;
    wire N__29273;
    wire N__29272;
    wire N__29269;
    wire N__29268;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29260;
    wire N__29259;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29245;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29237;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29222;
    wire N__29219;
    wire N__29218;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29196;
    wire N__29195;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29181;
    wire N__29174;
    wire N__29169;
    wire N__29166;
    wire N__29161;
    wire N__29158;
    wire N__29153;
    wire N__29148;
    wire N__29143;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29098;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29066;
    wire N__29063;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28954;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28918;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28879;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28704;
    wire N__28703;
    wire N__28702;
    wire N__28701;
    wire N__28700;
    wire N__28699;
    wire N__28694;
    wire N__28691;
    wire N__28690;
    wire N__28687;
    wire N__28686;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28674;
    wire N__28673;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28663;
    wire N__28660;
    wire N__28659;
    wire N__28658;
    wire N__28657;
    wire N__28654;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28606;
    wire N__28603;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28573;
    wire N__28570;
    wire N__28569;
    wire N__28568;
    wire N__28567;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28518;
    wire N__28515;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28497;
    wire N__28490;
    wire N__28487;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28468;
    wire N__28465;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28403;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28391;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28355;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28307;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28295;
    wire N__28292;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28277;
    wire N__28276;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28240;
    wire N__28239;
    wire N__28238;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28220;
    wire N__28217;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28205;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28177;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28169;
    wire N__28166;
    wire N__28161;
    wire N__28158;
    wire N__28153;
    wire N__28148;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28100;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28092;
    wire N__28087;
    wire N__28084;
    wire N__28079;
    wire N__28078;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28042;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28004;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27973;
    wire N__27972;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27958;
    wire N__27957;
    wire N__27956;
    wire N__27955;
    wire N__27950;
    wire N__27949;
    wire N__27948;
    wire N__27947;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27930;
    wire N__27927;
    wire N__27926;
    wire N__27925;
    wire N__27924;
    wire N__27923;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27907;
    wire N__27902;
    wire N__27899;
    wire N__27898;
    wire N__27897;
    wire N__27896;
    wire N__27895;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27877;
    wire N__27874;
    wire N__27867;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27839;
    wire N__27838;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27694;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27661;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27601;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27558;
    wire N__27557;
    wire N__27554;
    wire N__27549;
    wire N__27546;
    wire N__27541;
    wire N__27536;
    wire N__27533;
    wire N__27532;
    wire N__27531;
    wire N__27528;
    wire N__27527;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27504;
    wire N__27503;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27485;
    wire N__27482;
    wire N__27481;
    wire N__27478;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27455;
    wire N__27452;
    wire N__27451;
    wire N__27448;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27425;
    wire N__27422;
    wire N__27421;
    wire N__27418;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27302;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27121;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27117;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27109;
    wire N__27108;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27098;
    wire N__27093;
    wire N__27080;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27060;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26983;
    wire N__26980;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26944;
    wire N__26943;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26927;
    wire N__26924;
    wire N__26923;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26763;
    wire N__26762;
    wire N__26759;
    wire N__26754;
    wire N__26751;
    wire N__26746;
    wire N__26741;
    wire N__26740;
    wire N__26739;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26719;
    wire N__26716;
    wire N__26711;
    wire N__26708;
    wire N__26707;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26696;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26678;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26666;
    wire N__26663;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26578;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26488;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26443;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26260;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26231;
    wire N__26230;
    wire N__26229;
    wire N__26226;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26090;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26082;
    wire N__26081;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26051;
    wire N__26050;
    wire N__26047;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26009;
    wire N__26006;
    wire N__26005;
    wire N__26004;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25964;
    wire N__25963;
    wire N__25962;
    wire N__25959;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25923;
    wire N__25916;
    wire N__25913;
    wire N__25912;
    wire N__25911;
    wire N__25910;
    wire N__25907;
    wire N__25902;
    wire N__25901;
    wire N__25898;
    wire N__25897;
    wire N__25892;
    wire N__25885;
    wire N__25882;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25852;
    wire N__25847;
    wire N__25844;
    wire N__25843;
    wire N__25842;
    wire N__25841;
    wire N__25832;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25817;
    wire N__25814;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25756;
    wire N__25755;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25709;
    wire N__25706;
    wire N__25705;
    wire N__25704;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25660;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25637;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25619;
    wire N__25618;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25485;
    wire N__25482;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25460;
    wire N__25457;
    wire N__25456;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25397;
    wire N__25396;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25382;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25364;
    wire N__25363;
    wire N__25362;
    wire N__25359;
    wire N__25358;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25334;
    wire N__25333;
    wire N__25330;
    wire N__25325;
    wire N__25320;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25279;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25238;
    wire N__25237;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25229;
    wire N__25226;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25215;
    wire N__25210;
    wire N__25207;
    wire N__25202;
    wire N__25199;
    wire N__25190;
    wire N__25187;
    wire N__25186;
    wire N__25185;
    wire N__25184;
    wire N__25181;
    wire N__25176;
    wire N__25173;
    wire N__25168;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25141;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25058;
    wire N__25055;
    wire N__25054;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25004;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24997;
    wire N__24996;
    wire N__24993;
    wire N__24992;
    wire N__24991;
    wire N__24988;
    wire N__24987;
    wire N__24986;
    wire N__24985;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24981;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24957;
    wire N__24948;
    wire N__24947;
    wire N__24946;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24942;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24938;
    wire N__24937;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24921;
    wire N__24914;
    wire N__24909;
    wire N__24902;
    wire N__24897;
    wire N__24894;
    wire N__24883;
    wire N__24880;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24860;
    wire N__24859;
    wire N__24858;
    wire N__24855;
    wire N__24850;
    wire N__24841;
    wire N__24836;
    wire N__24831;
    wire N__24826;
    wire N__24823;
    wire N__24816;
    wire N__24801;
    wire N__24796;
    wire N__24793;
    wire N__24786;
    wire N__24773;
    wire N__24770;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24739;
    wire N__24738;
    wire N__24737;
    wire N__24734;
    wire N__24729;
    wire N__24726;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24618;
    wire N__24613;
    wire N__24608;
    wire N__24607;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24595;
    wire N__24592;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24573;
    wire N__24568;
    wire N__24565;
    wire N__24560;
    wire N__24559;
    wire N__24556;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24544;
    wire N__24541;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24515;
    wire N__24514;
    wire N__24509;
    wire N__24508;
    wire N__24507;
    wire N__24504;
    wire N__24499;
    wire N__24496;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24385;
    wire N__24382;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24352;
    wire N__24349;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24328;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24244;
    wire N__24241;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24225;
    wire N__24222;
    wire N__24217;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24153;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24137;
    wire N__24134;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24064;
    wire N__24063;
    wire N__24062;
    wire N__24059;
    wire N__24054;
    wire N__24051;
    wire N__24044;
    wire N__24041;
    wire N__24040;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23964;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23953;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23932;
    wire N__23917;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23909;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23853;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23787;
    wire N__23780;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23762;
    wire N__23759;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23741;
    wire N__23738;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23693;
    wire N__23690;
    wire N__23689;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23650;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23418;
    wire N__23413;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23361;
    wire N__23358;
    wire N__23353;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23296;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23284;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23264;
    wire N__23261;
    wire N__23254;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23237;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23212;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23194;
    wire N__23193;
    wire N__23192;
    wire N__23191;
    wire N__23188;
    wire N__23183;
    wire N__23178;
    wire N__23173;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23156;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23137;
    wire N__23132;
    wire N__23129;
    wire N__23122;
    wire N__23119;
    wire N__23114;
    wire N__23105;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23085;
    wire N__23084;
    wire N__23083;
    wire N__23082;
    wire N__23081;
    wire N__23080;
    wire N__23077;
    wire N__23076;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23064;
    wire N__23063;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23059;
    wire N__23056;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23041;
    wire N__23036;
    wire N__23031;
    wire N__23030;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23018;
    wire N__23011;
    wire N__23002;
    wire N__22997;
    wire N__22994;
    wire N__22989;
    wire N__22986;
    wire N__22985;
    wire N__22984;
    wire N__22983;
    wire N__22982;
    wire N__22979;
    wire N__22978;
    wire N__22971;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22948;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22944;
    wire N__22943;
    wire N__22942;
    wire N__22937;
    wire N__22928;
    wire N__22921;
    wire N__22916;
    wire N__22909;
    wire N__22902;
    wire N__22893;
    wire N__22888;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22788;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22628;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22610;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22585;
    wire N__22580;
    wire N__22577;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22539;
    wire N__22534;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22505;
    wire N__22504;
    wire N__22501;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22484;
    wire N__22483;
    wire N__22482;
    wire N__22481;
    wire N__22478;
    wire N__22473;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22451;
    wire N__22450;
    wire N__22447;
    wire N__22446;
    wire N__22443;
    wire N__22438;
    wire N__22433;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22421;
    wire N__22418;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22407;
    wire N__22406;
    wire N__22405;
    wire N__22402;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22361;
    wire N__22360;
    wire N__22359;
    wire N__22358;
    wire N__22355;
    wire N__22354;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22338;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22291;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22228;
    wire N__22225;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22199;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22179;
    wire N__22176;
    wire N__22163;
    wire N__22160;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22110;
    wire N__22107;
    wire N__22106;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22082;
    wire N__22079;
    wire N__22078;
    wire N__22075;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22048;
    wire N__22031;
    wire N__22030;
    wire N__22027;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22006;
    wire N__22003;
    wire N__22002;
    wire N__22001;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21963;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21937;
    wire N__21936;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21909;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21883;
    wire N__21882;
    wire N__21875;
    wire N__21872;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21829;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21701;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21689;
    wire N__21686;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21641;
    wire N__21638;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21628;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21624;
    wire N__21623;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21579;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21574;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21446;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21416;
    wire N__21415;
    wire N__21412;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21295;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21070;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21012;
    wire N__21009;
    wire N__21004;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20992;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20950;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20929;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20885;
    wire N__20882;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20874;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20862;
    wire N__20861;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20846;
    wire N__20845;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20817;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20789;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20775;
    wire N__20772;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20590;
    wire N__20585;
    wire N__20582;
    wire N__20581;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20508;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20435;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20399;
    wire N__20398;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20367;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20311;
    wire N__20310;
    wire N__20309;
    wire N__20308;
    wire N__20307;
    wire N__20306;
    wire N__20305;
    wire N__20304;
    wire N__20303;
    wire N__20302;
    wire N__20301;
    wire N__20300;
    wire N__20299;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20263;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20235;
    wire N__20230;
    wire N__20225;
    wire N__20224;
    wire N__20223;
    wire N__20222;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20197;
    wire N__20192;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20129;
    wire N__20126;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20121;
    wire N__20114;
    wire N__20109;
    wire N__20108;
    wire N__20107;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20101;
    wire N__20100;
    wire N__20095;
    wire N__20092;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20079;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20054;
    wire N__20049;
    wire N__20042;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20007;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19938;
    wire N__19937;
    wire N__19936;
    wire N__19935;
    wire N__19930;
    wire N__19923;
    wire N__19922;
    wire N__19921;
    wire N__19918;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19906;
    wire N__19901;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19833;
    wire N__19830;
    wire N__19825;
    wire N__19822;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19593;
    wire N__19588;
    wire N__19585;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19489;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19456;
    wire N__19451;
    wire N__19448;
    wire N__19447;
    wire N__19442;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19426;
    wire N__19425;
    wire N__19420;
    wire N__19419;
    wire N__19416;
    wire N__19415;
    wire N__19414;
    wire N__19413;
    wire N__19410;
    wire N__19403;
    wire N__19402;
    wire N__19399;
    wire N__19398;
    wire N__19395;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19342;
    wire N__19337;
    wire N__19336;
    wire N__19335;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19323;
    wire N__19322;
    wire N__19319;
    wire N__19310;
    wire N__19307;
    wire N__19302;
    wire N__19297;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19265;
    wire N__19262;
    wire N__19261;
    wire N__19260;
    wire N__19257;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19223;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19199;
    wire N__19198;
    wire N__19197;
    wire N__19192;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19169;
    wire N__19166;
    wire N__19165;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19146;
    wire N__19143;
    wire N__19138;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19013;
    wire N__19010;
    wire N__19009;
    wire N__19006;
    wire N__19005;
    wire N__19002;
    wire N__19001;
    wire N__19000;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18975;
    wire N__18968;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18953;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18870;
    wire N__18865;
    wire N__18862;
    wire N__18861;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18849;
    wire N__18846;
    wire N__18841;
    wire N__18836;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18817;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18803;
    wire N__18802;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18771;
    wire N__18766;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18680;
    wire N__18677;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18651;
    wire N__18646;
    wire N__18641;
    wire N__18638;
    wire N__18637;
    wire N__18636;
    wire N__18633;
    wire N__18628;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18597;
    wire N__18596;
    wire N__18591;
    wire N__18586;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18552;
    wire N__18549;
    wire N__18544;
    wire N__18539;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18509;
    wire N__18508;
    wire N__18507;
    wire N__18504;
    wire N__18499;
    wire N__18498;
    wire N__18493;
    wire N__18490;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18413;
    wire N__18412;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18371;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18357;
    wire N__18352;
    wire N__18349;
    wire N__18344;
    wire N__18343;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18312;
    wire N__18307;
    wire N__18304;
    wire N__18299;
    wire N__18298;
    wire N__18297;
    wire N__18296;
    wire N__18295;
    wire N__18294;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18264;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18248;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18203;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18144;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18119;
    wire N__18110;
    wire N__18109;
    wire N__18108;
    wire N__18105;
    wire N__18100;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18081;
    wire N__18076;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18064;
    wire N__18063;
    wire N__18060;
    wire N__18055;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18022;
    wire N__18019;
    wire N__18014;
    wire N__18011;
    wire N__18010;
    wire N__18009;
    wire N__18006;
    wire N__18001;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17986;
    wire N__17985;
    wire N__17982;
    wire N__17977;
    wire N__17972;
    wire N__17971;
    wire N__17968;
    wire N__17967;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17939;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17931;
    wire N__17928;
    wire N__17923;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17908;
    wire N__17907;
    wire N__17904;
    wire N__17899;
    wire N__17894;
    wire N__17893;
    wire N__17892;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17858;
    wire N__17857;
    wire N__17854;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17842;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17826;
    wire N__17823;
    wire N__17818;
    wire N__17813;
    wire N__17812;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17780;
    wire N__17777;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17741;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17692;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17656;
    wire N__17655;
    wire N__17652;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17622;
    wire N__17619;
    wire N__17614;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17587;
    wire N__17586;
    wire N__17583;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17553;
    wire N__17550;
    wire N__17545;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17512;
    wire N__17511;
    wire N__17508;
    wire N__17503;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17490;
    wire N__17487;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17471;
    wire N__17470;
    wire N__17467;
    wire N__17466;
    wire N__17465;
    wire N__17464;
    wire N__17461;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17442;
    wire N__17437;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17420;
    wire N__17417;
    wire N__17416;
    wire N__17415;
    wire N__17412;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17385;
    wire N__17378;
    wire N__17377;
    wire N__17374;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17345;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17329;
    wire N__17326;
    wire N__17325;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17313;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17296;
    wire N__17295;
    wire N__17292;
    wire N__17287;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17268;
    wire N__17265;
    wire N__17260;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17244;
    wire N__17241;
    wire N__17236;
    wire N__17231;
    wire N__17230;
    wire N__17227;
    wire N__17226;
    wire N__17225;
    wire N__17222;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17192;
    wire N__17189;
    wire N__17188;
    wire N__17187;
    wire N__17184;
    wire N__17179;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17115;
    wire N__17110;
    wire N__17105;
    wire N__17102;
    wire N__17101;
    wire N__17100;
    wire N__17097;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16910;
    wire N__16907;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16892;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16877;
    wire N__16874;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16866;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16274;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16219;
    wire N__16218;
    wire N__16211;
    wire N__16208;
    wire N__16207;
    wire N__16206;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16183;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16168;
    wire N__16165;
    wire N__16160;
    wire N__16159;
    wire N__16158;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16135;
    wire N__16134;
    wire N__16127;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16108;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16075;
    wire N__16074;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15329;
    wire N__15328;
    wire N__15327;
    wire N__15326;
    wire N__15325;
    wire N__15314;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15293;
    wire N__15290;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15261;
    wire N__15260;
    wire N__15255;
    wire N__15250;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15217;
    wire N__15216;
    wire N__15213;
    wire N__15212;
    wire N__15209;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15185;
    wire N__15180;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15159;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15095;
    wire N__15094;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15053;
    wire N__15050;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14822;
    wire N__14819;
    wire N__14818;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14780;
    wire N__14777;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14696;
    wire N__14693;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14500;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14434;
    wire N__14433;
    wire N__14430;
    wire N__14425;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14397;
    wire N__14392;
    wire N__14387;
    wire N__14384;
    wire N__14383;
    wire N__14382;
    wire N__14379;
    wire N__14374;
    wire N__14369;
    wire N__14368;
    wire N__14367;
    wire N__14364;
    wire N__14359;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14287;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14263;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14126;
    wire N__14125;
    wire N__14122;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14102;
    wire N__14101;
    wire N__14100;
    wire N__14097;
    wire N__14092;
    wire N__14087;
    wire N__14086;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14071;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14044;
    wire N__14043;
    wire N__14040;
    wire N__14035;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14020;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13948;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13834;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13810;
    wire N__13809;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13714;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire VCCG0;
    wire GNDG0;
    wire \pid_alt.O_0_6 ;
    wire \pid_alt.O_0_14 ;
    wire \pid_alt.O_0_12 ;
    wire \pid_alt.O_0_21 ;
    wire \pid_alt.O_0_7 ;
    wire \pid_alt.O_0_17 ;
    wire \pid_alt.O_0_15 ;
    wire \pid_alt.O_0_16 ;
    wire \pid_alt.O_0_5 ;
    wire \pid_alt.O_0_22 ;
    wire \pid_alt.O_0_4 ;
    wire \pid_alt.O_0_10 ;
    wire \pid_alt.O_0_23 ;
    wire \pid_alt.O_0_11 ;
    wire \pid_alt.O_0_13 ;
    wire \pid_alt.O_0_24 ;
    wire \pid_alt.O_0_19 ;
    wire \pid_alt.O_0_20 ;
    wire \pid_alt.O_0_18 ;
    wire \pid_alt.O_0_9 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.O_18 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.O_23 ;
    wire \pid_alt.O_4 ;
    wire \pid_alt.O_17 ;
    wire \pid_alt.O_19 ;
    wire \pid_alt.O_20 ;
    wire \pid_alt.O_21 ;
    wire \pid_alt.O_22 ;
    wire \pid_alt.O_6 ;
    wire \pid_alt.O_24 ;
    wire \pid_alt.O_15 ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_ ;
    wire \pid_alt.O_16 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.O_14 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.O_5 ;
    wire \pid_alt.O_7 ;
    wire \pid_alt.O_9 ;
    wire \pid_alt.O_8 ;
    wire \pid_alt.N_62_mux_cascade_ ;
    wire \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5 ;
    wire \pid_alt.N_37_cascade_ ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.N_37 ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire alt_ki_0;
    wire bfn_1_22_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire throttle_command_6;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_1_23_0_;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire scaler_2_data_5;
    wire \ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire throttle_command_9;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ;
    wire \pid_alt.O_0_8 ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire alt_kp_2;
    wire alt_ki_4;
    wire alt_ki_1;
    wire alt_ki_2;
    wire alt_ki_3;
    wire alt_ki_5;
    wire alt_ki_6;
    wire \pid_alt.O_12 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_ ;
    wire \pid_alt.O_13 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire bfn_2_11_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_2_12_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.m35_e_2_cascade_ ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5 ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.m21_e_2_cascade_ ;
    wire \pid_alt.m21_e_0_cascade_ ;
    wire \pid_alt.m21_e_8 ;
    wire bfn_2_14_0_;
    wire \scaler_2.un3_source_data_0_cry_0 ;
    wire \scaler_2.un3_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_7 ;
    wire bfn_2_15_0_;
    wire \scaler_2.un3_source_data_0_cry_8 ;
    wire \pid_alt.drone_altitude_i_0 ;
    wire drone_altitude_0;
    wire \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ;
    wire \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14 ;
    wire \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_ ;
    wire \pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_ ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.N_9_0_cascade_ ;
    wire \pid_alt.m21_e_10 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_ ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_alt.un1_reset_1_0_i_cascade_ ;
    wire \pid_alt.N_60_i_0 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire bfn_2_17_0_;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1 ;
    wire \pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2 ;
    wire \pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3 ;
    wire \pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5 ;
    wire \pid_alt.error_p_reg_esr_RNI91H61Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5 ;
    wire \pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire bfn_2_18_0_;
    wire \pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8 ;
    wire \pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9 ;
    wire \pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10 ;
    wire \pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12 ;
    wire \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13 ;
    wire \pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14 ;
    wire \pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire \pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14 ;
    wire \pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14 ;
    wire bfn_2_19_0_;
    wire \pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15 ;
    wire \pid_alt.error_p_reg_esr_RNIKU581Z0Z_15 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.error_p_reg_esr_RNIO2681Z0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_p_reg_esr_RNID23KZ0Z_17 ;
    wire \pid_alt.error_p_reg_esr_RNIS6681Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_p_reg_esr_RNI0B681Z0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.error_p_reg_esr_RNIIU781Z0Z_19 ;
    wire \pid_alt.error_p_reg_esr_RNIH63KZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.error_p_reg_esr_RNI2G981Z0Z_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_ ;
    wire \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_3 ;
    wire \pid_alt.source_pid_9_0_0_4 ;
    wire throttle_command_5;
    wire \ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.N_303_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire throttle_command_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.N_299_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_command_7;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5 ;
    wire \ppm_encoder_1.throttle_RNIN3352Z0Z_0 ;
    wire bfn_2_25_0_;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.throttle_RNIJII96Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire bfn_2_26_0_;
    wire \ppm_encoder_1.throttle_RNITSI96Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_2_27_0_;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ;
    wire bfn_2_28_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire bfn_2_29_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_2_30_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire alt_kp_3;
    wire alt_kp_6;
    wire alt_kp_5;
    wire alt_kp_1;
    wire alt_kp_0;
    wire drone_altitude_15;
    wire alt_command_2;
    wire alt_command_3;
    wire alt_command_1;
    wire \Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire alt_command_0;
    wire drone_altitude_i_7;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire drone_altitude_i_8;
    wire drone_altitude_i_9;
    wire drone_altitude_i_10;
    wire drone_altitude_i_11;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire drone_altitude_1;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire drone_altitude_12;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire drone_altitude_13;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire bfn_3_13_0_;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire bfn_3_14_0_;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire bfn_3_15_0_;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.state_0_g_0 ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire \pid_alt.error_p_reg_esr_RNIB03KZ0Z_16 ;
    wire \ppm_encoder_1.N_306 ;
    wire \dron_frame_decoder_1.N_194_4_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.m7_e_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO ;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.source_pid_9_0_tz_6 ;
    wire \pid_alt.source_pid_9_0_tz_6_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ;
    wire \pid_alt.N_92_cascade_ ;
    wire \pid_alt.un1_reset_1_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ;
    wire \pid_alt.un1_reset_0_i_cascade_ ;
    wire bfn_3_21_0_;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire bfn_3_22_0_;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6 ;
    wire \pid_alt.N_88 ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.N_88_cascade_ ;
    wire \pid_alt.N_90 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.N_90_cascade_ ;
    wire \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ;
    wire \pid_alt.N_60_i_1 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.N_130 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIALN65Z0Z_1 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ;
    wire \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.throttle_RNI5V123Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.throttle_RNI82223Z0Z_3 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0 ;
    wire \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.N_319_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire alt_kp_7;
    wire alt_kp_4;
    wire \pid_alt.O_10 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6 ;
    wire \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_ ;
    wire \pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7 ;
    wire \pid_alt.O_11 ;
    wire \pid_alt.N_422_0_g ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7 ;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire drone_altitude_14;
    wire drone_altitude_2;
    wire drone_altitude_3;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_p_reg_esr_RNIF43KZ0Z_18 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20 ;
    wire frame_decoder_CH2data_1;
    wire frame_decoder_CH2data_2;
    wire frame_decoder_CH2data_3;
    wire frame_decoder_CH2data_4;
    wire frame_decoder_CH2data_5;
    wire frame_decoder_CH2data_6;
    wire \scaler_2.N_881_i_l_ofxZ0 ;
    wire frame_decoder_CH2data_7;
    wire \scaler_2.un3_source_data_0_axb_7 ;
    wire \scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_4_16_0_;
    wire \scaler_2.un2_source_data_0 ;
    wire \scaler_2.un2_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_1_c_RNI14IK ;
    wire scaler_2_data_7;
    wire \scaler_2.un2_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_2_c_RNI48JK ;
    wire \scaler_2.un2_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ;
    wire scaler_2_data_9;
    wire \scaler_2.un2_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ;
    wire \scaler_2.un2_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ;
    wire scaler_2_data_11;
    wire \scaler_2.un2_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ;
    wire \scaler_2.un2_source_data_0_cry_7 ;
    wire \scaler_2.un2_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ;
    wire \scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ;
    wire bfn_4_17_0_;
    wire \scaler_2.un2_source_data_0_cry_9 ;
    wire scaler_2_data_14;
    wire alt_ki_7;
    wire \pid_alt.un1_pid_prereg_0_axb_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0_THRU_CO ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire N_423_g;
    wire \pid_alt.N_422_0 ;
    wire \pid_alt.state_1_0_0 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire throttle_command_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire throttle_command_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_command_2;
    wire throttle_command_4;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.N_304_cascade_ ;
    wire scaler_2_data_12;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire throttle_command_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIONI96Z0Z_8 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8 ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire throttle_command_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire scaler_2_data_8;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.N_296 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4 ;
    wire \ppm_encoder_1.N_227 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.N_302_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ;
    wire \ppm_encoder_1.N_145_17_cascade_ ;
    wire \ppm_encoder_1.N_145_17 ;
    wire \ppm_encoder_1.N_238_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.N_300 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.N_301 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire drone_altitude_i_4;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire drone_altitude_i_5;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire drone_altitude_i_6;
    wire alt_command_4;
    wire alt_command_5;
    wire alt_command_6;
    wire alt_command_7;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire frame_decoder_OFF2data_1;
    wire frame_decoder_OFF2data_2;
    wire frame_decoder_OFF2data_3;
    wire frame_decoder_OFF2data_4;
    wire frame_decoder_OFF2data_5;
    wire frame_decoder_OFF2data_6;
    wire frame_decoder_OFF2data_7;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.state_RNO_1Z0Z_0 ;
    wire \dron_frame_decoder_1.N_194_4 ;
    wire \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ;
    wire \dron_frame_decoder_1.state_RNO_0Z0Z_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_1 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3 ;
    wire debug_CH1_0A_c;
    wire \pid_alt.N_60_i ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire frame_decoder_OFF2data_0;
    wire frame_decoder_CH2data_0;
    wire scaler_2_data_4;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire scaler_2_data_10;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire scaler_2_data_13;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire bfn_5_22_0_;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire bfn_5_23_0_;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire scaler_2_data_6;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire throttle_command_0;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_command_1;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire throttle_command_3;
    wire pid_altitude_dv;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.N_140_0_cascade_ ;
    wire \ppm_encoder_1.N_145 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_5_27_0_;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_5_28_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.N_238 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire bfn_5_29_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_5_30_0_;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \dron_frame_decoder_1.N_390_0 ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ;
    wire \dron_frame_decoder_1.N_382_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_3_2 ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire uart_drone_data_0;
    wire uart_drone_data_1;
    wire uart_drone_data_2;
    wire uart_drone_data_3;
    wire uart_drone_data_4;
    wire uart_drone_data_5;
    wire uart_drone_data_6;
    wire uart_drone_data_7;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire bfn_7_19_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_OFF4data_2;
    wire frame_decoder_CH4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_OFF4data_4;
    wire frame_decoder_CH4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire bfn_7_20_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.N_905_i_l_ofxZ0 ;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNO_1 ;
    wire bfn_7_21_0_;
    wire scaler_4_data_6;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire scaler_4_data_7;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire scaler_4_data_8;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire scaler_4_data_9;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire scaler_4_data_10;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire scaler_4_data_11;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire scaler_4_data_12;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire scaler_4_data_13;
    wire bfn_7_22_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire \scaler_4.un2_source_data_0 ;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_CH4data_0;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire scaler_4_data_4;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire scaler_4_data_5;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.N_1014_0 ;
    wire \ppm_encoder_1.N_1014_i ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_7_26_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire bfn_7_27_0_;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_7_28_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_320_g ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_1_1_0 ;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ;
    wire frame_decoder_OFF4data_7;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire bfn_8_20_0_;
    wire frame_decoder_CH3data_1;
    wire frame_decoder_OFF3data_1;
    wire \scaler_3.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH3data_2;
    wire frame_decoder_OFF3data_2;
    wire \scaler_3.un3_source_data_0_cry_1 ;
    wire frame_decoder_OFF3data_3;
    wire frame_decoder_CH3data_3;
    wire \scaler_3.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH3data_4;
    wire frame_decoder_OFF3data_4;
    wire \scaler_3.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH3data_5;
    wire frame_decoder_OFF3data_5;
    wire \scaler_3.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH3data_6;
    wire frame_decoder_OFF3data_6;
    wire \scaler_3.un3_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_axb_7 ;
    wire \scaler_3.un3_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_7 ;
    wire CONSTANT_ONE_NET;
    wire bfn_8_21_0_;
    wire \scaler_3.un3_source_data_0_cry_8 ;
    wire frame_decoder_OFF3data_7;
    wire frame_decoder_CH3data_7;
    wire \scaler_3.N_893_i_l_ofxZ0 ;
    wire \scaler_3.un2_source_data_0_cry_1_c_RNO_0 ;
    wire bfn_8_22_0_;
    wire scaler_3_data_6;
    wire \scaler_3.un2_source_data_0_cry_1 ;
    wire \scaler_3.un3_source_data_0_cry_1_c_RNI44VK ;
    wire scaler_3_data_7;
    wire \scaler_3.un2_source_data_0_cry_2 ;
    wire \scaler_3.un3_source_data_0_cry_2_c_RNI780L ;
    wire scaler_3_data_8;
    wire \scaler_3.un2_source_data_0_cry_3 ;
    wire \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ;
    wire scaler_3_data_9;
    wire \scaler_3.un2_source_data_0_cry_4 ;
    wire \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ;
    wire scaler_3_data_10;
    wire \scaler_3.un2_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ;
    wire scaler_3_data_11;
    wire \scaler_3.un2_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_6_c_RNILUAN ;
    wire scaler_3_data_12;
    wire \scaler_3.un2_source_data_0_cry_7 ;
    wire \scaler_3.un2_source_data_0_cry_8 ;
    wire \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ;
    wire \scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ;
    wire scaler_3_data_13;
    wire bfn_8_23_0_;
    wire \scaler_3.un2_source_data_0_cry_9 ;
    wire scaler_3_data_14;
    wire \scaler_3.un2_source_data_0 ;
    wire scaler_3_data_5;
    wire debug_CH3_20A_c_0_g;
    wire \ppm_encoder_1.N_305 ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.N_320 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_159_d ;
    wire \ppm_encoder_1.PPM_STATE_59_d ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ;
    wire \Commands_frame_decoder.N_338 ;
    wire \Commands_frame_decoder.N_309_cascade_ ;
    wire uart_pc_data_7;
    wire uart_pc_data_2;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ;
    wire uart_pc_data_5;
    wire \Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ;
    wire \Commands_frame_decoder.N_342 ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.N_308_2 ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.N_308_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_1_0 ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_0 ;
    wire uart_pc_data_0;
    wire uart_pc_data_6;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire uart_pc_data_3;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire uart_pc_data_1;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire uart_pc_data_4;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lto13_1 ;
    wire \dron_frame_decoder_1.WDT10lt14_0 ;
    wire \dron_frame_decoder_1.WDT10lt14_0_cascade_ ;
    wire \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire frame_decoder_OFF3data_0;
    wire frame_decoder_CH3data_0;
    wire scaler_3_data_4;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire bfn_10_11_0_;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire uart_drone_data_rdy;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire \Commands_frame_decoder.state_ns_i_a3_1_0_0 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.N_143_cascade_ ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_pc.state_srsts_i_0_2 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.N_145 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_144_1_cascade_ ;
    wire \uart_drone.N_144_1 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_pc.un1_state_2_0_cascade_ ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \Commands_frame_decoder.WDT8lto13_1_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ;
    wire \Commands_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.N_303_0 ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.N_335 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_10_19_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire bfn_10_20_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_1 ;
    wire \Commands_frame_decoder.CO0_cascade_ ;
    wire \Commands_frame_decoder.CO0 ;
    wire \Commands_frame_decoder.countZ0Z_1 ;
    wire \Commands_frame_decoder.countZ0Z_2 ;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.count_RNIDLVE1Z0Z_2 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_11_15_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire bfn_11_16_0_;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.un1_state51_iZ0 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.data_rdyc_1 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.CO0 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.un1_state_2_0 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.state_0_0 ;
    wire \reset_module_System.reset6_15_cascade_ ;
    wire bfn_12_13_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire bfn_12_14_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_12_15_0_;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire bfn_12_17_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire reset_system;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.reset6_3_cascade_ ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_11 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_drone.un1_state_7_0_cascade_ ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.CO0 ;
    wire \uart_drone.N_152 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire debug_CH3_20A_c;
    wire reset_system_g;
    wire debug_CH3_20A_c_0;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;

    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28718),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28717),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__14840,N__14867,N__14891,N__14915,N__14942,N__14969,N__14996,N__15023,N__14636,N__14666,N__14693,N__14722,N__14750,N__14777,N__14804,N__15362}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__20501,N__16982,N__16970,N__20489,N__16772,N__14483,N__16958,N__16946}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_0_24 ,\pid_alt.O_0_23 ,\pid_alt.O_0_22 ,\pid_alt.O_0_21 ,\pid_alt.O_0_20 ,\pid_alt.O_0_19 ,\pid_alt.O_0_18 ,\pid_alt.O_0_17 ,\pid_alt.O_0_16 ,\pid_alt.O_0_15 ,\pid_alt.O_0_14 ,\pid_alt.O_0_13 ,\pid_alt.O_0_12 ,\pid_alt.O_0_11 ,\pid_alt.O_0_10 ,\pid_alt.O_0_9 ,\pid_alt.O_0_8 ,\pid_alt.O_0_7 ,\pid_alt.O_0_6 ,\pid_alt.O_0_5 ,\pid_alt.O_0_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28699),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28704),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__14833,N__14860,N__14884,N__14908,N__14935,N__14965,N__14992,N__15019,N__14632,N__14662,N__14692,N__14723,N__14749,N__14776,N__14803,N__15358}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__21149,N__14567,N__14579,N__14471,N__14591,N__14606,N__14459,N__14144}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_24 ,\pid_alt.O_23 ,\pid_alt.O_22 ,\pid_alt.O_21 ,\pid_alt.O_20 ,\pid_alt.O_19 ,\pid_alt.O_18 ,\pid_alt.O_17 ,\pid_alt.O_16 ,\pid_alt.O_15 ,\pid_alt.O_14 ,\pid_alt.O_13 ,\pid_alt.O_12 ,\pid_alt.O_11 ,\pid_alt.O_10 ,\pid_alt.O_9 ,\pid_alt.O_8 ,\pid_alt.O_7 ,\pid_alt.O_6 ,\pid_alt.O_5 ,\pid_alt.O_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__37455),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__37457),
            .DIN(N__37456),
            .DOUT(N__37455),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__37457),
            .PADOUT(N__37456),
            .PADIN(N__37455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__37446),
            .DIN(N__37445),
            .DOUT(N__37444),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__37446),
            .PADOUT(N__37445),
            .PADIN(N__37444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__37437),
            .DIN(N__37436),
            .DOUT(N__37435),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__37437),
            .PADOUT(N__37436),
            .PADIN(N__37435),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__37428),
            .DIN(N__37427),
            .DOUT(N__37426),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__37428),
            .PADOUT(N__37427),
            .PADIN(N__37426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36338),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__37419),
            .DIN(N__37418),
            .DOUT(N__37417),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__37419),
            .PADOUT(N__37418),
            .PADIN(N__37417),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__37410),
            .DIN(N__37409),
            .DOUT(N__37408),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__37410),
            .PADOUT(N__37409),
            .PADIN(N__37408),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__37401),
            .DIN(N__37400),
            .DOUT(N__37399),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__37401),
            .PADOUT(N__37400),
            .PADIN(N__37399),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__37392),
            .DIN(N__37391),
            .DOUT(N__37390),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__37392),
            .PADOUT(N__37391),
            .PADIN(N__37390),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__37383),
            .DIN(N__37382),
            .DOUT(N__37381),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__37383),
            .PADOUT(N__37382),
            .PADIN(N__37381),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__37374),
            .DIN(N__37373),
            .DOUT(N__37372),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__37374),
            .PADOUT(N__37373),
            .PADIN(N__37372),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24710),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__37365),
            .DIN(N__37364),
            .DOUT(N__37363),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__37365),
            .PADOUT(N__37364),
            .PADIN(N__37363),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36976),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__9045 (
            .O(N__37346),
            .I(\uart_drone.un1_state_7_0_cascade_ ));
    CascadeMux I__9044 (
            .O(N__37343),
            .I(N__37340));
    InMux I__9043 (
            .O(N__37340),
            .I(N__37337));
    LocalMux I__9042 (
            .O(N__37337),
            .I(\uart_drone.un1_state_7_0 ));
    InMux I__9041 (
            .O(N__37334),
            .I(N__37331));
    LocalMux I__9040 (
            .O(N__37331),
            .I(\uart_drone.CO0 ));
    InMux I__9039 (
            .O(N__37328),
            .I(N__37322));
    InMux I__9038 (
            .O(N__37327),
            .I(N__37319));
    InMux I__9037 (
            .O(N__37326),
            .I(N__37316));
    InMux I__9036 (
            .O(N__37325),
            .I(N__37313));
    LocalMux I__9035 (
            .O(N__37322),
            .I(N__37310));
    LocalMux I__9034 (
            .O(N__37319),
            .I(N__37307));
    LocalMux I__9033 (
            .O(N__37316),
            .I(N__37304));
    LocalMux I__9032 (
            .O(N__37313),
            .I(N__37299));
    Span4Mux_h I__9031 (
            .O(N__37310),
            .I(N__37299));
    Span4Mux_h I__9030 (
            .O(N__37307),
            .I(N__37296));
    Odrv4 I__9029 (
            .O(N__37304),
            .I(\uart_drone.N_152 ));
    Odrv4 I__9028 (
            .O(N__37299),
            .I(\uart_drone.N_152 ));
    Odrv4 I__9027 (
            .O(N__37296),
            .I(\uart_drone.N_152 ));
    InMux I__9026 (
            .O(N__37289),
            .I(N__37283));
    InMux I__9025 (
            .O(N__37288),
            .I(N__37278));
    InMux I__9024 (
            .O(N__37287),
            .I(N__37278));
    InMux I__9023 (
            .O(N__37286),
            .I(N__37275));
    LocalMux I__9022 (
            .O(N__37283),
            .I(N__37272));
    LocalMux I__9021 (
            .O(N__37278),
            .I(N__37267));
    LocalMux I__9020 (
            .O(N__37275),
            .I(N__37267));
    Span4Mux_v I__9019 (
            .O(N__37272),
            .I(N__37264));
    Span4Mux_h I__9018 (
            .O(N__37267),
            .I(N__37261));
    Odrv4 I__9017 (
            .O(N__37264),
            .I(\uart_drone.un1_state_4_0 ));
    Odrv4 I__9016 (
            .O(N__37261),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__9015 (
            .O(N__37256),
            .I(N__37252));
    InMux I__9014 (
            .O(N__37255),
            .I(N__37248));
    LocalMux I__9013 (
            .O(N__37252),
            .I(N__37244));
    InMux I__9012 (
            .O(N__37251),
            .I(N__37241));
    LocalMux I__9011 (
            .O(N__37248),
            .I(N__37237));
    InMux I__9010 (
            .O(N__37247),
            .I(N__37233));
    Span4Mux_v I__9009 (
            .O(N__37244),
            .I(N__37228));
    LocalMux I__9008 (
            .O(N__37241),
            .I(N__37228));
    CascadeMux I__9007 (
            .O(N__37240),
            .I(N__37223));
    Span4Mux_h I__9006 (
            .O(N__37237),
            .I(N__37220));
    InMux I__9005 (
            .O(N__37236),
            .I(N__37217));
    LocalMux I__9004 (
            .O(N__37233),
            .I(N__37212));
    Span4Mux_h I__9003 (
            .O(N__37228),
            .I(N__37212));
    InMux I__9002 (
            .O(N__37227),
            .I(N__37209));
    InMux I__9001 (
            .O(N__37226),
            .I(N__37204));
    InMux I__9000 (
            .O(N__37223),
            .I(N__37204));
    Odrv4 I__8999 (
            .O(N__37220),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__8998 (
            .O(N__37217),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__8997 (
            .O(N__37212),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__8996 (
            .O(N__37209),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__8995 (
            .O(N__37204),
            .I(\uart_drone.stateZ0Z_3 ));
    InMux I__8994 (
            .O(N__37193),
            .I(N__37186));
    InMux I__8993 (
            .O(N__37192),
            .I(N__37176));
    InMux I__8992 (
            .O(N__37191),
            .I(N__37176));
    InMux I__8991 (
            .O(N__37190),
            .I(N__37176));
    InMux I__8990 (
            .O(N__37189),
            .I(N__37176));
    LocalMux I__8989 (
            .O(N__37186),
            .I(N__37171));
    InMux I__8988 (
            .O(N__37185),
            .I(N__37168));
    LocalMux I__8987 (
            .O(N__37176),
            .I(N__37165));
    InMux I__8986 (
            .O(N__37175),
            .I(N__37162));
    InMux I__8985 (
            .O(N__37174),
            .I(N__37158));
    Span4Mux_v I__8984 (
            .O(N__37171),
            .I(N__37149));
    LocalMux I__8983 (
            .O(N__37168),
            .I(N__37149));
    Span4Mux_v I__8982 (
            .O(N__37165),
            .I(N__37149));
    LocalMux I__8981 (
            .O(N__37162),
            .I(N__37149));
    InMux I__8980 (
            .O(N__37161),
            .I(N__37146));
    LocalMux I__8979 (
            .O(N__37158),
            .I(N__37143));
    Span4Mux_h I__8978 (
            .O(N__37149),
            .I(N__37140));
    LocalMux I__8977 (
            .O(N__37146),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__8976 (
            .O(N__37143),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__8975 (
            .O(N__37140),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__8974 (
            .O(N__37133),
            .I(N__37128));
    CascadeMux I__8973 (
            .O(N__37132),
            .I(N__37123));
    CascadeMux I__8972 (
            .O(N__37131),
            .I(N__37120));
    LocalMux I__8971 (
            .O(N__37128),
            .I(N__37114));
    InMux I__8970 (
            .O(N__37127),
            .I(N__37111));
    InMux I__8969 (
            .O(N__37126),
            .I(N__37108));
    InMux I__8968 (
            .O(N__37123),
            .I(N__37097));
    InMux I__8967 (
            .O(N__37120),
            .I(N__37097));
    InMux I__8966 (
            .O(N__37119),
            .I(N__37097));
    InMux I__8965 (
            .O(N__37118),
            .I(N__37097));
    InMux I__8964 (
            .O(N__37117),
            .I(N__37094));
    Span4Mux_v I__8963 (
            .O(N__37114),
            .I(N__37087));
    LocalMux I__8962 (
            .O(N__37111),
            .I(N__37087));
    LocalMux I__8961 (
            .O(N__37108),
            .I(N__37087));
    InMux I__8960 (
            .O(N__37107),
            .I(N__37082));
    InMux I__8959 (
            .O(N__37106),
            .I(N__37082));
    LocalMux I__8958 (
            .O(N__37097),
            .I(N__37079));
    LocalMux I__8957 (
            .O(N__37094),
            .I(N__37076));
    Span4Mux_h I__8956 (
            .O(N__37087),
            .I(N__37073));
    LocalMux I__8955 (
            .O(N__37082),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__8954 (
            .O(N__37079),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__8953 (
            .O(N__37076),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__8952 (
            .O(N__37073),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__8951 (
            .O(N__37064),
            .I(N__37052));
    InMux I__8950 (
            .O(N__37063),
            .I(N__37052));
    InMux I__8949 (
            .O(N__37062),
            .I(N__37052));
    InMux I__8948 (
            .O(N__37061),
            .I(N__37052));
    LocalMux I__8947 (
            .O(N__37052),
            .I(N__37047));
    InMux I__8946 (
            .O(N__37051),
            .I(N__37044));
    CascadeMux I__8945 (
            .O(N__37050),
            .I(N__37038));
    Span4Mux_v I__8944 (
            .O(N__37047),
            .I(N__37033));
    LocalMux I__8943 (
            .O(N__37044),
            .I(N__37033));
    InMux I__8942 (
            .O(N__37043),
            .I(N__37030));
    InMux I__8941 (
            .O(N__37042),
            .I(N__37025));
    InMux I__8940 (
            .O(N__37041),
            .I(N__37022));
    InMux I__8939 (
            .O(N__37038),
            .I(N__37019));
    Span4Mux_h I__8938 (
            .O(N__37033),
            .I(N__37016));
    LocalMux I__8937 (
            .O(N__37030),
            .I(N__37013));
    InMux I__8936 (
            .O(N__37029),
            .I(N__37010));
    InMux I__8935 (
            .O(N__37028),
            .I(N__37007));
    LocalMux I__8934 (
            .O(N__37025),
            .I(N__37004));
    LocalMux I__8933 (
            .O(N__37022),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__8932 (
            .O(N__37019),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__8931 (
            .O(N__37016),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv12 I__8930 (
            .O(N__37013),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__8929 (
            .O(N__37010),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__8928 (
            .O(N__37007),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv12 I__8927 (
            .O(N__37004),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__8926 (
            .O(N__36989),
            .I(N__36986));
    LocalMux I__8925 (
            .O(N__36986),
            .I(N__36983));
    Span4Mux_h I__8924 (
            .O(N__36983),
            .I(N__36980));
    Odrv4 I__8923 (
            .O(N__36980),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__8922 (
            .O(N__36977),
            .I(N__36973));
    IoInMux I__8921 (
            .O(N__36976),
            .I(N__36970));
    LocalMux I__8920 (
            .O(N__36973),
            .I(N__36966));
    LocalMux I__8919 (
            .O(N__36970),
            .I(N__36962));
    InMux I__8918 (
            .O(N__36969),
            .I(N__36959));
    Span4Mux_v I__8917 (
            .O(N__36966),
            .I(N__36955));
    InMux I__8916 (
            .O(N__36965),
            .I(N__36952));
    Span12Mux_s11_v I__8915 (
            .O(N__36962),
            .I(N__36949));
    LocalMux I__8914 (
            .O(N__36959),
            .I(N__36946));
    InMux I__8913 (
            .O(N__36958),
            .I(N__36943));
    Span4Mux_v I__8912 (
            .O(N__36955),
            .I(N__36939));
    LocalMux I__8911 (
            .O(N__36952),
            .I(N__36936));
    Span12Mux_h I__8910 (
            .O(N__36949),
            .I(N__36929));
    Span12Mux_h I__8909 (
            .O(N__36946),
            .I(N__36929));
    LocalMux I__8908 (
            .O(N__36943),
            .I(N__36929));
    InMux I__8907 (
            .O(N__36942),
            .I(N__36926));
    Sp12to4 I__8906 (
            .O(N__36939),
            .I(N__36921));
    Span12Mux_v I__8905 (
            .O(N__36936),
            .I(N__36921));
    Odrv12 I__8904 (
            .O(N__36929),
            .I(debug_CH3_20A_c));
    LocalMux I__8903 (
            .O(N__36926),
            .I(debug_CH3_20A_c));
    Odrv12 I__8902 (
            .O(N__36921),
            .I(debug_CH3_20A_c));
    CascadeMux I__8901 (
            .O(N__36914),
            .I(N__36906));
    CascadeMux I__8900 (
            .O(N__36913),
            .I(N__36903));
    InMux I__8899 (
            .O(N__36912),
            .I(N__36870));
    InMux I__8898 (
            .O(N__36911),
            .I(N__36867));
    InMux I__8897 (
            .O(N__36910),
            .I(N__36864));
    InMux I__8896 (
            .O(N__36909),
            .I(N__36851));
    InMux I__8895 (
            .O(N__36906),
            .I(N__36851));
    InMux I__8894 (
            .O(N__36903),
            .I(N__36851));
    InMux I__8893 (
            .O(N__36902),
            .I(N__36851));
    InMux I__8892 (
            .O(N__36901),
            .I(N__36851));
    InMux I__8891 (
            .O(N__36900),
            .I(N__36851));
    InMux I__8890 (
            .O(N__36899),
            .I(N__36846));
    InMux I__8889 (
            .O(N__36898),
            .I(N__36846));
    InMux I__8888 (
            .O(N__36897),
            .I(N__36843));
    InMux I__8887 (
            .O(N__36896),
            .I(N__36840));
    InMux I__8886 (
            .O(N__36895),
            .I(N__36837));
    InMux I__8885 (
            .O(N__36894),
            .I(N__36834));
    InMux I__8884 (
            .O(N__36893),
            .I(N__36831));
    InMux I__8883 (
            .O(N__36892),
            .I(N__36828));
    InMux I__8882 (
            .O(N__36891),
            .I(N__36825));
    InMux I__8881 (
            .O(N__36890),
            .I(N__36822));
    InMux I__8880 (
            .O(N__36889),
            .I(N__36817));
    InMux I__8879 (
            .O(N__36888),
            .I(N__36817));
    InMux I__8878 (
            .O(N__36887),
            .I(N__36814));
    InMux I__8877 (
            .O(N__36886),
            .I(N__36811));
    InMux I__8876 (
            .O(N__36885),
            .I(N__36808));
    InMux I__8875 (
            .O(N__36884),
            .I(N__36805));
    InMux I__8874 (
            .O(N__36883),
            .I(N__36802));
    InMux I__8873 (
            .O(N__36882),
            .I(N__36799));
    InMux I__8872 (
            .O(N__36881),
            .I(N__36794));
    InMux I__8871 (
            .O(N__36880),
            .I(N__36794));
    InMux I__8870 (
            .O(N__36879),
            .I(N__36791));
    InMux I__8869 (
            .O(N__36878),
            .I(N__36788));
    InMux I__8868 (
            .O(N__36877),
            .I(N__36785));
    InMux I__8867 (
            .O(N__36876),
            .I(N__36782));
    InMux I__8866 (
            .O(N__36875),
            .I(N__36779));
    InMux I__8865 (
            .O(N__36874),
            .I(N__36774));
    InMux I__8864 (
            .O(N__36873),
            .I(N__36774));
    LocalMux I__8863 (
            .O(N__36870),
            .I(N__36686));
    LocalMux I__8862 (
            .O(N__36867),
            .I(N__36683));
    LocalMux I__8861 (
            .O(N__36864),
            .I(N__36680));
    LocalMux I__8860 (
            .O(N__36851),
            .I(N__36677));
    LocalMux I__8859 (
            .O(N__36846),
            .I(N__36674));
    LocalMux I__8858 (
            .O(N__36843),
            .I(N__36671));
    LocalMux I__8857 (
            .O(N__36840),
            .I(N__36668));
    LocalMux I__8856 (
            .O(N__36837),
            .I(N__36665));
    LocalMux I__8855 (
            .O(N__36834),
            .I(N__36662));
    LocalMux I__8854 (
            .O(N__36831),
            .I(N__36659));
    LocalMux I__8853 (
            .O(N__36828),
            .I(N__36656));
    LocalMux I__8852 (
            .O(N__36825),
            .I(N__36653));
    LocalMux I__8851 (
            .O(N__36822),
            .I(N__36650));
    LocalMux I__8850 (
            .O(N__36817),
            .I(N__36647));
    LocalMux I__8849 (
            .O(N__36814),
            .I(N__36644));
    LocalMux I__8848 (
            .O(N__36811),
            .I(N__36641));
    LocalMux I__8847 (
            .O(N__36808),
            .I(N__36638));
    LocalMux I__8846 (
            .O(N__36805),
            .I(N__36635));
    LocalMux I__8845 (
            .O(N__36802),
            .I(N__36632));
    LocalMux I__8844 (
            .O(N__36799),
            .I(N__36629));
    LocalMux I__8843 (
            .O(N__36794),
            .I(N__36626));
    LocalMux I__8842 (
            .O(N__36791),
            .I(N__36623));
    LocalMux I__8841 (
            .O(N__36788),
            .I(N__36620));
    LocalMux I__8840 (
            .O(N__36785),
            .I(N__36617));
    LocalMux I__8839 (
            .O(N__36782),
            .I(N__36614));
    LocalMux I__8838 (
            .O(N__36779),
            .I(N__36611));
    LocalMux I__8837 (
            .O(N__36774),
            .I(N__36608));
    SRMux I__8836 (
            .O(N__36773),
            .I(N__36383));
    SRMux I__8835 (
            .O(N__36772),
            .I(N__36383));
    SRMux I__8834 (
            .O(N__36771),
            .I(N__36383));
    SRMux I__8833 (
            .O(N__36770),
            .I(N__36383));
    SRMux I__8832 (
            .O(N__36769),
            .I(N__36383));
    SRMux I__8831 (
            .O(N__36768),
            .I(N__36383));
    SRMux I__8830 (
            .O(N__36767),
            .I(N__36383));
    SRMux I__8829 (
            .O(N__36766),
            .I(N__36383));
    SRMux I__8828 (
            .O(N__36765),
            .I(N__36383));
    SRMux I__8827 (
            .O(N__36764),
            .I(N__36383));
    SRMux I__8826 (
            .O(N__36763),
            .I(N__36383));
    SRMux I__8825 (
            .O(N__36762),
            .I(N__36383));
    SRMux I__8824 (
            .O(N__36761),
            .I(N__36383));
    SRMux I__8823 (
            .O(N__36760),
            .I(N__36383));
    SRMux I__8822 (
            .O(N__36759),
            .I(N__36383));
    SRMux I__8821 (
            .O(N__36758),
            .I(N__36383));
    SRMux I__8820 (
            .O(N__36757),
            .I(N__36383));
    SRMux I__8819 (
            .O(N__36756),
            .I(N__36383));
    SRMux I__8818 (
            .O(N__36755),
            .I(N__36383));
    SRMux I__8817 (
            .O(N__36754),
            .I(N__36383));
    SRMux I__8816 (
            .O(N__36753),
            .I(N__36383));
    SRMux I__8815 (
            .O(N__36752),
            .I(N__36383));
    SRMux I__8814 (
            .O(N__36751),
            .I(N__36383));
    SRMux I__8813 (
            .O(N__36750),
            .I(N__36383));
    SRMux I__8812 (
            .O(N__36749),
            .I(N__36383));
    SRMux I__8811 (
            .O(N__36748),
            .I(N__36383));
    SRMux I__8810 (
            .O(N__36747),
            .I(N__36383));
    SRMux I__8809 (
            .O(N__36746),
            .I(N__36383));
    SRMux I__8808 (
            .O(N__36745),
            .I(N__36383));
    SRMux I__8807 (
            .O(N__36744),
            .I(N__36383));
    SRMux I__8806 (
            .O(N__36743),
            .I(N__36383));
    SRMux I__8805 (
            .O(N__36742),
            .I(N__36383));
    SRMux I__8804 (
            .O(N__36741),
            .I(N__36383));
    SRMux I__8803 (
            .O(N__36740),
            .I(N__36383));
    SRMux I__8802 (
            .O(N__36739),
            .I(N__36383));
    SRMux I__8801 (
            .O(N__36738),
            .I(N__36383));
    SRMux I__8800 (
            .O(N__36737),
            .I(N__36383));
    SRMux I__8799 (
            .O(N__36736),
            .I(N__36383));
    SRMux I__8798 (
            .O(N__36735),
            .I(N__36383));
    SRMux I__8797 (
            .O(N__36734),
            .I(N__36383));
    SRMux I__8796 (
            .O(N__36733),
            .I(N__36383));
    SRMux I__8795 (
            .O(N__36732),
            .I(N__36383));
    SRMux I__8794 (
            .O(N__36731),
            .I(N__36383));
    SRMux I__8793 (
            .O(N__36730),
            .I(N__36383));
    SRMux I__8792 (
            .O(N__36729),
            .I(N__36383));
    SRMux I__8791 (
            .O(N__36728),
            .I(N__36383));
    SRMux I__8790 (
            .O(N__36727),
            .I(N__36383));
    SRMux I__8789 (
            .O(N__36726),
            .I(N__36383));
    SRMux I__8788 (
            .O(N__36725),
            .I(N__36383));
    SRMux I__8787 (
            .O(N__36724),
            .I(N__36383));
    SRMux I__8786 (
            .O(N__36723),
            .I(N__36383));
    SRMux I__8785 (
            .O(N__36722),
            .I(N__36383));
    SRMux I__8784 (
            .O(N__36721),
            .I(N__36383));
    SRMux I__8783 (
            .O(N__36720),
            .I(N__36383));
    SRMux I__8782 (
            .O(N__36719),
            .I(N__36383));
    SRMux I__8781 (
            .O(N__36718),
            .I(N__36383));
    SRMux I__8780 (
            .O(N__36717),
            .I(N__36383));
    SRMux I__8779 (
            .O(N__36716),
            .I(N__36383));
    SRMux I__8778 (
            .O(N__36715),
            .I(N__36383));
    SRMux I__8777 (
            .O(N__36714),
            .I(N__36383));
    SRMux I__8776 (
            .O(N__36713),
            .I(N__36383));
    SRMux I__8775 (
            .O(N__36712),
            .I(N__36383));
    SRMux I__8774 (
            .O(N__36711),
            .I(N__36383));
    SRMux I__8773 (
            .O(N__36710),
            .I(N__36383));
    SRMux I__8772 (
            .O(N__36709),
            .I(N__36383));
    SRMux I__8771 (
            .O(N__36708),
            .I(N__36383));
    SRMux I__8770 (
            .O(N__36707),
            .I(N__36383));
    SRMux I__8769 (
            .O(N__36706),
            .I(N__36383));
    SRMux I__8768 (
            .O(N__36705),
            .I(N__36383));
    SRMux I__8767 (
            .O(N__36704),
            .I(N__36383));
    SRMux I__8766 (
            .O(N__36703),
            .I(N__36383));
    SRMux I__8765 (
            .O(N__36702),
            .I(N__36383));
    SRMux I__8764 (
            .O(N__36701),
            .I(N__36383));
    SRMux I__8763 (
            .O(N__36700),
            .I(N__36383));
    SRMux I__8762 (
            .O(N__36699),
            .I(N__36383));
    SRMux I__8761 (
            .O(N__36698),
            .I(N__36383));
    SRMux I__8760 (
            .O(N__36697),
            .I(N__36383));
    SRMux I__8759 (
            .O(N__36696),
            .I(N__36383));
    SRMux I__8758 (
            .O(N__36695),
            .I(N__36383));
    SRMux I__8757 (
            .O(N__36694),
            .I(N__36383));
    SRMux I__8756 (
            .O(N__36693),
            .I(N__36383));
    SRMux I__8755 (
            .O(N__36692),
            .I(N__36383));
    SRMux I__8754 (
            .O(N__36691),
            .I(N__36383));
    SRMux I__8753 (
            .O(N__36690),
            .I(N__36383));
    SRMux I__8752 (
            .O(N__36689),
            .I(N__36383));
    Glb2LocalMux I__8751 (
            .O(N__36686),
            .I(N__36383));
    Glb2LocalMux I__8750 (
            .O(N__36683),
            .I(N__36383));
    Glb2LocalMux I__8749 (
            .O(N__36680),
            .I(N__36383));
    Glb2LocalMux I__8748 (
            .O(N__36677),
            .I(N__36383));
    Glb2LocalMux I__8747 (
            .O(N__36674),
            .I(N__36383));
    Glb2LocalMux I__8746 (
            .O(N__36671),
            .I(N__36383));
    Glb2LocalMux I__8745 (
            .O(N__36668),
            .I(N__36383));
    Glb2LocalMux I__8744 (
            .O(N__36665),
            .I(N__36383));
    Glb2LocalMux I__8743 (
            .O(N__36662),
            .I(N__36383));
    Glb2LocalMux I__8742 (
            .O(N__36659),
            .I(N__36383));
    Glb2LocalMux I__8741 (
            .O(N__36656),
            .I(N__36383));
    Glb2LocalMux I__8740 (
            .O(N__36653),
            .I(N__36383));
    Glb2LocalMux I__8739 (
            .O(N__36650),
            .I(N__36383));
    Glb2LocalMux I__8738 (
            .O(N__36647),
            .I(N__36383));
    Glb2LocalMux I__8737 (
            .O(N__36644),
            .I(N__36383));
    Glb2LocalMux I__8736 (
            .O(N__36641),
            .I(N__36383));
    Glb2LocalMux I__8735 (
            .O(N__36638),
            .I(N__36383));
    Glb2LocalMux I__8734 (
            .O(N__36635),
            .I(N__36383));
    Glb2LocalMux I__8733 (
            .O(N__36632),
            .I(N__36383));
    Glb2LocalMux I__8732 (
            .O(N__36629),
            .I(N__36383));
    Glb2LocalMux I__8731 (
            .O(N__36626),
            .I(N__36383));
    Glb2LocalMux I__8730 (
            .O(N__36623),
            .I(N__36383));
    Glb2LocalMux I__8729 (
            .O(N__36620),
            .I(N__36383));
    Glb2LocalMux I__8728 (
            .O(N__36617),
            .I(N__36383));
    Glb2LocalMux I__8727 (
            .O(N__36614),
            .I(N__36383));
    Glb2LocalMux I__8726 (
            .O(N__36611),
            .I(N__36383));
    Glb2LocalMux I__8725 (
            .O(N__36608),
            .I(N__36383));
    GlobalMux I__8724 (
            .O(N__36383),
            .I(N__36380));
    gio2CtrlBuf I__8723 (
            .O(N__36380),
            .I(reset_system_g));
    IoInMux I__8722 (
            .O(N__36377),
            .I(N__36374));
    LocalMux I__8721 (
            .O(N__36374),
            .I(N__36371));
    Odrv12 I__8720 (
            .O(N__36371),
            .I(debug_CH3_20A_c_0));
    InMux I__8719 (
            .O(N__36368),
            .I(N__36365));
    LocalMux I__8718 (
            .O(N__36365),
            .I(N__36362));
    Span4Mux_h I__8717 (
            .O(N__36362),
            .I(N__36359));
    Odrv4 I__8716 (
            .O(N__36359),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__8715 (
            .O(N__36356),
            .I(N__36353));
    InMux I__8714 (
            .O(N__36353),
            .I(N__36346));
    InMux I__8713 (
            .O(N__36352),
            .I(N__36346));
    InMux I__8712 (
            .O(N__36351),
            .I(N__36340));
    LocalMux I__8711 (
            .O(N__36346),
            .I(N__36335));
    InMux I__8710 (
            .O(N__36345),
            .I(N__36332));
    InMux I__8709 (
            .O(N__36344),
            .I(N__36329));
    InMux I__8708 (
            .O(N__36343),
            .I(N__36321));
    LocalMux I__8707 (
            .O(N__36340),
            .I(N__36318));
    InMux I__8706 (
            .O(N__36339),
            .I(N__36315));
    IoInMux I__8705 (
            .O(N__36338),
            .I(N__36311));
    Span4Mux_h I__8704 (
            .O(N__36335),
            .I(N__36308));
    LocalMux I__8703 (
            .O(N__36332),
            .I(N__36303));
    LocalMux I__8702 (
            .O(N__36329),
            .I(N__36303));
    InMux I__8701 (
            .O(N__36328),
            .I(N__36294));
    InMux I__8700 (
            .O(N__36327),
            .I(N__36294));
    InMux I__8699 (
            .O(N__36326),
            .I(N__36294));
    InMux I__8698 (
            .O(N__36325),
            .I(N__36294));
    InMux I__8697 (
            .O(N__36324),
            .I(N__36291));
    LocalMux I__8696 (
            .O(N__36321),
            .I(N__36284));
    Span4Mux_v I__8695 (
            .O(N__36318),
            .I(N__36284));
    LocalMux I__8694 (
            .O(N__36315),
            .I(N__36284));
    InMux I__8693 (
            .O(N__36314),
            .I(N__36281));
    LocalMux I__8692 (
            .O(N__36311),
            .I(N__36278));
    Span4Mux_v I__8691 (
            .O(N__36308),
            .I(N__36275));
    Span4Mux_h I__8690 (
            .O(N__36303),
            .I(N__36270));
    LocalMux I__8689 (
            .O(N__36294),
            .I(N__36270));
    LocalMux I__8688 (
            .O(N__36291),
            .I(N__36263));
    Span4Mux_h I__8687 (
            .O(N__36284),
            .I(N__36263));
    LocalMux I__8686 (
            .O(N__36281),
            .I(N__36263));
    Span4Mux_s1_v I__8685 (
            .O(N__36278),
            .I(N__36260));
    Sp12to4 I__8684 (
            .O(N__36275),
            .I(N__36255));
    Sp12to4 I__8683 (
            .O(N__36270),
            .I(N__36255));
    Sp12to4 I__8682 (
            .O(N__36263),
            .I(N__36252));
    Span4Mux_h I__8681 (
            .O(N__36260),
            .I(N__36249));
    Span12Mux_v I__8680 (
            .O(N__36255),
            .I(N__36246));
    Span12Mux_v I__8679 (
            .O(N__36252),
            .I(N__36243));
    Odrv4 I__8678 (
            .O(N__36249),
            .I(debug_CH2_18A_c));
    Odrv12 I__8677 (
            .O(N__36246),
            .I(debug_CH2_18A_c));
    Odrv12 I__8676 (
            .O(N__36243),
            .I(debug_CH2_18A_c));
    InMux I__8675 (
            .O(N__36236),
            .I(N__36231));
    InMux I__8674 (
            .O(N__36235),
            .I(N__36225));
    InMux I__8673 (
            .O(N__36234),
            .I(N__36225));
    LocalMux I__8672 (
            .O(N__36231),
            .I(N__36222));
    InMux I__8671 (
            .O(N__36230),
            .I(N__36219));
    LocalMux I__8670 (
            .O(N__36225),
            .I(N__36213));
    Span4Mux_h I__8669 (
            .O(N__36222),
            .I(N__36208));
    LocalMux I__8668 (
            .O(N__36219),
            .I(N__36208));
    InMux I__8667 (
            .O(N__36218),
            .I(N__36201));
    InMux I__8666 (
            .O(N__36217),
            .I(N__36201));
    InMux I__8665 (
            .O(N__36216),
            .I(N__36201));
    Odrv4 I__8664 (
            .O(N__36213),
            .I(\uart_pc.un1_state_2_0 ));
    Odrv4 I__8663 (
            .O(N__36208),
            .I(\uart_pc.un1_state_2_0 ));
    LocalMux I__8662 (
            .O(N__36201),
            .I(\uart_pc.un1_state_2_0 ));
    CascadeMux I__8661 (
            .O(N__36194),
            .I(N__36191));
    InMux I__8660 (
            .O(N__36191),
            .I(N__36188));
    LocalMux I__8659 (
            .O(N__36188),
            .I(N__36185));
    Span4Mux_h I__8658 (
            .O(N__36185),
            .I(N__36181));
    CascadeMux I__8657 (
            .O(N__36184),
            .I(N__36178));
    Span4Mux_h I__8656 (
            .O(N__36181),
            .I(N__36175));
    InMux I__8655 (
            .O(N__36178),
            .I(N__36172));
    Odrv4 I__8654 (
            .O(N__36175),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__8653 (
            .O(N__36172),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    ClkMux I__8652 (
            .O(N__36167),
            .I(N__35690));
    ClkMux I__8651 (
            .O(N__36166),
            .I(N__35690));
    ClkMux I__8650 (
            .O(N__36165),
            .I(N__35690));
    ClkMux I__8649 (
            .O(N__36164),
            .I(N__35690));
    ClkMux I__8648 (
            .O(N__36163),
            .I(N__35690));
    ClkMux I__8647 (
            .O(N__36162),
            .I(N__35690));
    ClkMux I__8646 (
            .O(N__36161),
            .I(N__35690));
    ClkMux I__8645 (
            .O(N__36160),
            .I(N__35690));
    ClkMux I__8644 (
            .O(N__36159),
            .I(N__35690));
    ClkMux I__8643 (
            .O(N__36158),
            .I(N__35690));
    ClkMux I__8642 (
            .O(N__36157),
            .I(N__35690));
    ClkMux I__8641 (
            .O(N__36156),
            .I(N__35690));
    ClkMux I__8640 (
            .O(N__36155),
            .I(N__35690));
    ClkMux I__8639 (
            .O(N__36154),
            .I(N__35690));
    ClkMux I__8638 (
            .O(N__36153),
            .I(N__35690));
    ClkMux I__8637 (
            .O(N__36152),
            .I(N__35690));
    ClkMux I__8636 (
            .O(N__36151),
            .I(N__35690));
    ClkMux I__8635 (
            .O(N__36150),
            .I(N__35690));
    ClkMux I__8634 (
            .O(N__36149),
            .I(N__35690));
    ClkMux I__8633 (
            .O(N__36148),
            .I(N__35690));
    ClkMux I__8632 (
            .O(N__36147),
            .I(N__35690));
    ClkMux I__8631 (
            .O(N__36146),
            .I(N__35690));
    ClkMux I__8630 (
            .O(N__36145),
            .I(N__35690));
    ClkMux I__8629 (
            .O(N__36144),
            .I(N__35690));
    ClkMux I__8628 (
            .O(N__36143),
            .I(N__35690));
    ClkMux I__8627 (
            .O(N__36142),
            .I(N__35690));
    ClkMux I__8626 (
            .O(N__36141),
            .I(N__35690));
    ClkMux I__8625 (
            .O(N__36140),
            .I(N__35690));
    ClkMux I__8624 (
            .O(N__36139),
            .I(N__35690));
    ClkMux I__8623 (
            .O(N__36138),
            .I(N__35690));
    ClkMux I__8622 (
            .O(N__36137),
            .I(N__35690));
    ClkMux I__8621 (
            .O(N__36136),
            .I(N__35690));
    ClkMux I__8620 (
            .O(N__36135),
            .I(N__35690));
    ClkMux I__8619 (
            .O(N__36134),
            .I(N__35690));
    ClkMux I__8618 (
            .O(N__36133),
            .I(N__35690));
    ClkMux I__8617 (
            .O(N__36132),
            .I(N__35690));
    ClkMux I__8616 (
            .O(N__36131),
            .I(N__35690));
    ClkMux I__8615 (
            .O(N__36130),
            .I(N__35690));
    ClkMux I__8614 (
            .O(N__36129),
            .I(N__35690));
    ClkMux I__8613 (
            .O(N__36128),
            .I(N__35690));
    ClkMux I__8612 (
            .O(N__36127),
            .I(N__35690));
    ClkMux I__8611 (
            .O(N__36126),
            .I(N__35690));
    ClkMux I__8610 (
            .O(N__36125),
            .I(N__35690));
    ClkMux I__8609 (
            .O(N__36124),
            .I(N__35690));
    ClkMux I__8608 (
            .O(N__36123),
            .I(N__35690));
    ClkMux I__8607 (
            .O(N__36122),
            .I(N__35690));
    ClkMux I__8606 (
            .O(N__36121),
            .I(N__35690));
    ClkMux I__8605 (
            .O(N__36120),
            .I(N__35690));
    ClkMux I__8604 (
            .O(N__36119),
            .I(N__35690));
    ClkMux I__8603 (
            .O(N__36118),
            .I(N__35690));
    ClkMux I__8602 (
            .O(N__36117),
            .I(N__35690));
    ClkMux I__8601 (
            .O(N__36116),
            .I(N__35690));
    ClkMux I__8600 (
            .O(N__36115),
            .I(N__35690));
    ClkMux I__8599 (
            .O(N__36114),
            .I(N__35690));
    ClkMux I__8598 (
            .O(N__36113),
            .I(N__35690));
    ClkMux I__8597 (
            .O(N__36112),
            .I(N__35690));
    ClkMux I__8596 (
            .O(N__36111),
            .I(N__35690));
    ClkMux I__8595 (
            .O(N__36110),
            .I(N__35690));
    ClkMux I__8594 (
            .O(N__36109),
            .I(N__35690));
    ClkMux I__8593 (
            .O(N__36108),
            .I(N__35690));
    ClkMux I__8592 (
            .O(N__36107),
            .I(N__35690));
    ClkMux I__8591 (
            .O(N__36106),
            .I(N__35690));
    ClkMux I__8590 (
            .O(N__36105),
            .I(N__35690));
    ClkMux I__8589 (
            .O(N__36104),
            .I(N__35690));
    ClkMux I__8588 (
            .O(N__36103),
            .I(N__35690));
    ClkMux I__8587 (
            .O(N__36102),
            .I(N__35690));
    ClkMux I__8586 (
            .O(N__36101),
            .I(N__35690));
    ClkMux I__8585 (
            .O(N__36100),
            .I(N__35690));
    ClkMux I__8584 (
            .O(N__36099),
            .I(N__35690));
    ClkMux I__8583 (
            .O(N__36098),
            .I(N__35690));
    ClkMux I__8582 (
            .O(N__36097),
            .I(N__35690));
    ClkMux I__8581 (
            .O(N__36096),
            .I(N__35690));
    ClkMux I__8580 (
            .O(N__36095),
            .I(N__35690));
    ClkMux I__8579 (
            .O(N__36094),
            .I(N__35690));
    ClkMux I__8578 (
            .O(N__36093),
            .I(N__35690));
    ClkMux I__8577 (
            .O(N__36092),
            .I(N__35690));
    ClkMux I__8576 (
            .O(N__36091),
            .I(N__35690));
    ClkMux I__8575 (
            .O(N__36090),
            .I(N__35690));
    ClkMux I__8574 (
            .O(N__36089),
            .I(N__35690));
    ClkMux I__8573 (
            .O(N__36088),
            .I(N__35690));
    ClkMux I__8572 (
            .O(N__36087),
            .I(N__35690));
    ClkMux I__8571 (
            .O(N__36086),
            .I(N__35690));
    ClkMux I__8570 (
            .O(N__36085),
            .I(N__35690));
    ClkMux I__8569 (
            .O(N__36084),
            .I(N__35690));
    ClkMux I__8568 (
            .O(N__36083),
            .I(N__35690));
    ClkMux I__8567 (
            .O(N__36082),
            .I(N__35690));
    ClkMux I__8566 (
            .O(N__36081),
            .I(N__35690));
    ClkMux I__8565 (
            .O(N__36080),
            .I(N__35690));
    ClkMux I__8564 (
            .O(N__36079),
            .I(N__35690));
    ClkMux I__8563 (
            .O(N__36078),
            .I(N__35690));
    ClkMux I__8562 (
            .O(N__36077),
            .I(N__35690));
    ClkMux I__8561 (
            .O(N__36076),
            .I(N__35690));
    ClkMux I__8560 (
            .O(N__36075),
            .I(N__35690));
    ClkMux I__8559 (
            .O(N__36074),
            .I(N__35690));
    ClkMux I__8558 (
            .O(N__36073),
            .I(N__35690));
    ClkMux I__8557 (
            .O(N__36072),
            .I(N__35690));
    ClkMux I__8556 (
            .O(N__36071),
            .I(N__35690));
    ClkMux I__8555 (
            .O(N__36070),
            .I(N__35690));
    ClkMux I__8554 (
            .O(N__36069),
            .I(N__35690));
    ClkMux I__8553 (
            .O(N__36068),
            .I(N__35690));
    ClkMux I__8552 (
            .O(N__36067),
            .I(N__35690));
    ClkMux I__8551 (
            .O(N__36066),
            .I(N__35690));
    ClkMux I__8550 (
            .O(N__36065),
            .I(N__35690));
    ClkMux I__8549 (
            .O(N__36064),
            .I(N__35690));
    ClkMux I__8548 (
            .O(N__36063),
            .I(N__35690));
    ClkMux I__8547 (
            .O(N__36062),
            .I(N__35690));
    ClkMux I__8546 (
            .O(N__36061),
            .I(N__35690));
    ClkMux I__8545 (
            .O(N__36060),
            .I(N__35690));
    ClkMux I__8544 (
            .O(N__36059),
            .I(N__35690));
    ClkMux I__8543 (
            .O(N__36058),
            .I(N__35690));
    ClkMux I__8542 (
            .O(N__36057),
            .I(N__35690));
    ClkMux I__8541 (
            .O(N__36056),
            .I(N__35690));
    ClkMux I__8540 (
            .O(N__36055),
            .I(N__35690));
    ClkMux I__8539 (
            .O(N__36054),
            .I(N__35690));
    ClkMux I__8538 (
            .O(N__36053),
            .I(N__35690));
    ClkMux I__8537 (
            .O(N__36052),
            .I(N__35690));
    ClkMux I__8536 (
            .O(N__36051),
            .I(N__35690));
    ClkMux I__8535 (
            .O(N__36050),
            .I(N__35690));
    ClkMux I__8534 (
            .O(N__36049),
            .I(N__35690));
    ClkMux I__8533 (
            .O(N__36048),
            .I(N__35690));
    ClkMux I__8532 (
            .O(N__36047),
            .I(N__35690));
    ClkMux I__8531 (
            .O(N__36046),
            .I(N__35690));
    ClkMux I__8530 (
            .O(N__36045),
            .I(N__35690));
    ClkMux I__8529 (
            .O(N__36044),
            .I(N__35690));
    ClkMux I__8528 (
            .O(N__36043),
            .I(N__35690));
    ClkMux I__8527 (
            .O(N__36042),
            .I(N__35690));
    ClkMux I__8526 (
            .O(N__36041),
            .I(N__35690));
    ClkMux I__8525 (
            .O(N__36040),
            .I(N__35690));
    ClkMux I__8524 (
            .O(N__36039),
            .I(N__35690));
    ClkMux I__8523 (
            .O(N__36038),
            .I(N__35690));
    ClkMux I__8522 (
            .O(N__36037),
            .I(N__35690));
    ClkMux I__8521 (
            .O(N__36036),
            .I(N__35690));
    ClkMux I__8520 (
            .O(N__36035),
            .I(N__35690));
    ClkMux I__8519 (
            .O(N__36034),
            .I(N__35690));
    ClkMux I__8518 (
            .O(N__36033),
            .I(N__35690));
    ClkMux I__8517 (
            .O(N__36032),
            .I(N__35690));
    ClkMux I__8516 (
            .O(N__36031),
            .I(N__35690));
    ClkMux I__8515 (
            .O(N__36030),
            .I(N__35690));
    ClkMux I__8514 (
            .O(N__36029),
            .I(N__35690));
    ClkMux I__8513 (
            .O(N__36028),
            .I(N__35690));
    ClkMux I__8512 (
            .O(N__36027),
            .I(N__35690));
    ClkMux I__8511 (
            .O(N__36026),
            .I(N__35690));
    ClkMux I__8510 (
            .O(N__36025),
            .I(N__35690));
    ClkMux I__8509 (
            .O(N__36024),
            .I(N__35690));
    ClkMux I__8508 (
            .O(N__36023),
            .I(N__35690));
    ClkMux I__8507 (
            .O(N__36022),
            .I(N__35690));
    ClkMux I__8506 (
            .O(N__36021),
            .I(N__35690));
    ClkMux I__8505 (
            .O(N__36020),
            .I(N__35690));
    ClkMux I__8504 (
            .O(N__36019),
            .I(N__35690));
    ClkMux I__8503 (
            .O(N__36018),
            .I(N__35690));
    ClkMux I__8502 (
            .O(N__36017),
            .I(N__35690));
    ClkMux I__8501 (
            .O(N__36016),
            .I(N__35690));
    ClkMux I__8500 (
            .O(N__36015),
            .I(N__35690));
    ClkMux I__8499 (
            .O(N__36014),
            .I(N__35690));
    ClkMux I__8498 (
            .O(N__36013),
            .I(N__35690));
    ClkMux I__8497 (
            .O(N__36012),
            .I(N__35690));
    ClkMux I__8496 (
            .O(N__36011),
            .I(N__35690));
    ClkMux I__8495 (
            .O(N__36010),
            .I(N__35690));
    ClkMux I__8494 (
            .O(N__36009),
            .I(N__35690));
    GlobalMux I__8493 (
            .O(N__35690),
            .I(N__35687));
    gio2CtrlBuf I__8492 (
            .O(N__35687),
            .I(clk_system_c_g));
    SRMux I__8491 (
            .O(N__35684),
            .I(N__35680));
    SRMux I__8490 (
            .O(N__35683),
            .I(N__35676));
    LocalMux I__8489 (
            .O(N__35680),
            .I(N__35672));
    SRMux I__8488 (
            .O(N__35679),
            .I(N__35669));
    LocalMux I__8487 (
            .O(N__35676),
            .I(N__35666));
    SRMux I__8486 (
            .O(N__35675),
            .I(N__35663));
    Span4Mux_h I__8485 (
            .O(N__35672),
            .I(N__35660));
    LocalMux I__8484 (
            .O(N__35669),
            .I(N__35657));
    Span4Mux_v I__8483 (
            .O(N__35666),
            .I(N__35652));
    LocalMux I__8482 (
            .O(N__35663),
            .I(N__35652));
    Odrv4 I__8481 (
            .O(N__35660),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv12 I__8480 (
            .O(N__35657),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv4 I__8479 (
            .O(N__35652),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__8478 (
            .O(N__35645),
            .I(N__35641));
    InMux I__8477 (
            .O(N__35644),
            .I(N__35638));
    LocalMux I__8476 (
            .O(N__35641),
            .I(N__35635));
    LocalMux I__8475 (
            .O(N__35638),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__8474 (
            .O(N__35635),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__8473 (
            .O(N__35630),
            .I(N__35626));
    InMux I__8472 (
            .O(N__35629),
            .I(N__35623));
    LocalMux I__8471 (
            .O(N__35626),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__8470 (
            .O(N__35623),
            .I(\reset_module_System.countZ0Z_16 ));
    CascadeMux I__8469 (
            .O(N__35618),
            .I(\reset_module_System.reset6_3_cascade_ ));
    InMux I__8468 (
            .O(N__35615),
            .I(N__35612));
    LocalMux I__8467 (
            .O(N__35612),
            .I(\reset_module_System.reset6_13 ));
    InMux I__8466 (
            .O(N__35609),
            .I(N__35606));
    LocalMux I__8465 (
            .O(N__35606),
            .I(N__35602));
    InMux I__8464 (
            .O(N__35605),
            .I(N__35599));
    Odrv4 I__8463 (
            .O(N__35602),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__8462 (
            .O(N__35599),
            .I(\reset_module_System.countZ0Z_12 ));
    CascadeMux I__8461 (
            .O(N__35594),
            .I(\reset_module_System.reset6_17_cascade_ ));
    CascadeMux I__8460 (
            .O(N__35591),
            .I(\reset_module_System.reset6_19_cascade_ ));
    CascadeMux I__8459 (
            .O(N__35588),
            .I(N__35582));
    InMux I__8458 (
            .O(N__35587),
            .I(N__35575));
    InMux I__8457 (
            .O(N__35586),
            .I(N__35575));
    InMux I__8456 (
            .O(N__35585),
            .I(N__35575));
    InMux I__8455 (
            .O(N__35582),
            .I(N__35572));
    LocalMux I__8454 (
            .O(N__35575),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__8453 (
            .O(N__35572),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__8452 (
            .O(N__35567),
            .I(N__35560));
    InMux I__8451 (
            .O(N__35566),
            .I(N__35560));
    InMux I__8450 (
            .O(N__35565),
            .I(N__35557));
    LocalMux I__8449 (
            .O(N__35560),
            .I(\reset_module_System.reset6_15 ));
    LocalMux I__8448 (
            .O(N__35557),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__8447 (
            .O(N__35552),
            .I(\reset_module_System.count_1_1_cascade_ ));
    InMux I__8446 (
            .O(N__35549),
            .I(N__35544));
    InMux I__8445 (
            .O(N__35548),
            .I(N__35539));
    InMux I__8444 (
            .O(N__35547),
            .I(N__35539));
    LocalMux I__8443 (
            .O(N__35544),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__8442 (
            .O(N__35539),
            .I(\reset_module_System.reset6_19 ));
    InMux I__8441 (
            .O(N__35534),
            .I(N__35529));
    InMux I__8440 (
            .O(N__35533),
            .I(N__35524));
    InMux I__8439 (
            .O(N__35532),
            .I(N__35524));
    LocalMux I__8438 (
            .O(N__35529),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__8437 (
            .O(N__35524),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__8436 (
            .O(N__35519),
            .I(N__35515));
    InMux I__8435 (
            .O(N__35518),
            .I(N__35512));
    LocalMux I__8434 (
            .O(N__35515),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__8433 (
            .O(N__35512),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__8432 (
            .O(N__35507),
            .I(N__35503));
    InMux I__8431 (
            .O(N__35506),
            .I(N__35500));
    LocalMux I__8430 (
            .O(N__35503),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__8429 (
            .O(N__35500),
            .I(\reset_module_System.countZ0Z_11 ));
    CascadeMux I__8428 (
            .O(N__35495),
            .I(N__35492));
    InMux I__8427 (
            .O(N__35492),
            .I(N__35488));
    InMux I__8426 (
            .O(N__35491),
            .I(N__35485));
    LocalMux I__8425 (
            .O(N__35488),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__8424 (
            .O(N__35485),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__8423 (
            .O(N__35480),
            .I(N__35476));
    InMux I__8422 (
            .O(N__35479),
            .I(N__35473));
    LocalMux I__8421 (
            .O(N__35476),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__8420 (
            .O(N__35473),
            .I(\reset_module_System.countZ0Z_10 ));
    CascadeMux I__8419 (
            .O(N__35468),
            .I(N__35465));
    InMux I__8418 (
            .O(N__35465),
            .I(N__35457));
    InMux I__8417 (
            .O(N__35464),
            .I(N__35457));
    InMux I__8416 (
            .O(N__35463),
            .I(N__35454));
    InMux I__8415 (
            .O(N__35462),
            .I(N__35451));
    LocalMux I__8414 (
            .O(N__35457),
            .I(N__35448));
    LocalMux I__8413 (
            .O(N__35454),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__8412 (
            .O(N__35451),
            .I(\reset_module_System.reset6_14 ));
    Odrv4 I__8411 (
            .O(N__35448),
            .I(\reset_module_System.reset6_14 ));
    InMux I__8410 (
            .O(N__35441),
            .I(N__35437));
    InMux I__8409 (
            .O(N__35440),
            .I(N__35434));
    LocalMux I__8408 (
            .O(N__35437),
            .I(\reset_module_System.countZ0Z_19 ));
    LocalMux I__8407 (
            .O(N__35434),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__8406 (
            .O(N__35429),
            .I(N__35425));
    InMux I__8405 (
            .O(N__35428),
            .I(N__35422));
    LocalMux I__8404 (
            .O(N__35425),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__8403 (
            .O(N__35422),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__8402 (
            .O(N__35417),
            .I(N__35413));
    InMux I__8401 (
            .O(N__35416),
            .I(N__35410));
    InMux I__8400 (
            .O(N__35413),
            .I(N__35407));
    LocalMux I__8399 (
            .O(N__35410),
            .I(\reset_module_System.countZ0Z_21 ));
    LocalMux I__8398 (
            .O(N__35407),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__8397 (
            .O(N__35402),
            .I(N__35398));
    InMux I__8396 (
            .O(N__35401),
            .I(N__35395));
    LocalMux I__8395 (
            .O(N__35398),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__8394 (
            .O(N__35395),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__8393 (
            .O(N__35390),
            .I(N__35387));
    LocalMux I__8392 (
            .O(N__35387),
            .I(\reset_module_System.reset6_11 ));
    InMux I__8391 (
            .O(N__35384),
            .I(N__35381));
    LocalMux I__8390 (
            .O(N__35381),
            .I(N__35378));
    Span4Mux_h I__8389 (
            .O(N__35378),
            .I(N__35375));
    Odrv4 I__8388 (
            .O(N__35375),
            .I(\uart_pc.data_Auxce_0_3 ));
    CascadeMux I__8387 (
            .O(N__35372),
            .I(N__35369));
    InMux I__8386 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__8385 (
            .O(N__35366),
            .I(N__35362));
    CascadeMux I__8384 (
            .O(N__35365),
            .I(N__35359));
    Span4Mux_h I__8383 (
            .O(N__35362),
            .I(N__35356));
    InMux I__8382 (
            .O(N__35359),
            .I(N__35353));
    Odrv4 I__8381 (
            .O(N__35356),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__8380 (
            .O(N__35353),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__8379 (
            .O(N__35348),
            .I(N__35345));
    LocalMux I__8378 (
            .O(N__35345),
            .I(N__35341));
    InMux I__8377 (
            .O(N__35344),
            .I(N__35338));
    Span4Mux_h I__8376 (
            .O(N__35341),
            .I(N__35332));
    LocalMux I__8375 (
            .O(N__35338),
            .I(N__35332));
    InMux I__8374 (
            .O(N__35337),
            .I(N__35329));
    Sp12to4 I__8373 (
            .O(N__35332),
            .I(N__35319));
    LocalMux I__8372 (
            .O(N__35329),
            .I(N__35319));
    InMux I__8371 (
            .O(N__35328),
            .I(N__35314));
    InMux I__8370 (
            .O(N__35327),
            .I(N__35314));
    InMux I__8369 (
            .O(N__35326),
            .I(N__35309));
    InMux I__8368 (
            .O(N__35325),
            .I(N__35309));
    InMux I__8367 (
            .O(N__35324),
            .I(N__35306));
    Odrv12 I__8366 (
            .O(N__35319),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__8365 (
            .O(N__35314),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__8364 (
            .O(N__35309),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__8363 (
            .O(N__35306),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__8362 (
            .O(N__35297),
            .I(N__35294));
    LocalMux I__8361 (
            .O(N__35294),
            .I(N__35289));
    InMux I__8360 (
            .O(N__35293),
            .I(N__35284));
    InMux I__8359 (
            .O(N__35292),
            .I(N__35284));
    Span4Mux_h I__8358 (
            .O(N__35289),
            .I(N__35279));
    LocalMux I__8357 (
            .O(N__35284),
            .I(N__35279));
    Odrv4 I__8356 (
            .O(N__35279),
            .I(\uart_pc.N_126_li ));
    InMux I__8355 (
            .O(N__35276),
            .I(N__35273));
    LocalMux I__8354 (
            .O(N__35273),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    InMux I__8353 (
            .O(N__35270),
            .I(N__35265));
    InMux I__8352 (
            .O(N__35269),
            .I(N__35260));
    InMux I__8351 (
            .O(N__35268),
            .I(N__35257));
    LocalMux I__8350 (
            .O(N__35265),
            .I(N__35253));
    CascadeMux I__8349 (
            .O(N__35264),
            .I(N__35250));
    CascadeMux I__8348 (
            .O(N__35263),
            .I(N__35247));
    LocalMux I__8347 (
            .O(N__35260),
            .I(N__35241));
    LocalMux I__8346 (
            .O(N__35257),
            .I(N__35241));
    CascadeMux I__8345 (
            .O(N__35256),
            .I(N__35237));
    Span4Mux_h I__8344 (
            .O(N__35253),
            .I(N__35233));
    InMux I__8343 (
            .O(N__35250),
            .I(N__35228));
    InMux I__8342 (
            .O(N__35247),
            .I(N__35228));
    CascadeMux I__8341 (
            .O(N__35246),
            .I(N__35225));
    Span4Mux_h I__8340 (
            .O(N__35241),
            .I(N__35222));
    InMux I__8339 (
            .O(N__35240),
            .I(N__35217));
    InMux I__8338 (
            .O(N__35237),
            .I(N__35217));
    InMux I__8337 (
            .O(N__35236),
            .I(N__35214));
    Span4Mux_v I__8336 (
            .O(N__35233),
            .I(N__35209));
    LocalMux I__8335 (
            .O(N__35228),
            .I(N__35209));
    InMux I__8334 (
            .O(N__35225),
            .I(N__35206));
    Odrv4 I__8333 (
            .O(N__35222),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__8332 (
            .O(N__35217),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__8331 (
            .O(N__35214),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__8330 (
            .O(N__35209),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__8329 (
            .O(N__35206),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__8328 (
            .O(N__35195),
            .I(N__35192));
    LocalMux I__8327 (
            .O(N__35192),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    CascadeMux I__8326 (
            .O(N__35189),
            .I(N__35186));
    InMux I__8325 (
            .O(N__35186),
            .I(N__35179));
    InMux I__8324 (
            .O(N__35185),
            .I(N__35179));
    InMux I__8323 (
            .O(N__35184),
            .I(N__35176));
    LocalMux I__8322 (
            .O(N__35179),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__8321 (
            .O(N__35176),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    CascadeMux I__8320 (
            .O(N__35171),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ));
    InMux I__8319 (
            .O(N__35168),
            .I(N__35164));
    InMux I__8318 (
            .O(N__35167),
            .I(N__35161));
    LocalMux I__8317 (
            .O(N__35164),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__8316 (
            .O(N__35161),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    CascadeMux I__8315 (
            .O(N__35156),
            .I(N__35149));
    CascadeMux I__8314 (
            .O(N__35155),
            .I(N__35146));
    InMux I__8313 (
            .O(N__35154),
            .I(N__35140));
    InMux I__8312 (
            .O(N__35153),
            .I(N__35140));
    InMux I__8311 (
            .O(N__35152),
            .I(N__35135));
    InMux I__8310 (
            .O(N__35149),
            .I(N__35135));
    InMux I__8309 (
            .O(N__35146),
            .I(N__35130));
    InMux I__8308 (
            .O(N__35145),
            .I(N__35130));
    LocalMux I__8307 (
            .O(N__35140),
            .I(N__35127));
    LocalMux I__8306 (
            .O(N__35135),
            .I(\uart_pc.N_143 ));
    LocalMux I__8305 (
            .O(N__35130),
            .I(\uart_pc.N_143 ));
    Odrv4 I__8304 (
            .O(N__35127),
            .I(\uart_pc.N_143 ));
    CascadeMux I__8303 (
            .O(N__35120),
            .I(N__35116));
    InMux I__8302 (
            .O(N__35119),
            .I(N__35109));
    InMux I__8301 (
            .O(N__35116),
            .I(N__35109));
    CascadeMux I__8300 (
            .O(N__35115),
            .I(N__35105));
    InMux I__8299 (
            .O(N__35114),
            .I(N__35102));
    LocalMux I__8298 (
            .O(N__35109),
            .I(N__35099));
    InMux I__8297 (
            .O(N__35108),
            .I(N__35094));
    InMux I__8296 (
            .O(N__35105),
            .I(N__35094));
    LocalMux I__8295 (
            .O(N__35102),
            .I(N__35091));
    Span4Mux_v I__8294 (
            .O(N__35099),
            .I(N__35084));
    LocalMux I__8293 (
            .O(N__35094),
            .I(N__35084));
    Span4Mux_h I__8292 (
            .O(N__35091),
            .I(N__35084));
    Odrv4 I__8291 (
            .O(N__35084),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__8290 (
            .O(N__35081),
            .I(N__35072));
    InMux I__8289 (
            .O(N__35080),
            .I(N__35069));
    IoInMux I__8288 (
            .O(N__35079),
            .I(N__35066));
    InMux I__8287 (
            .O(N__35078),
            .I(N__35060));
    InMux I__8286 (
            .O(N__35077),
            .I(N__35051));
    InMux I__8285 (
            .O(N__35076),
            .I(N__35048));
    InMux I__8284 (
            .O(N__35075),
            .I(N__35045));
    LocalMux I__8283 (
            .O(N__35072),
            .I(N__35042));
    LocalMux I__8282 (
            .O(N__35069),
            .I(N__35039));
    LocalMux I__8281 (
            .O(N__35066),
            .I(N__35036));
    CascadeMux I__8280 (
            .O(N__35065),
            .I(N__35029));
    CascadeMux I__8279 (
            .O(N__35064),
            .I(N__35026));
    InMux I__8278 (
            .O(N__35063),
            .I(N__35017));
    LocalMux I__8277 (
            .O(N__35060),
            .I(N__35014));
    InMux I__8276 (
            .O(N__35059),
            .I(N__35011));
    InMux I__8275 (
            .O(N__35058),
            .I(N__35008));
    InMux I__8274 (
            .O(N__35057),
            .I(N__34999));
    InMux I__8273 (
            .O(N__35056),
            .I(N__34999));
    InMux I__8272 (
            .O(N__35055),
            .I(N__34999));
    InMux I__8271 (
            .O(N__35054),
            .I(N__34999));
    LocalMux I__8270 (
            .O(N__35051),
            .I(N__34994));
    LocalMux I__8269 (
            .O(N__35048),
            .I(N__34994));
    LocalMux I__8268 (
            .O(N__35045),
            .I(N__34991));
    Span4Mux_v I__8267 (
            .O(N__35042),
            .I(N__34986));
    Span4Mux_h I__8266 (
            .O(N__35039),
            .I(N__34986));
    IoSpan4Mux I__8265 (
            .O(N__35036),
            .I(N__34983));
    InMux I__8264 (
            .O(N__35035),
            .I(N__34980));
    InMux I__8263 (
            .O(N__35034),
            .I(N__34975));
    InMux I__8262 (
            .O(N__35033),
            .I(N__34975));
    InMux I__8261 (
            .O(N__35032),
            .I(N__34972));
    InMux I__8260 (
            .O(N__35029),
            .I(N__34969));
    InMux I__8259 (
            .O(N__35026),
            .I(N__34966));
    InMux I__8258 (
            .O(N__35025),
            .I(N__34963));
    InMux I__8257 (
            .O(N__35024),
            .I(N__34960));
    InMux I__8256 (
            .O(N__35023),
            .I(N__34955));
    InMux I__8255 (
            .O(N__35022),
            .I(N__34955));
    InMux I__8254 (
            .O(N__35021),
            .I(N__34952));
    InMux I__8253 (
            .O(N__35020),
            .I(N__34949));
    LocalMux I__8252 (
            .O(N__35017),
            .I(N__34944));
    Span4Mux_v I__8251 (
            .O(N__35014),
            .I(N__34944));
    LocalMux I__8250 (
            .O(N__35011),
            .I(N__34941));
    LocalMux I__8249 (
            .O(N__35008),
            .I(N__34938));
    LocalMux I__8248 (
            .O(N__34999),
            .I(N__34931));
    Span4Mux_v I__8247 (
            .O(N__34994),
            .I(N__34931));
    Span4Mux_v I__8246 (
            .O(N__34991),
            .I(N__34931));
    Span4Mux_h I__8245 (
            .O(N__34986),
            .I(N__34928));
    Span4Mux_s3_v I__8244 (
            .O(N__34983),
            .I(N__34925));
    LocalMux I__8243 (
            .O(N__34980),
            .I(N__34922));
    LocalMux I__8242 (
            .O(N__34975),
            .I(N__34919));
    LocalMux I__8241 (
            .O(N__34972),
            .I(N__34916));
    LocalMux I__8240 (
            .O(N__34969),
            .I(N__34913));
    LocalMux I__8239 (
            .O(N__34966),
            .I(N__34902));
    LocalMux I__8238 (
            .O(N__34963),
            .I(N__34902));
    LocalMux I__8237 (
            .O(N__34960),
            .I(N__34902));
    LocalMux I__8236 (
            .O(N__34955),
            .I(N__34902));
    LocalMux I__8235 (
            .O(N__34952),
            .I(N__34902));
    LocalMux I__8234 (
            .O(N__34949),
            .I(N__34899));
    Sp12to4 I__8233 (
            .O(N__34944),
            .I(N__34894));
    Span12Mux_s6_v I__8232 (
            .O(N__34941),
            .I(N__34894));
    Span4Mux_v I__8231 (
            .O(N__34938),
            .I(N__34887));
    Span4Mux_h I__8230 (
            .O(N__34931),
            .I(N__34887));
    Span4Mux_h I__8229 (
            .O(N__34928),
            .I(N__34887));
    Span4Mux_v I__8228 (
            .O(N__34925),
            .I(N__34884));
    Span4Mux_v I__8227 (
            .O(N__34922),
            .I(N__34879));
    Span4Mux_v I__8226 (
            .O(N__34919),
            .I(N__34879));
    Span4Mux_h I__8225 (
            .O(N__34916),
            .I(N__34874));
    Span4Mux_h I__8224 (
            .O(N__34913),
            .I(N__34874));
    Span4Mux_v I__8223 (
            .O(N__34902),
            .I(N__34869));
    Span4Mux_h I__8222 (
            .O(N__34899),
            .I(N__34869));
    Span12Mux_v I__8221 (
            .O(N__34894),
            .I(N__34866));
    Span4Mux_v I__8220 (
            .O(N__34887),
            .I(N__34861));
    Span4Mux_h I__8219 (
            .O(N__34884),
            .I(N__34861));
    Odrv4 I__8218 (
            .O(N__34879),
            .I(reset_system));
    Odrv4 I__8217 (
            .O(N__34874),
            .I(reset_system));
    Odrv4 I__8216 (
            .O(N__34869),
            .I(reset_system));
    Odrv12 I__8215 (
            .O(N__34866),
            .I(reset_system));
    Odrv4 I__8214 (
            .O(N__34861),
            .I(reset_system));
    CascadeMux I__8213 (
            .O(N__34850),
            .I(N__34844));
    InMux I__8212 (
            .O(N__34849),
            .I(N__34841));
    InMux I__8211 (
            .O(N__34848),
            .I(N__34838));
    InMux I__8210 (
            .O(N__34847),
            .I(N__34833));
    InMux I__8209 (
            .O(N__34844),
            .I(N__34833));
    LocalMux I__8208 (
            .O(N__34841),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__8207 (
            .O(N__34838),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__8206 (
            .O(N__34833),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__8205 (
            .O(N__34826),
            .I(N__34822));
    InMux I__8204 (
            .O(N__34825),
            .I(N__34819));
    LocalMux I__8203 (
            .O(N__34822),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__8202 (
            .O(N__34819),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__8201 (
            .O(N__34814),
            .I(N__34810));
    InMux I__8200 (
            .O(N__34813),
            .I(N__34807));
    LocalMux I__8199 (
            .O(N__34810),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__8198 (
            .O(N__34807),
            .I(\reset_module_System.countZ0Z_7 ));
    CascadeMux I__8197 (
            .O(N__34802),
            .I(N__34799));
    InMux I__8196 (
            .O(N__34799),
            .I(N__34795));
    InMux I__8195 (
            .O(N__34798),
            .I(N__34792));
    LocalMux I__8194 (
            .O(N__34795),
            .I(N__34789));
    LocalMux I__8193 (
            .O(N__34792),
            .I(\reset_module_System.countZ0Z_5 ));
    Odrv4 I__8192 (
            .O(N__34789),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__8191 (
            .O(N__34784),
            .I(N__34780));
    InMux I__8190 (
            .O(N__34783),
            .I(N__34777));
    LocalMux I__8189 (
            .O(N__34780),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__8188 (
            .O(N__34777),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__8187 (
            .O(N__34772),
            .I(N__34768));
    InMux I__8186 (
            .O(N__34771),
            .I(N__34765));
    LocalMux I__8185 (
            .O(N__34768),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__8184 (
            .O(N__34765),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__8183 (
            .O(N__34760),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__8182 (
            .O(N__34757),
            .I(N__34753));
    CascadeMux I__8181 (
            .O(N__34756),
            .I(N__34748));
    LocalMux I__8180 (
            .O(N__34753),
            .I(N__34743));
    InMux I__8179 (
            .O(N__34752),
            .I(N__34738));
    InMux I__8178 (
            .O(N__34751),
            .I(N__34738));
    InMux I__8177 (
            .O(N__34748),
            .I(N__34733));
    InMux I__8176 (
            .O(N__34747),
            .I(N__34733));
    InMux I__8175 (
            .O(N__34746),
            .I(N__34730));
    Odrv4 I__8174 (
            .O(N__34743),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__8173 (
            .O(N__34738),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__8172 (
            .O(N__34733),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__8171 (
            .O(N__34730),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__8170 (
            .O(N__34721),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__8169 (
            .O(N__34718),
            .I(N__34715));
    InMux I__8168 (
            .O(N__34715),
            .I(N__34712));
    LocalMux I__8167 (
            .O(N__34712),
            .I(N__34709));
    Span4Mux_v I__8166 (
            .O(N__34709),
            .I(N__34705));
    InMux I__8165 (
            .O(N__34708),
            .I(N__34702));
    Odrv4 I__8164 (
            .O(N__34705),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__8163 (
            .O(N__34702),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__8162 (
            .O(N__34697),
            .I(N__34694));
    InMux I__8161 (
            .O(N__34694),
            .I(N__34691));
    LocalMux I__8160 (
            .O(N__34691),
            .I(N__34688));
    Span4Mux_h I__8159 (
            .O(N__34688),
            .I(N__34685));
    Odrv4 I__8158 (
            .O(N__34685),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__8157 (
            .O(N__34682),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__8156 (
            .O(N__34679),
            .I(N__34676));
    LocalMux I__8155 (
            .O(N__34676),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    InMux I__8154 (
            .O(N__34673),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__8153 (
            .O(N__34670),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__8152 (
            .O(N__34667),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__8151 (
            .O(N__34664),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__8150 (
            .O(N__34661),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__8149 (
            .O(N__34658),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__8148 (
            .O(N__34655),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__8147 (
            .O(N__34652),
            .I(bfn_12_15_0_));
    InMux I__8146 (
            .O(N__34649),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__8145 (
            .O(N__34646),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__8144 (
            .O(N__34643),
            .I(N__34640));
    InMux I__8143 (
            .O(N__34640),
            .I(N__34636));
    InMux I__8142 (
            .O(N__34639),
            .I(N__34633));
    LocalMux I__8141 (
            .O(N__34636),
            .I(N__34630));
    LocalMux I__8140 (
            .O(N__34633),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__8139 (
            .O(N__34630),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__8138 (
            .O(N__34625),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__8137 (
            .O(N__34622),
            .I(N__34618));
    InMux I__8136 (
            .O(N__34621),
            .I(N__34615));
    LocalMux I__8135 (
            .O(N__34618),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__8134 (
            .O(N__34615),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__8133 (
            .O(N__34610),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__8132 (
            .O(N__34607),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__8131 (
            .O(N__34604),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__8130 (
            .O(N__34601),
            .I(N__34597));
    InMux I__8129 (
            .O(N__34600),
            .I(N__34594));
    LocalMux I__8128 (
            .O(N__34597),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__8127 (
            .O(N__34594),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__8126 (
            .O(N__34589),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__8125 (
            .O(N__34586),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__8124 (
            .O(N__34583),
            .I(\reset_module_System.count_1_cry_7 ));
    InMux I__8123 (
            .O(N__34580),
            .I(bfn_12_14_0_));
    InMux I__8122 (
            .O(N__34577),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__8121 (
            .O(N__34574),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__8120 (
            .O(N__34571),
            .I(N__34567));
    CascadeMux I__8119 (
            .O(N__34570),
            .I(N__34562));
    LocalMux I__8118 (
            .O(N__34567),
            .I(N__34555));
    InMux I__8117 (
            .O(N__34566),
            .I(N__34552));
    InMux I__8116 (
            .O(N__34565),
            .I(N__34549));
    InMux I__8115 (
            .O(N__34562),
            .I(N__34543));
    InMux I__8114 (
            .O(N__34561),
            .I(N__34540));
    InMux I__8113 (
            .O(N__34560),
            .I(N__34533));
    InMux I__8112 (
            .O(N__34559),
            .I(N__34533));
    InMux I__8111 (
            .O(N__34558),
            .I(N__34533));
    Span4Mux_h I__8110 (
            .O(N__34555),
            .I(N__34530));
    LocalMux I__8109 (
            .O(N__34552),
            .I(N__34525));
    LocalMux I__8108 (
            .O(N__34549),
            .I(N__34525));
    InMux I__8107 (
            .O(N__34548),
            .I(N__34518));
    InMux I__8106 (
            .O(N__34547),
            .I(N__34518));
    InMux I__8105 (
            .O(N__34546),
            .I(N__34518));
    LocalMux I__8104 (
            .O(N__34543),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__8103 (
            .O(N__34540),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__8102 (
            .O(N__34533),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv4 I__8101 (
            .O(N__34530),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv12 I__8100 (
            .O(N__34525),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__8099 (
            .O(N__34518),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CascadeMux I__8098 (
            .O(N__34505),
            .I(N__34501));
    InMux I__8097 (
            .O(N__34504),
            .I(N__34494));
    InMux I__8096 (
            .O(N__34501),
            .I(N__34494));
    InMux I__8095 (
            .O(N__34500),
            .I(N__34491));
    InMux I__8094 (
            .O(N__34499),
            .I(N__34488));
    LocalMux I__8093 (
            .O(N__34494),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__8092 (
            .O(N__34491),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__8091 (
            .O(N__34488),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__8090 (
            .O(N__34481),
            .I(N__34475));
    InMux I__8089 (
            .O(N__34480),
            .I(N__34475));
    LocalMux I__8088 (
            .O(N__34475),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__8087 (
            .O(N__34472),
            .I(N__34468));
    CascadeMux I__8086 (
            .O(N__34471),
            .I(N__34463));
    LocalMux I__8085 (
            .O(N__34468),
            .I(N__34459));
    InMux I__8084 (
            .O(N__34467),
            .I(N__34456));
    InMux I__8083 (
            .O(N__34466),
            .I(N__34453));
    InMux I__8082 (
            .O(N__34463),
            .I(N__34443));
    InMux I__8081 (
            .O(N__34462),
            .I(N__34443));
    Span4Mux_h I__8080 (
            .O(N__34459),
            .I(N__34440));
    LocalMux I__8079 (
            .O(N__34456),
            .I(N__34435));
    LocalMux I__8078 (
            .O(N__34453),
            .I(N__34435));
    InMux I__8077 (
            .O(N__34452),
            .I(N__34430));
    InMux I__8076 (
            .O(N__34451),
            .I(N__34430));
    InMux I__8075 (
            .O(N__34450),
            .I(N__34427));
    InMux I__8074 (
            .O(N__34449),
            .I(N__34422));
    InMux I__8073 (
            .O(N__34448),
            .I(N__34422));
    LocalMux I__8072 (
            .O(N__34443),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv4 I__8071 (
            .O(N__34440),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv12 I__8070 (
            .O(N__34435),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__8069 (
            .O(N__34430),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__8068 (
            .O(N__34427),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__8067 (
            .O(N__34422),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__8066 (
            .O(N__34409),
            .I(N__34406));
    LocalMux I__8065 (
            .O(N__34406),
            .I(N__34402));
    CascadeMux I__8064 (
            .O(N__34405),
            .I(N__34399));
    Span4Mux_h I__8063 (
            .O(N__34402),
            .I(N__34396));
    InMux I__8062 (
            .O(N__34399),
            .I(N__34393));
    Odrv4 I__8061 (
            .O(N__34396),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__8060 (
            .O(N__34393),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    IoInMux I__8059 (
            .O(N__34388),
            .I(N__34385));
    LocalMux I__8058 (
            .O(N__34385),
            .I(N__34382));
    IoSpan4Mux I__8057 (
            .O(N__34382),
            .I(N__34374));
    CascadeMux I__8056 (
            .O(N__34381),
            .I(N__34371));
    CascadeMux I__8055 (
            .O(N__34380),
            .I(N__34368));
    CascadeMux I__8054 (
            .O(N__34379),
            .I(N__34365));
    InMux I__8053 (
            .O(N__34378),
            .I(N__34359));
    InMux I__8052 (
            .O(N__34377),
            .I(N__34356));
    Span4Mux_s0_v I__8051 (
            .O(N__34374),
            .I(N__34353));
    InMux I__8050 (
            .O(N__34371),
            .I(N__34339));
    InMux I__8049 (
            .O(N__34368),
            .I(N__34339));
    InMux I__8048 (
            .O(N__34365),
            .I(N__34339));
    InMux I__8047 (
            .O(N__34364),
            .I(N__34339));
    InMux I__8046 (
            .O(N__34363),
            .I(N__34339));
    InMux I__8045 (
            .O(N__34362),
            .I(N__34339));
    LocalMux I__8044 (
            .O(N__34359),
            .I(N__34336));
    LocalMux I__8043 (
            .O(N__34356),
            .I(N__34332));
    Sp12to4 I__8042 (
            .O(N__34353),
            .I(N__34328));
    CascadeMux I__8041 (
            .O(N__34352),
            .I(N__34325));
    LocalMux I__8040 (
            .O(N__34339),
            .I(N__34318));
    Span4Mux_h I__8039 (
            .O(N__34336),
            .I(N__34318));
    InMux I__8038 (
            .O(N__34335),
            .I(N__34315));
    Span4Mux_h I__8037 (
            .O(N__34332),
            .I(N__34312));
    InMux I__8036 (
            .O(N__34331),
            .I(N__34309));
    Span12Mux_v I__8035 (
            .O(N__34328),
            .I(N__34306));
    InMux I__8034 (
            .O(N__34325),
            .I(N__34303));
    InMux I__8033 (
            .O(N__34324),
            .I(N__34300));
    InMux I__8032 (
            .O(N__34323),
            .I(N__34297));
    Span4Mux_v I__8031 (
            .O(N__34318),
            .I(N__34294));
    LocalMux I__8030 (
            .O(N__34315),
            .I(N__34287));
    Sp12to4 I__8029 (
            .O(N__34312),
            .I(N__34287));
    LocalMux I__8028 (
            .O(N__34309),
            .I(N__34287));
    Odrv12 I__8027 (
            .O(N__34306),
            .I(debug_CH0_16A_c));
    LocalMux I__8026 (
            .O(N__34303),
            .I(debug_CH0_16A_c));
    LocalMux I__8025 (
            .O(N__34300),
            .I(debug_CH0_16A_c));
    LocalMux I__8024 (
            .O(N__34297),
            .I(debug_CH0_16A_c));
    Odrv4 I__8023 (
            .O(N__34294),
            .I(debug_CH0_16A_c));
    Odrv12 I__8022 (
            .O(N__34287),
            .I(debug_CH0_16A_c));
    InMux I__8021 (
            .O(N__34274),
            .I(N__34271));
    LocalMux I__8020 (
            .O(N__34271),
            .I(N__34261));
    InMux I__8019 (
            .O(N__34270),
            .I(N__34258));
    InMux I__8018 (
            .O(N__34269),
            .I(N__34245));
    InMux I__8017 (
            .O(N__34268),
            .I(N__34245));
    InMux I__8016 (
            .O(N__34267),
            .I(N__34245));
    InMux I__8015 (
            .O(N__34266),
            .I(N__34245));
    InMux I__8014 (
            .O(N__34265),
            .I(N__34245));
    InMux I__8013 (
            .O(N__34264),
            .I(N__34245));
    Span4Mux_v I__8012 (
            .O(N__34261),
            .I(N__34240));
    LocalMux I__8011 (
            .O(N__34258),
            .I(N__34240));
    LocalMux I__8010 (
            .O(N__34245),
            .I(N__34237));
    Span4Mux_v I__8009 (
            .O(N__34240),
            .I(N__34234));
    Span4Mux_v I__8008 (
            .O(N__34237),
            .I(N__34231));
    Odrv4 I__8007 (
            .O(N__34234),
            .I(\uart_drone.un1_state_2_0 ));
    Odrv4 I__8006 (
            .O(N__34231),
            .I(\uart_drone.un1_state_2_0 ));
    InMux I__8005 (
            .O(N__34226),
            .I(N__34223));
    LocalMux I__8004 (
            .O(N__34223),
            .I(N__34220));
    Span4Mux_h I__8003 (
            .O(N__34220),
            .I(N__34216));
    CascadeMux I__8002 (
            .O(N__34219),
            .I(N__34213));
    Span4Mux_v I__8001 (
            .O(N__34216),
            .I(N__34210));
    InMux I__8000 (
            .O(N__34213),
            .I(N__34207));
    Odrv4 I__7999 (
            .O(N__34210),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__7998 (
            .O(N__34207),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    SRMux I__7997 (
            .O(N__34202),
            .I(N__34198));
    SRMux I__7996 (
            .O(N__34201),
            .I(N__34195));
    LocalMux I__7995 (
            .O(N__34198),
            .I(N__34192));
    LocalMux I__7994 (
            .O(N__34195),
            .I(N__34189));
    Span4Mux_v I__7993 (
            .O(N__34192),
            .I(N__34186));
    Span4Mux_h I__7992 (
            .O(N__34189),
            .I(N__34183));
    Span4Mux_h I__7991 (
            .O(N__34186),
            .I(N__34179));
    Span4Mux_v I__7990 (
            .O(N__34183),
            .I(N__34176));
    SRMux I__7989 (
            .O(N__34182),
            .I(N__34173));
    Odrv4 I__7988 (
            .O(N__34179),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    Odrv4 I__7987 (
            .O(N__34176),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    LocalMux I__7986 (
            .O(N__34173),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__7985 (
            .O(N__34166),
            .I(N__34155));
    InMux I__7984 (
            .O(N__34165),
            .I(N__34144));
    InMux I__7983 (
            .O(N__34164),
            .I(N__34144));
    InMux I__7982 (
            .O(N__34163),
            .I(N__34144));
    InMux I__7981 (
            .O(N__34162),
            .I(N__34144));
    InMux I__7980 (
            .O(N__34161),
            .I(N__34144));
    InMux I__7979 (
            .O(N__34160),
            .I(N__34137));
    InMux I__7978 (
            .O(N__34159),
            .I(N__34137));
    InMux I__7977 (
            .O(N__34158),
            .I(N__34137));
    LocalMux I__7976 (
            .O(N__34155),
            .I(N__34134));
    LocalMux I__7975 (
            .O(N__34144),
            .I(N__34124));
    LocalMux I__7974 (
            .O(N__34137),
            .I(N__34124));
    Span4Mux_h I__7973 (
            .O(N__34134),
            .I(N__34121));
    InMux I__7972 (
            .O(N__34133),
            .I(N__34114));
    InMux I__7971 (
            .O(N__34132),
            .I(N__34114));
    InMux I__7970 (
            .O(N__34131),
            .I(N__34114));
    CascadeMux I__7969 (
            .O(N__34130),
            .I(N__34111));
    InMux I__7968 (
            .O(N__34129),
            .I(N__34108));
    Span4Mux_v I__7967 (
            .O(N__34124),
            .I(N__34105));
    Span4Mux_v I__7966 (
            .O(N__34121),
            .I(N__34102));
    LocalMux I__7965 (
            .O(N__34114),
            .I(N__34099));
    InMux I__7964 (
            .O(N__34111),
            .I(N__34096));
    LocalMux I__7963 (
            .O(N__34108),
            .I(N__34091));
    Span4Mux_v I__7962 (
            .O(N__34105),
            .I(N__34091));
    Span4Mux_h I__7961 (
            .O(N__34102),
            .I(N__34088));
    Sp12to4 I__7960 (
            .O(N__34099),
            .I(N__34083));
    LocalMux I__7959 (
            .O(N__34096),
            .I(N__34083));
    Odrv4 I__7958 (
            .O(N__34091),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__7957 (
            .O(N__34088),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv12 I__7956 (
            .O(N__34083),
            .I(\pid_alt.stateZ0Z_0 ));
    IoInMux I__7955 (
            .O(N__34076),
            .I(N__34073));
    LocalMux I__7954 (
            .O(N__34073),
            .I(N__34070));
    Odrv4 I__7953 (
            .O(N__34070),
            .I(\pid_alt.state_0_0 ));
    CascadeMux I__7952 (
            .O(N__34067),
            .I(\reset_module_System.reset6_15_cascade_ ));
    InMux I__7951 (
            .O(N__34064),
            .I(N__34060));
    InMux I__7950 (
            .O(N__34063),
            .I(N__34057));
    LocalMux I__7949 (
            .O(N__34060),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__7948 (
            .O(N__34057),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__7947 (
            .O(N__34052),
            .I(N__34049));
    LocalMux I__7946 (
            .O(N__34049),
            .I(\reset_module_System.count_1_2 ));
    InMux I__7945 (
            .O(N__34046),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__7944 (
            .O(N__34043),
            .I(N__34037));
    InMux I__7943 (
            .O(N__34042),
            .I(N__34032));
    InMux I__7942 (
            .O(N__34041),
            .I(N__34032));
    InMux I__7941 (
            .O(N__34040),
            .I(N__34029));
    LocalMux I__7940 (
            .O(N__34037),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__7939 (
            .O(N__34032),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__7938 (
            .O(N__34029),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__7937 (
            .O(N__34022),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__7936 (
            .O(N__34019),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    CascadeMux I__7935 (
            .O(N__34016),
            .I(N__34012));
    InMux I__7934 (
            .O(N__34015),
            .I(N__34007));
    InMux I__7933 (
            .O(N__34012),
            .I(N__34000));
    InMux I__7932 (
            .O(N__34011),
            .I(N__34000));
    InMux I__7931 (
            .O(N__34010),
            .I(N__34000));
    LocalMux I__7930 (
            .O(N__34007),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__7929 (
            .O(N__34000),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    SRMux I__7928 (
            .O(N__33995),
            .I(N__33992));
    LocalMux I__7927 (
            .O(N__33992),
            .I(N__33988));
    SRMux I__7926 (
            .O(N__33991),
            .I(N__33985));
    Span4Mux_v I__7925 (
            .O(N__33988),
            .I(N__33980));
    LocalMux I__7924 (
            .O(N__33985),
            .I(N__33980));
    Span4Mux_v I__7923 (
            .O(N__33980),
            .I(N__33977));
    Span4Mux_h I__7922 (
            .O(N__33977),
            .I(N__33974));
    Odrv4 I__7921 (
            .O(N__33974),
            .I(\Commands_frame_decoder.un1_state51_iZ0 ));
    InMux I__7920 (
            .O(N__33971),
            .I(N__33967));
    InMux I__7919 (
            .O(N__33970),
            .I(N__33964));
    LocalMux I__7918 (
            .O(N__33967),
            .I(N__33961));
    LocalMux I__7917 (
            .O(N__33964),
            .I(\uart_pc.N_144_1 ));
    Odrv4 I__7916 (
            .O(N__33961),
            .I(\uart_pc.N_144_1 ));
    InMux I__7915 (
            .O(N__33956),
            .I(N__33950));
    InMux I__7914 (
            .O(N__33955),
            .I(N__33947));
    InMux I__7913 (
            .O(N__33954),
            .I(N__33944));
    InMux I__7912 (
            .O(N__33953),
            .I(N__33941));
    LocalMux I__7911 (
            .O(N__33950),
            .I(N__33938));
    LocalMux I__7910 (
            .O(N__33947),
            .I(N__33935));
    LocalMux I__7909 (
            .O(N__33944),
            .I(N__33932));
    LocalMux I__7908 (
            .O(N__33941),
            .I(N__33929));
    Span4Mux_h I__7907 (
            .O(N__33938),
            .I(N__33926));
    Span4Mux_h I__7906 (
            .O(N__33935),
            .I(N__33923));
    Span4Mux_h I__7905 (
            .O(N__33932),
            .I(N__33918));
    Span4Mux_h I__7904 (
            .O(N__33929),
            .I(N__33918));
    Odrv4 I__7903 (
            .O(N__33926),
            .I(\uart_pc.data_rdyc_1 ));
    Odrv4 I__7902 (
            .O(N__33923),
            .I(\uart_pc.data_rdyc_1 ));
    Odrv4 I__7901 (
            .O(N__33918),
            .I(\uart_pc.data_rdyc_1 ));
    InMux I__7900 (
            .O(N__33911),
            .I(N__33908));
    LocalMux I__7899 (
            .O(N__33908),
            .I(N__33898));
    InMux I__7898 (
            .O(N__33907),
            .I(N__33893));
    InMux I__7897 (
            .O(N__33906),
            .I(N__33893));
    InMux I__7896 (
            .O(N__33905),
            .I(N__33888));
    InMux I__7895 (
            .O(N__33904),
            .I(N__33888));
    InMux I__7894 (
            .O(N__33903),
            .I(N__33885));
    InMux I__7893 (
            .O(N__33902),
            .I(N__33882));
    InMux I__7892 (
            .O(N__33901),
            .I(N__33879));
    Span4Mux_v I__7891 (
            .O(N__33898),
            .I(N__33874));
    LocalMux I__7890 (
            .O(N__33893),
            .I(N__33874));
    LocalMux I__7889 (
            .O(N__33888),
            .I(N__33871));
    LocalMux I__7888 (
            .O(N__33885),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__7887 (
            .O(N__33882),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__7886 (
            .O(N__33879),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__7885 (
            .O(N__33874),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__7884 (
            .O(N__33871),
            .I(\uart_pc.stateZ0Z_3 ));
    InMux I__7883 (
            .O(N__33860),
            .I(N__33854));
    InMux I__7882 (
            .O(N__33859),
            .I(N__33851));
    InMux I__7881 (
            .O(N__33858),
            .I(N__33848));
    InMux I__7880 (
            .O(N__33857),
            .I(N__33845));
    LocalMux I__7879 (
            .O(N__33854),
            .I(\uart_pc.N_152 ));
    LocalMux I__7878 (
            .O(N__33851),
            .I(\uart_pc.N_152 ));
    LocalMux I__7877 (
            .O(N__33848),
            .I(\uart_pc.N_152 ));
    LocalMux I__7876 (
            .O(N__33845),
            .I(\uart_pc.N_152 ));
    InMux I__7875 (
            .O(N__33836),
            .I(N__33833));
    LocalMux I__7874 (
            .O(N__33833),
            .I(\uart_pc.CO0 ));
    InMux I__7873 (
            .O(N__33830),
            .I(N__33827));
    LocalMux I__7872 (
            .O(N__33827),
            .I(N__33821));
    InMux I__7871 (
            .O(N__33826),
            .I(N__33818));
    InMux I__7870 (
            .O(N__33825),
            .I(N__33815));
    InMux I__7869 (
            .O(N__33824),
            .I(N__33807));
    Span4Mux_h I__7868 (
            .O(N__33821),
            .I(N__33804));
    LocalMux I__7867 (
            .O(N__33818),
            .I(N__33799));
    LocalMux I__7866 (
            .O(N__33815),
            .I(N__33799));
    InMux I__7865 (
            .O(N__33814),
            .I(N__33792));
    InMux I__7864 (
            .O(N__33813),
            .I(N__33792));
    InMux I__7863 (
            .O(N__33812),
            .I(N__33792));
    InMux I__7862 (
            .O(N__33811),
            .I(N__33787));
    InMux I__7861 (
            .O(N__33810),
            .I(N__33787));
    LocalMux I__7860 (
            .O(N__33807),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    Odrv4 I__7859 (
            .O(N__33804),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    Odrv12 I__7858 (
            .O(N__33799),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__7857 (
            .O(N__33792),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__7856 (
            .O(N__33787),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__7855 (
            .O(N__33776),
            .I(N__33772));
    InMux I__7854 (
            .O(N__33775),
            .I(N__33769));
    LocalMux I__7853 (
            .O(N__33772),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__7852 (
            .O(N__33769),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__7851 (
            .O(N__33764),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__7850 (
            .O(N__33761),
            .I(N__33757));
    InMux I__7849 (
            .O(N__33760),
            .I(N__33754));
    LocalMux I__7848 (
            .O(N__33757),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__7847 (
            .O(N__33754),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__7846 (
            .O(N__33749),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__7845 (
            .O(N__33746),
            .I(N__33742));
    InMux I__7844 (
            .O(N__33745),
            .I(N__33739));
    LocalMux I__7843 (
            .O(N__33742),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__7842 (
            .O(N__33739),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__7841 (
            .O(N__33734),
            .I(bfn_11_16_0_));
    CascadeMux I__7840 (
            .O(N__33731),
            .I(N__33727));
    InMux I__7839 (
            .O(N__33730),
            .I(N__33724));
    InMux I__7838 (
            .O(N__33727),
            .I(N__33721));
    LocalMux I__7837 (
            .O(N__33724),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__7836 (
            .O(N__33721),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__7835 (
            .O(N__33716),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__7834 (
            .O(N__33713),
            .I(N__33709));
    InMux I__7833 (
            .O(N__33712),
            .I(N__33706));
    LocalMux I__7832 (
            .O(N__33709),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__7831 (
            .O(N__33706),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__7830 (
            .O(N__33701),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__7829 (
            .O(N__33698),
            .I(N__33693));
    InMux I__7828 (
            .O(N__33697),
            .I(N__33688));
    InMux I__7827 (
            .O(N__33696),
            .I(N__33688));
    LocalMux I__7826 (
            .O(N__33693),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__7825 (
            .O(N__33688),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__7824 (
            .O(N__33683),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__7823 (
            .O(N__33680),
            .I(N__33675));
    InMux I__7822 (
            .O(N__33679),
            .I(N__33670));
    InMux I__7821 (
            .O(N__33678),
            .I(N__33670));
    LocalMux I__7820 (
            .O(N__33675),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__7819 (
            .O(N__33670),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__7818 (
            .O(N__33665),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    CascadeMux I__7817 (
            .O(N__33662),
            .I(N__33658));
    InMux I__7816 (
            .O(N__33661),
            .I(N__33655));
    InMux I__7815 (
            .O(N__33658),
            .I(N__33652));
    LocalMux I__7814 (
            .O(N__33655),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__7813 (
            .O(N__33652),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__7812 (
            .O(N__33647),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__7811 (
            .O(N__33644),
            .I(N__33637));
    InMux I__7810 (
            .O(N__33643),
            .I(N__33634));
    CascadeMux I__7809 (
            .O(N__33642),
            .I(N__33625));
    CascadeMux I__7808 (
            .O(N__33641),
            .I(N__33618));
    CascadeMux I__7807 (
            .O(N__33640),
            .I(N__33614));
    LocalMux I__7806 (
            .O(N__33637),
            .I(N__33609));
    LocalMux I__7805 (
            .O(N__33634),
            .I(N__33606));
    InMux I__7804 (
            .O(N__33633),
            .I(N__33603));
    InMux I__7803 (
            .O(N__33632),
            .I(N__33600));
    InMux I__7802 (
            .O(N__33631),
            .I(N__33597));
    InMux I__7801 (
            .O(N__33630),
            .I(N__33592));
    InMux I__7800 (
            .O(N__33629),
            .I(N__33592));
    InMux I__7799 (
            .O(N__33628),
            .I(N__33589));
    InMux I__7798 (
            .O(N__33625),
            .I(N__33580));
    InMux I__7797 (
            .O(N__33624),
            .I(N__33580));
    InMux I__7796 (
            .O(N__33623),
            .I(N__33580));
    InMux I__7795 (
            .O(N__33622),
            .I(N__33580));
    InMux I__7794 (
            .O(N__33621),
            .I(N__33577));
    InMux I__7793 (
            .O(N__33618),
            .I(N__33570));
    InMux I__7792 (
            .O(N__33617),
            .I(N__33570));
    InMux I__7791 (
            .O(N__33614),
            .I(N__33570));
    InMux I__7790 (
            .O(N__33613),
            .I(N__33567));
    InMux I__7789 (
            .O(N__33612),
            .I(N__33564));
    Span4Mux_h I__7788 (
            .O(N__33609),
            .I(N__33549));
    Span4Mux_v I__7787 (
            .O(N__33606),
            .I(N__33549));
    LocalMux I__7786 (
            .O(N__33603),
            .I(N__33549));
    LocalMux I__7785 (
            .O(N__33600),
            .I(N__33549));
    LocalMux I__7784 (
            .O(N__33597),
            .I(N__33549));
    LocalMux I__7783 (
            .O(N__33592),
            .I(N__33546));
    LocalMux I__7782 (
            .O(N__33589),
            .I(N__33543));
    LocalMux I__7781 (
            .O(N__33580),
            .I(N__33538));
    LocalMux I__7780 (
            .O(N__33577),
            .I(N__33538));
    LocalMux I__7779 (
            .O(N__33570),
            .I(N__33535));
    LocalMux I__7778 (
            .O(N__33567),
            .I(N__33530));
    LocalMux I__7777 (
            .O(N__33564),
            .I(N__33530));
    InMux I__7776 (
            .O(N__33563),
            .I(N__33527));
    InMux I__7775 (
            .O(N__33562),
            .I(N__33524));
    InMux I__7774 (
            .O(N__33561),
            .I(N__33519));
    InMux I__7773 (
            .O(N__33560),
            .I(N__33519));
    Span4Mux_v I__7772 (
            .O(N__33549),
            .I(N__33514));
    Span4Mux_h I__7771 (
            .O(N__33546),
            .I(N__33514));
    Span4Mux_h I__7770 (
            .O(N__33543),
            .I(N__33507));
    Span4Mux_h I__7769 (
            .O(N__33538),
            .I(N__33507));
    Span4Mux_h I__7768 (
            .O(N__33535),
            .I(N__33507));
    Odrv4 I__7767 (
            .O(N__33530),
            .I(uart_pc_data_rdy));
    LocalMux I__7766 (
            .O(N__33527),
            .I(uart_pc_data_rdy));
    LocalMux I__7765 (
            .O(N__33524),
            .I(uart_pc_data_rdy));
    LocalMux I__7764 (
            .O(N__33519),
            .I(uart_pc_data_rdy));
    Odrv4 I__7763 (
            .O(N__33514),
            .I(uart_pc_data_rdy));
    Odrv4 I__7762 (
            .O(N__33507),
            .I(uart_pc_data_rdy));
    InMux I__7761 (
            .O(N__33494),
            .I(N__33485));
    InMux I__7760 (
            .O(N__33493),
            .I(N__33485));
    InMux I__7759 (
            .O(N__33492),
            .I(N__33482));
    InMux I__7758 (
            .O(N__33491),
            .I(N__33477));
    InMux I__7757 (
            .O(N__33490),
            .I(N__33477));
    LocalMux I__7756 (
            .O(N__33485),
            .I(N__33474));
    LocalMux I__7755 (
            .O(N__33482),
            .I(N__33471));
    LocalMux I__7754 (
            .O(N__33477),
            .I(N__33468));
    Span4Mux_h I__7753 (
            .O(N__33474),
            .I(N__33462));
    Span4Mux_v I__7752 (
            .O(N__33471),
            .I(N__33462));
    Span4Mux_h I__7751 (
            .O(N__33468),
            .I(N__33459));
    InMux I__7750 (
            .O(N__33467),
            .I(N__33456));
    Odrv4 I__7749 (
            .O(N__33462),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    Odrv4 I__7748 (
            .O(N__33459),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    LocalMux I__7747 (
            .O(N__33456),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    InMux I__7746 (
            .O(N__33449),
            .I(N__33440));
    InMux I__7745 (
            .O(N__33448),
            .I(N__33440));
    InMux I__7744 (
            .O(N__33447),
            .I(N__33440));
    LocalMux I__7743 (
            .O(N__33440),
            .I(\Commands_frame_decoder.count_RNIDLVE1Z0Z_2 ));
    CascadeMux I__7742 (
            .O(N__33437),
            .I(N__33434));
    InMux I__7741 (
            .O(N__33434),
            .I(N__33428));
    InMux I__7740 (
            .O(N__33433),
            .I(N__33428));
    LocalMux I__7739 (
            .O(N__33428),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    CascadeMux I__7738 (
            .O(N__33425),
            .I(N__33421));
    InMux I__7737 (
            .O(N__33424),
            .I(N__33414));
    InMux I__7736 (
            .O(N__33421),
            .I(N__33414));
    CascadeMux I__7735 (
            .O(N__33420),
            .I(N__33411));
    CascadeMux I__7734 (
            .O(N__33419),
            .I(N__33408));
    LocalMux I__7733 (
            .O(N__33414),
            .I(N__33405));
    InMux I__7732 (
            .O(N__33411),
            .I(N__33402));
    InMux I__7731 (
            .O(N__33408),
            .I(N__33399));
    Odrv4 I__7730 (
            .O(N__33405),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__7729 (
            .O(N__33402),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__7728 (
            .O(N__33399),
            .I(\uart_pc.stateZ0Z_2 ));
    CascadeMux I__7727 (
            .O(N__33392),
            .I(N__33388));
    InMux I__7726 (
            .O(N__33391),
            .I(N__33385));
    InMux I__7725 (
            .O(N__33388),
            .I(N__33382));
    LocalMux I__7724 (
            .O(N__33385),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__7723 (
            .O(N__33382),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__7722 (
            .O(N__33377),
            .I(N__33374));
    LocalMux I__7721 (
            .O(N__33374),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__7720 (
            .O(N__33371),
            .I(N__33368));
    LocalMux I__7719 (
            .O(N__33368),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__7718 (
            .O(N__33365),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__7717 (
            .O(N__33362),
            .I(N__33359));
    LocalMux I__7716 (
            .O(N__33359),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__7715 (
            .O(N__33356),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__7714 (
            .O(N__33353),
            .I(N__33350));
    LocalMux I__7713 (
            .O(N__33350),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__7712 (
            .O(N__33347),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__7711 (
            .O(N__33344),
            .I(N__33340));
    InMux I__7710 (
            .O(N__33343),
            .I(N__33337));
    LocalMux I__7709 (
            .O(N__33340),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__7708 (
            .O(N__33337),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__7707 (
            .O(N__33332),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__7706 (
            .O(N__33329),
            .I(N__33325));
    InMux I__7705 (
            .O(N__33328),
            .I(N__33322));
    LocalMux I__7704 (
            .O(N__33325),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__7703 (
            .O(N__33322),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    InMux I__7702 (
            .O(N__33317),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__7701 (
            .O(N__33314),
            .I(N__33309));
    InMux I__7700 (
            .O(N__33313),
            .I(N__33304));
    InMux I__7699 (
            .O(N__33312),
            .I(N__33304));
    LocalMux I__7698 (
            .O(N__33309),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__7697 (
            .O(N__33304),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__7696 (
            .O(N__33299),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__7695 (
            .O(N__33296),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    InMux I__7694 (
            .O(N__33293),
            .I(N__33288));
    InMux I__7693 (
            .O(N__33292),
            .I(N__33283));
    InMux I__7692 (
            .O(N__33291),
            .I(N__33283));
    LocalMux I__7691 (
            .O(N__33288),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__7690 (
            .O(N__33283),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    SRMux I__7689 (
            .O(N__33278),
            .I(N__33274));
    SRMux I__7688 (
            .O(N__33277),
            .I(N__33271));
    LocalMux I__7687 (
            .O(N__33274),
            .I(N__33268));
    LocalMux I__7686 (
            .O(N__33271),
            .I(N__33265));
    Span4Mux_v I__7685 (
            .O(N__33268),
            .I(N__33262));
    Span4Mux_h I__7684 (
            .O(N__33265),
            .I(N__33259));
    Span4Mux_v I__7683 (
            .O(N__33262),
            .I(N__33254));
    Span4Mux_v I__7682 (
            .O(N__33259),
            .I(N__33254));
    Odrv4 I__7681 (
            .O(N__33254),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    CascadeMux I__7680 (
            .O(N__33251),
            .I(N__33246));
    InMux I__7679 (
            .O(N__33250),
            .I(N__33243));
    InMux I__7678 (
            .O(N__33249),
            .I(N__33240));
    InMux I__7677 (
            .O(N__33246),
            .I(N__33237));
    LocalMux I__7676 (
            .O(N__33243),
            .I(N__33234));
    LocalMux I__7675 (
            .O(N__33240),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__7674 (
            .O(N__33237),
            .I(\uart_pc.stateZ0Z_1 ));
    Odrv12 I__7673 (
            .O(N__33234),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__7672 (
            .O(N__33227),
            .I(N__33221));
    InMux I__7671 (
            .O(N__33226),
            .I(N__33218));
    InMux I__7670 (
            .O(N__33225),
            .I(N__33215));
    InMux I__7669 (
            .O(N__33224),
            .I(N__33210));
    InMux I__7668 (
            .O(N__33221),
            .I(N__33210));
    LocalMux I__7667 (
            .O(N__33218),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__7666 (
            .O(N__33215),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__7665 (
            .O(N__33210),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    InMux I__7664 (
            .O(N__33203),
            .I(N__33199));
    InMux I__7663 (
            .O(N__33202),
            .I(N__33196));
    LocalMux I__7662 (
            .O(N__33199),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__7661 (
            .O(N__33196),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    InMux I__7660 (
            .O(N__33191),
            .I(N__33188));
    LocalMux I__7659 (
            .O(N__33188),
            .I(\uart_drone.timer_Count_RNO_0_0_1 ));
    CascadeMux I__7658 (
            .O(N__33185),
            .I(\Commands_frame_decoder.CO0_cascade_ ));
    InMux I__7657 (
            .O(N__33182),
            .I(N__33179));
    LocalMux I__7656 (
            .O(N__33179),
            .I(\Commands_frame_decoder.CO0 ));
    InMux I__7655 (
            .O(N__33176),
            .I(N__33170));
    InMux I__7654 (
            .O(N__33175),
            .I(N__33170));
    LocalMux I__7653 (
            .O(N__33170),
            .I(\Commands_frame_decoder.countZ0Z_1 ));
    CascadeMux I__7652 (
            .O(N__33167),
            .I(N__33163));
    InMux I__7651 (
            .O(N__33166),
            .I(N__33160));
    InMux I__7650 (
            .O(N__33163),
            .I(N__33156));
    LocalMux I__7649 (
            .O(N__33160),
            .I(N__33153));
    CascadeMux I__7648 (
            .O(N__33159),
            .I(N__33150));
    LocalMux I__7647 (
            .O(N__33156),
            .I(N__33144));
    Span4Mux_v I__7646 (
            .O(N__33153),
            .I(N__33144));
    InMux I__7645 (
            .O(N__33150),
            .I(N__33139));
    InMux I__7644 (
            .O(N__33149),
            .I(N__33139));
    Odrv4 I__7643 (
            .O(N__33144),
            .I(\Commands_frame_decoder.countZ0Z_2 ));
    LocalMux I__7642 (
            .O(N__33139),
            .I(\Commands_frame_decoder.countZ0Z_2 ));
    InMux I__7641 (
            .O(N__33134),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__7640 (
            .O(N__33131),
            .I(N__33127));
    InMux I__7639 (
            .O(N__33130),
            .I(N__33124));
    LocalMux I__7638 (
            .O(N__33127),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    LocalMux I__7637 (
            .O(N__33124),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__7636 (
            .O(N__33119),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__7635 (
            .O(N__33116),
            .I(N__33112));
    InMux I__7634 (
            .O(N__33115),
            .I(N__33109));
    LocalMux I__7633 (
            .O(N__33112),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    LocalMux I__7632 (
            .O(N__33109),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    InMux I__7631 (
            .O(N__33104),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__7630 (
            .O(N__33101),
            .I(N__33097));
    InMux I__7629 (
            .O(N__33100),
            .I(N__33094));
    LocalMux I__7628 (
            .O(N__33097),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__7627 (
            .O(N__33094),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__7626 (
            .O(N__33089),
            .I(bfn_10_20_0_));
    CascadeMux I__7625 (
            .O(N__33086),
            .I(N__33082));
    InMux I__7624 (
            .O(N__33085),
            .I(N__33079));
    InMux I__7623 (
            .O(N__33082),
            .I(N__33076));
    LocalMux I__7622 (
            .O(N__33079),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__7621 (
            .O(N__33076),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__7620 (
            .O(N__33071),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__7619 (
            .O(N__33068),
            .I(N__33064));
    InMux I__7618 (
            .O(N__33067),
            .I(N__33061));
    LocalMux I__7617 (
            .O(N__33064),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__7616 (
            .O(N__33061),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__7615 (
            .O(N__33056),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__7614 (
            .O(N__33053),
            .I(N__33048));
    InMux I__7613 (
            .O(N__33052),
            .I(N__33045));
    InMux I__7612 (
            .O(N__33051),
            .I(N__33042));
    LocalMux I__7611 (
            .O(N__33048),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__7610 (
            .O(N__33045),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__7609 (
            .O(N__33042),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__7608 (
            .O(N__33035),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__7607 (
            .O(N__33032),
            .I(N__33027));
    InMux I__7606 (
            .O(N__33031),
            .I(N__33024));
    InMux I__7605 (
            .O(N__33030),
            .I(N__33021));
    LocalMux I__7604 (
            .O(N__33027),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__7603 (
            .O(N__33024),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__7602 (
            .O(N__33021),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__7601 (
            .O(N__33014),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    CascadeMux I__7600 (
            .O(N__33011),
            .I(N__33007));
    InMux I__7599 (
            .O(N__33010),
            .I(N__33004));
    InMux I__7598 (
            .O(N__33007),
            .I(N__33001));
    LocalMux I__7597 (
            .O(N__33004),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__7596 (
            .O(N__33001),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__7595 (
            .O(N__32996),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__7594 (
            .O(N__32993),
            .I(N__32990));
    LocalMux I__7593 (
            .O(N__32990),
            .I(N__32987));
    Odrv4 I__7592 (
            .O(N__32987),
            .I(\uart_pc.data_Auxce_0_5 ));
    CascadeMux I__7591 (
            .O(N__32984),
            .I(N__32980));
    InMux I__7590 (
            .O(N__32983),
            .I(N__32977));
    InMux I__7589 (
            .O(N__32980),
            .I(N__32974));
    LocalMux I__7588 (
            .O(N__32977),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__7587 (
            .O(N__32974),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__7586 (
            .O(N__32969),
            .I(N__32966));
    LocalMux I__7585 (
            .O(N__32966),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__7584 (
            .O(N__32963),
            .I(N__32960));
    LocalMux I__7583 (
            .O(N__32960),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__7582 (
            .O(N__32957),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__7581 (
            .O(N__32954),
            .I(N__32951));
    LocalMux I__7580 (
            .O(N__32951),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__7579 (
            .O(N__32948),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__7578 (
            .O(N__32945),
            .I(N__32942));
    LocalMux I__7577 (
            .O(N__32942),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__7576 (
            .O(N__32939),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__7575 (
            .O(N__32936),
            .I(N__32932));
    InMux I__7574 (
            .O(N__32935),
            .I(N__32929));
    LocalMux I__7573 (
            .O(N__32932),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    LocalMux I__7572 (
            .O(N__32929),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__7571 (
            .O(N__32924),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__7570 (
            .O(N__32921),
            .I(N__32917));
    InMux I__7569 (
            .O(N__32920),
            .I(N__32914));
    LocalMux I__7568 (
            .O(N__32917),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    LocalMux I__7567 (
            .O(N__32914),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    InMux I__7566 (
            .O(N__32909),
            .I(N__32905));
    InMux I__7565 (
            .O(N__32908),
            .I(N__32902));
    LocalMux I__7564 (
            .O(N__32905),
            .I(N__32897));
    LocalMux I__7563 (
            .O(N__32902),
            .I(N__32897));
    Span4Mux_h I__7562 (
            .O(N__32897),
            .I(N__32894));
    Odrv4 I__7561 (
            .O(N__32894),
            .I(\Commands_frame_decoder.N_303_0 ));
    InMux I__7560 (
            .O(N__32891),
            .I(N__32885));
    InMux I__7559 (
            .O(N__32890),
            .I(N__32885));
    LocalMux I__7558 (
            .O(N__32885),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    InMux I__7557 (
            .O(N__32882),
            .I(N__32876));
    InMux I__7556 (
            .O(N__32881),
            .I(N__32876));
    LocalMux I__7555 (
            .O(N__32876),
            .I(N__32864));
    InMux I__7554 (
            .O(N__32875),
            .I(N__32857));
    InMux I__7553 (
            .O(N__32874),
            .I(N__32857));
    InMux I__7552 (
            .O(N__32873),
            .I(N__32857));
    InMux I__7551 (
            .O(N__32872),
            .I(N__32852));
    InMux I__7550 (
            .O(N__32871),
            .I(N__32852));
    InMux I__7549 (
            .O(N__32870),
            .I(N__32849));
    InMux I__7548 (
            .O(N__32869),
            .I(N__32842));
    InMux I__7547 (
            .O(N__32868),
            .I(N__32842));
    InMux I__7546 (
            .O(N__32867),
            .I(N__32842));
    Sp12to4 I__7545 (
            .O(N__32864),
            .I(N__32837));
    LocalMux I__7544 (
            .O(N__32857),
            .I(N__32837));
    LocalMux I__7543 (
            .O(N__32852),
            .I(N__32832));
    LocalMux I__7542 (
            .O(N__32849),
            .I(N__32832));
    LocalMux I__7541 (
            .O(N__32842),
            .I(N__32829));
    Span12Mux_v I__7540 (
            .O(N__32837),
            .I(N__32826));
    Span4Mux_v I__7539 (
            .O(N__32832),
            .I(N__32823));
    Span4Mux_h I__7538 (
            .O(N__32829),
            .I(N__32820));
    Odrv12 I__7537 (
            .O(N__32826),
            .I(\Commands_frame_decoder.N_335 ));
    Odrv4 I__7536 (
            .O(N__32823),
            .I(\Commands_frame_decoder.N_335 ));
    Odrv4 I__7535 (
            .O(N__32820),
            .I(\Commands_frame_decoder.N_335 ));
    CascadeMux I__7534 (
            .O(N__32813),
            .I(N__32810));
    InMux I__7533 (
            .O(N__32810),
            .I(N__32807));
    LocalMux I__7532 (
            .O(N__32807),
            .I(N__32802));
    InMux I__7531 (
            .O(N__32806),
            .I(N__32797));
    InMux I__7530 (
            .O(N__32805),
            .I(N__32797));
    Odrv12 I__7529 (
            .O(N__32802),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__7528 (
            .O(N__32797),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__7527 (
            .O(N__32792),
            .I(N__32789));
    LocalMux I__7526 (
            .O(N__32789),
            .I(\uart_pc.data_Auxce_0_6 ));
    InMux I__7525 (
            .O(N__32786),
            .I(N__32783));
    LocalMux I__7524 (
            .O(N__32783),
            .I(N__32780));
    Odrv4 I__7523 (
            .O(N__32780),
            .I(\uart_pc.data_Auxce_0_1 ));
    InMux I__7522 (
            .O(N__32777),
            .I(N__32774));
    LocalMux I__7521 (
            .O(N__32774),
            .I(N__32771));
    Odrv4 I__7520 (
            .O(N__32771),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__7519 (
            .O(N__32768),
            .I(N__32765));
    LocalMux I__7518 (
            .O(N__32765),
            .I(N__32762));
    Span4Mux_h I__7517 (
            .O(N__32762),
            .I(N__32759));
    Odrv4 I__7516 (
            .O(N__32759),
            .I(\uart_drone.data_Auxce_0_1 ));
    CascadeMux I__7515 (
            .O(N__32756),
            .I(\uart_pc.un1_state_2_0_cascade_ ));
    CascadeMux I__7514 (
            .O(N__32753),
            .I(N__32750));
    InMux I__7513 (
            .O(N__32750),
            .I(N__32746));
    InMux I__7512 (
            .O(N__32749),
            .I(N__32743));
    LocalMux I__7511 (
            .O(N__32746),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__7510 (
            .O(N__32743),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__7509 (
            .O(N__32738),
            .I(N__32735));
    LocalMux I__7508 (
            .O(N__32735),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    CascadeMux I__7507 (
            .O(N__32732),
            .I(N__32729));
    InMux I__7506 (
            .O(N__32729),
            .I(N__32725));
    CascadeMux I__7505 (
            .O(N__32728),
            .I(N__32722));
    LocalMux I__7504 (
            .O(N__32725),
            .I(N__32719));
    InMux I__7503 (
            .O(N__32722),
            .I(N__32716));
    Odrv4 I__7502 (
            .O(N__32719),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__7501 (
            .O(N__32716),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    CascadeMux I__7500 (
            .O(N__32711),
            .I(N__32707));
    InMux I__7499 (
            .O(N__32710),
            .I(N__32704));
    InMux I__7498 (
            .O(N__32707),
            .I(N__32701));
    LocalMux I__7497 (
            .O(N__32704),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__7496 (
            .O(N__32701),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__7495 (
            .O(N__32696),
            .I(N__32692));
    CascadeMux I__7494 (
            .O(N__32695),
            .I(N__32689));
    LocalMux I__7493 (
            .O(N__32692),
            .I(N__32686));
    InMux I__7492 (
            .O(N__32689),
            .I(N__32683));
    Odrv4 I__7491 (
            .O(N__32686),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__7490 (
            .O(N__32683),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__7489 (
            .O(N__32678),
            .I(\Commands_frame_decoder.WDT8lto13_1_cascade_ ));
    InMux I__7488 (
            .O(N__32675),
            .I(N__32672));
    LocalMux I__7487 (
            .O(N__32672),
            .I(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ));
    CascadeMux I__7486 (
            .O(N__32669),
            .I(\Commands_frame_decoder.WDT8lt14_0_cascade_ ));
    InMux I__7485 (
            .O(N__32666),
            .I(N__32663));
    LocalMux I__7484 (
            .O(N__32663),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    InMux I__7483 (
            .O(N__32660),
            .I(N__32657));
    LocalMux I__7482 (
            .O(N__32657),
            .I(\uart_pc.state_srsts_i_0_2 ));
    CascadeMux I__7481 (
            .O(N__32654),
            .I(\uart_pc.N_145_cascade_ ));
    InMux I__7480 (
            .O(N__32651),
            .I(N__32646));
    InMux I__7479 (
            .O(N__32650),
            .I(N__32637));
    InMux I__7478 (
            .O(N__32649),
            .I(N__32637));
    LocalMux I__7477 (
            .O(N__32646),
            .I(N__32634));
    InMux I__7476 (
            .O(N__32645),
            .I(N__32629));
    InMux I__7475 (
            .O(N__32644),
            .I(N__32629));
    InMux I__7474 (
            .O(N__32643),
            .I(N__32624));
    InMux I__7473 (
            .O(N__32642),
            .I(N__32621));
    LocalMux I__7472 (
            .O(N__32637),
            .I(N__32614));
    Span4Mux_h I__7471 (
            .O(N__32634),
            .I(N__32614));
    LocalMux I__7470 (
            .O(N__32629),
            .I(N__32614));
    InMux I__7469 (
            .O(N__32628),
            .I(N__32609));
    InMux I__7468 (
            .O(N__32627),
            .I(N__32609));
    LocalMux I__7467 (
            .O(N__32624),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7466 (
            .O(N__32621),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__7465 (
            .O(N__32614),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7464 (
            .O(N__32609),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__7463 (
            .O(N__32600),
            .I(N__32594));
    InMux I__7462 (
            .O(N__32599),
            .I(N__32591));
    InMux I__7461 (
            .O(N__32598),
            .I(N__32582));
    InMux I__7460 (
            .O(N__32597),
            .I(N__32582));
    LocalMux I__7459 (
            .O(N__32594),
            .I(N__32579));
    LocalMux I__7458 (
            .O(N__32591),
            .I(N__32576));
    InMux I__7457 (
            .O(N__32590),
            .I(N__32573));
    InMux I__7456 (
            .O(N__32589),
            .I(N__32568));
    InMux I__7455 (
            .O(N__32588),
            .I(N__32568));
    InMux I__7454 (
            .O(N__32587),
            .I(N__32565));
    LocalMux I__7453 (
            .O(N__32582),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__7452 (
            .O(N__32579),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__7451 (
            .O(N__32576),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7450 (
            .O(N__32573),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7449 (
            .O(N__32568),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7448 (
            .O(N__32565),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__7447 (
            .O(N__32552),
            .I(N__32549));
    LocalMux I__7446 (
            .O(N__32549),
            .I(N__32546));
    Odrv4 I__7445 (
            .O(N__32546),
            .I(\uart_drone.N_145 ));
    CascadeMux I__7444 (
            .O(N__32543),
            .I(N__32539));
    CascadeMux I__7443 (
            .O(N__32542),
            .I(N__32536));
    InMux I__7442 (
            .O(N__32539),
            .I(N__32531));
    InMux I__7441 (
            .O(N__32536),
            .I(N__32528));
    InMux I__7440 (
            .O(N__32535),
            .I(N__32525));
    InMux I__7439 (
            .O(N__32534),
            .I(N__32522));
    LocalMux I__7438 (
            .O(N__32531),
            .I(N__32517));
    LocalMux I__7437 (
            .O(N__32528),
            .I(N__32517));
    LocalMux I__7436 (
            .O(N__32525),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__7435 (
            .O(N__32522),
            .I(\uart_drone.stateZ0Z_2 ));
    Odrv4 I__7434 (
            .O(N__32517),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__7433 (
            .O(N__32510),
            .I(\uart_drone.N_144_1_cascade_ ));
    InMux I__7432 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__7431 (
            .O(N__32504),
            .I(\uart_drone.N_144_1 ));
    CascadeMux I__7430 (
            .O(N__32501),
            .I(N__32496));
    CascadeMux I__7429 (
            .O(N__32500),
            .I(N__32493));
    CascadeMux I__7428 (
            .O(N__32499),
            .I(N__32488));
    InMux I__7427 (
            .O(N__32496),
            .I(N__32479));
    InMux I__7426 (
            .O(N__32493),
            .I(N__32479));
    InMux I__7425 (
            .O(N__32492),
            .I(N__32479));
    InMux I__7424 (
            .O(N__32491),
            .I(N__32479));
    InMux I__7423 (
            .O(N__32488),
            .I(N__32476));
    LocalMux I__7422 (
            .O(N__32479),
            .I(\uart_drone.N_143 ));
    LocalMux I__7421 (
            .O(N__32476),
            .I(\uart_drone.N_143 ));
    InMux I__7420 (
            .O(N__32471),
            .I(N__32468));
    LocalMux I__7419 (
            .O(N__32468),
            .I(N__32461));
    CascadeMux I__7418 (
            .O(N__32467),
            .I(N__32457));
    InMux I__7417 (
            .O(N__32466),
            .I(N__32454));
    InMux I__7416 (
            .O(N__32465),
            .I(N__32449));
    InMux I__7415 (
            .O(N__32464),
            .I(N__32449));
    Span4Mux_h I__7414 (
            .O(N__32461),
            .I(N__32446));
    InMux I__7413 (
            .O(N__32460),
            .I(N__32443));
    InMux I__7412 (
            .O(N__32457),
            .I(N__32440));
    LocalMux I__7411 (
            .O(N__32454),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7410 (
            .O(N__32449),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__7409 (
            .O(N__32446),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7408 (
            .O(N__32443),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7407 (
            .O(N__32440),
            .I(\uart_drone.stateZ0Z_4 ));
    InMux I__7406 (
            .O(N__32429),
            .I(N__32426));
    LocalMux I__7405 (
            .O(N__32426),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    InMux I__7404 (
            .O(N__32423),
            .I(N__32418));
    InMux I__7403 (
            .O(N__32422),
            .I(N__32410));
    InMux I__7402 (
            .O(N__32421),
            .I(N__32407));
    LocalMux I__7401 (
            .O(N__32418),
            .I(N__32403));
    InMux I__7400 (
            .O(N__32417),
            .I(N__32400));
    InMux I__7399 (
            .O(N__32416),
            .I(N__32397));
    InMux I__7398 (
            .O(N__32415),
            .I(N__32390));
    InMux I__7397 (
            .O(N__32414),
            .I(N__32390));
    InMux I__7396 (
            .O(N__32413),
            .I(N__32390));
    LocalMux I__7395 (
            .O(N__32410),
            .I(N__32384));
    LocalMux I__7394 (
            .O(N__32407),
            .I(N__32384));
    InMux I__7393 (
            .O(N__32406),
            .I(N__32381));
    Span4Mux_v I__7392 (
            .O(N__32403),
            .I(N__32376));
    LocalMux I__7391 (
            .O(N__32400),
            .I(N__32376));
    LocalMux I__7390 (
            .O(N__32397),
            .I(N__32373));
    LocalMux I__7389 (
            .O(N__32390),
            .I(N__32370));
    InMux I__7388 (
            .O(N__32389),
            .I(N__32367));
    Span4Mux_v I__7387 (
            .O(N__32384),
            .I(N__32364));
    LocalMux I__7386 (
            .O(N__32381),
            .I(N__32357));
    Span4Mux_v I__7385 (
            .O(N__32376),
            .I(N__32357));
    Span4Mux_h I__7384 (
            .O(N__32373),
            .I(N__32357));
    Span4Mux_h I__7383 (
            .O(N__32370),
            .I(N__32353));
    LocalMux I__7382 (
            .O(N__32367),
            .I(N__32350));
    Span4Mux_h I__7381 (
            .O(N__32364),
            .I(N__32345));
    Span4Mux_v I__7380 (
            .O(N__32357),
            .I(N__32345));
    InMux I__7379 (
            .O(N__32356),
            .I(N__32342));
    Odrv4 I__7378 (
            .O(N__32353),
            .I(uart_drone_data_rdy));
    Odrv4 I__7377 (
            .O(N__32350),
            .I(uart_drone_data_rdy));
    Odrv4 I__7376 (
            .O(N__32345),
            .I(uart_drone_data_rdy));
    LocalMux I__7375 (
            .O(N__32342),
            .I(uart_drone_data_rdy));
    InMux I__7374 (
            .O(N__32333),
            .I(N__32330));
    LocalMux I__7373 (
            .O(N__32330),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__7372 (
            .O(N__32327),
            .I(N__32322));
    InMux I__7371 (
            .O(N__32326),
            .I(N__32319));
    InMux I__7370 (
            .O(N__32325),
            .I(N__32316));
    LocalMux I__7369 (
            .O(N__32322),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__7368 (
            .O(N__32319),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__7367 (
            .O(N__32316),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__7366 (
            .O(N__32309),
            .I(N__32306));
    LocalMux I__7365 (
            .O(N__32306),
            .I(N__32303));
    Odrv12 I__7364 (
            .O(N__32303),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    CascadeMux I__7363 (
            .O(N__32300),
            .I(N__32297));
    InMux I__7362 (
            .O(N__32297),
            .I(N__32294));
    LocalMux I__7361 (
            .O(N__32294),
            .I(N__32291));
    Span4Mux_h I__7360 (
            .O(N__32291),
            .I(N__32287));
    InMux I__7359 (
            .O(N__32290),
            .I(N__32284));
    Odrv4 I__7358 (
            .O(N__32287),
            .I(\Commands_frame_decoder.state_ns_i_a3_1_0_0 ));
    LocalMux I__7357 (
            .O(N__32284),
            .I(\Commands_frame_decoder.state_ns_i_a3_1_0_0 ));
    CascadeMux I__7356 (
            .O(N__32279),
            .I(N__32275));
    InMux I__7355 (
            .O(N__32278),
            .I(N__32271));
    InMux I__7354 (
            .O(N__32275),
            .I(N__32266));
    InMux I__7353 (
            .O(N__32274),
            .I(N__32266));
    LocalMux I__7352 (
            .O(N__32271),
            .I(\uart_drone.N_126_li ));
    LocalMux I__7351 (
            .O(N__32266),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__7350 (
            .O(N__32261),
            .I(N__32255));
    CascadeMux I__7349 (
            .O(N__32260),
            .I(N__32252));
    InMux I__7348 (
            .O(N__32259),
            .I(N__32243));
    InMux I__7347 (
            .O(N__32258),
            .I(N__32243));
    InMux I__7346 (
            .O(N__32255),
            .I(N__32243));
    InMux I__7345 (
            .O(N__32252),
            .I(N__32243));
    LocalMux I__7344 (
            .O(N__32243),
            .I(N__32239));
    InMux I__7343 (
            .O(N__32242),
            .I(N__32236));
    Odrv4 I__7342 (
            .O(N__32239),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__7341 (
            .O(N__32236),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__7340 (
            .O(N__32231),
            .I(\uart_drone.N_143_cascade_ ));
    InMux I__7339 (
            .O(N__32228),
            .I(N__32225));
    LocalMux I__7338 (
            .O(N__32225),
            .I(N__32222));
    Odrv12 I__7337 (
            .O(N__32222),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__7336 (
            .O(N__32219),
            .I(N__32216));
    LocalMux I__7335 (
            .O(N__32216),
            .I(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ));
    CascadeMux I__7334 (
            .O(N__32213),
            .I(N__32210));
    InMux I__7333 (
            .O(N__32210),
            .I(N__32207));
    LocalMux I__7332 (
            .O(N__32207),
            .I(N__32203));
    CascadeMux I__7331 (
            .O(N__32206),
            .I(N__32200));
    Span4Mux_h I__7330 (
            .O(N__32203),
            .I(N__32197));
    InMux I__7329 (
            .O(N__32200),
            .I(N__32194));
    Odrv4 I__7328 (
            .O(N__32197),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    LocalMux I__7327 (
            .O(N__32194),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    InMux I__7326 (
            .O(N__32189),
            .I(N__32179));
    InMux I__7325 (
            .O(N__32188),
            .I(N__32179));
    InMux I__7324 (
            .O(N__32187),
            .I(N__32179));
    InMux I__7323 (
            .O(N__32186),
            .I(N__32175));
    LocalMux I__7322 (
            .O(N__32179),
            .I(N__32171));
    InMux I__7321 (
            .O(N__32178),
            .I(N__32168));
    LocalMux I__7320 (
            .O(N__32175),
            .I(N__32165));
    InMux I__7319 (
            .O(N__32174),
            .I(N__32162));
    Span4Mux_h I__7318 (
            .O(N__32171),
            .I(N__32157));
    LocalMux I__7317 (
            .O(N__32168),
            .I(N__32154));
    Span4Mux_v I__7316 (
            .O(N__32165),
            .I(N__32149));
    LocalMux I__7315 (
            .O(N__32162),
            .I(N__32149));
    InMux I__7314 (
            .O(N__32161),
            .I(N__32146));
    InMux I__7313 (
            .O(N__32160),
            .I(N__32143));
    Span4Mux_v I__7312 (
            .O(N__32157),
            .I(N__32140));
    Span4Mux_v I__7311 (
            .O(N__32154),
            .I(N__32135));
    Span4Mux_h I__7310 (
            .O(N__32149),
            .I(N__32135));
    LocalMux I__7309 (
            .O(N__32146),
            .I(N__32132));
    LocalMux I__7308 (
            .O(N__32143),
            .I(N__32129));
    Odrv4 I__7307 (
            .O(N__32140),
            .I(\dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ));
    Odrv4 I__7306 (
            .O(N__32135),
            .I(\dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ));
    Odrv12 I__7305 (
            .O(N__32132),
            .I(\dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ));
    Odrv4 I__7304 (
            .O(N__32129),
            .I(\dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ));
    CascadeMux I__7303 (
            .O(N__32120),
            .I(N__32117));
    InMux I__7302 (
            .O(N__32117),
            .I(N__32114));
    LocalMux I__7301 (
            .O(N__32114),
            .I(N__32111));
    Span4Mux_h I__7300 (
            .O(N__32111),
            .I(N__32108));
    Span4Mux_v I__7299 (
            .O(N__32108),
            .I(N__32104));
    InMux I__7298 (
            .O(N__32107),
            .I(N__32101));
    Odrv4 I__7297 (
            .O(N__32104),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__7296 (
            .O(N__32101),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    InMux I__7295 (
            .O(N__32096),
            .I(N__32093));
    LocalMux I__7294 (
            .O(N__32093),
            .I(N__32087));
    InMux I__7293 (
            .O(N__32092),
            .I(N__32084));
    InMux I__7292 (
            .O(N__32091),
            .I(N__32081));
    CascadeMux I__7291 (
            .O(N__32090),
            .I(N__32078));
    Span4Mux_h I__7290 (
            .O(N__32087),
            .I(N__32071));
    LocalMux I__7289 (
            .O(N__32084),
            .I(N__32071));
    LocalMux I__7288 (
            .O(N__32081),
            .I(N__32071));
    InMux I__7287 (
            .O(N__32078),
            .I(N__32068));
    Span4Mux_v I__7286 (
            .O(N__32071),
            .I(N__32063));
    LocalMux I__7285 (
            .O(N__32068),
            .I(N__32063));
    Odrv4 I__7284 (
            .O(N__32063),
            .I(frame_decoder_OFF3data_0));
    InMux I__7283 (
            .O(N__32060),
            .I(N__32056));
    InMux I__7282 (
            .O(N__32059),
            .I(N__32052));
    LocalMux I__7281 (
            .O(N__32056),
            .I(N__32049));
    InMux I__7280 (
            .O(N__32055),
            .I(N__32046));
    LocalMux I__7279 (
            .O(N__32052),
            .I(N__32038));
    Span4Mux_h I__7278 (
            .O(N__32049),
            .I(N__32038));
    LocalMux I__7277 (
            .O(N__32046),
            .I(N__32038));
    InMux I__7276 (
            .O(N__32045),
            .I(N__32035));
    Span4Mux_v I__7275 (
            .O(N__32038),
            .I(N__32030));
    LocalMux I__7274 (
            .O(N__32035),
            .I(N__32030));
    Odrv4 I__7273 (
            .O(N__32030),
            .I(frame_decoder_CH3data_0));
    InMux I__7272 (
            .O(N__32027),
            .I(N__32023));
    CascadeMux I__7271 (
            .O(N__32026),
            .I(N__32020));
    LocalMux I__7270 (
            .O(N__32023),
            .I(N__32017));
    InMux I__7269 (
            .O(N__32020),
            .I(N__32014));
    Odrv4 I__7268 (
            .O(N__32017),
            .I(scaler_3_data_4));
    LocalMux I__7267 (
            .O(N__32014),
            .I(scaler_3_data_4));
    InMux I__7266 (
            .O(N__32009),
            .I(N__32005));
    InMux I__7265 (
            .O(N__32008),
            .I(N__32002));
    LocalMux I__7264 (
            .O(N__32005),
            .I(N__31999));
    LocalMux I__7263 (
            .O(N__32002),
            .I(N__31996));
    Span4Mux_v I__7262 (
            .O(N__31999),
            .I(N__31991));
    Span4Mux_v I__7261 (
            .O(N__31996),
            .I(N__31991));
    Odrv4 I__7260 (
            .O(N__31991),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa ));
    InMux I__7259 (
            .O(N__31988),
            .I(N__31984));
    InMux I__7258 (
            .O(N__31987),
            .I(N__31981));
    LocalMux I__7257 (
            .O(N__31984),
            .I(N__31978));
    LocalMux I__7256 (
            .O(N__31981),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    Odrv4 I__7255 (
            .O(N__31978),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    InMux I__7254 (
            .O(N__31973),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__7253 (
            .O(N__31970),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__7252 (
            .O(N__31967),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__7251 (
            .O(N__31964),
            .I(N__31960));
    CascadeMux I__7250 (
            .O(N__31963),
            .I(N__31957));
    LocalMux I__7249 (
            .O(N__31960),
            .I(N__31954));
    InMux I__7248 (
            .O(N__31957),
            .I(N__31951));
    Odrv4 I__7247 (
            .O(N__31954),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__7246 (
            .O(N__31951),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    CascadeMux I__7245 (
            .O(N__31946),
            .I(N__31943));
    InMux I__7244 (
            .O(N__31943),
            .I(N__31940));
    LocalMux I__7243 (
            .O(N__31940),
            .I(N__31936));
    InMux I__7242 (
            .O(N__31939),
            .I(N__31933));
    Odrv4 I__7241 (
            .O(N__31936),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__7240 (
            .O(N__31933),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    CEMux I__7239 (
            .O(N__31928),
            .I(N__31925));
    LocalMux I__7238 (
            .O(N__31925),
            .I(N__31922));
    Odrv4 I__7237 (
            .O(N__31922),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    InMux I__7236 (
            .O(N__31919),
            .I(N__31916));
    LocalMux I__7235 (
            .O(N__31916),
            .I(N__31913));
    Odrv4 I__7234 (
            .O(N__31913),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    CascadeMux I__7233 (
            .O(N__31910),
            .I(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ));
    InMux I__7232 (
            .O(N__31907),
            .I(N__31904));
    LocalMux I__7231 (
            .O(N__31904),
            .I(\dron_frame_decoder_1.WDT10lto13_1 ));
    InMux I__7230 (
            .O(N__31901),
            .I(N__31898));
    LocalMux I__7229 (
            .O(N__31898),
            .I(\dron_frame_decoder_1.WDT10lt14_0 ));
    CascadeMux I__7228 (
            .O(N__31895),
            .I(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ));
    InMux I__7227 (
            .O(N__31892),
            .I(N__31889));
    LocalMux I__7226 (
            .O(N__31889),
            .I(N__31886));
    Span4Mux_v I__7225 (
            .O(N__31886),
            .I(N__31883));
    Odrv4 I__7224 (
            .O(N__31883),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    InMux I__7223 (
            .O(N__31880),
            .I(N__31870));
    InMux I__7222 (
            .O(N__31879),
            .I(N__31870));
    CascadeMux I__7221 (
            .O(N__31878),
            .I(N__31867));
    InMux I__7220 (
            .O(N__31877),
            .I(N__31859));
    InMux I__7219 (
            .O(N__31876),
            .I(N__31859));
    InMux I__7218 (
            .O(N__31875),
            .I(N__31859));
    LocalMux I__7217 (
            .O(N__31870),
            .I(N__31856));
    InMux I__7216 (
            .O(N__31867),
            .I(N__31851));
    InMux I__7215 (
            .O(N__31866),
            .I(N__31851));
    LocalMux I__7214 (
            .O(N__31859),
            .I(N__31848));
    Odrv4 I__7213 (
            .O(N__31856),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__7212 (
            .O(N__31851),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    Odrv4 I__7211 (
            .O(N__31848),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__7210 (
            .O(N__31841),
            .I(N__31836));
    InMux I__7209 (
            .O(N__31840),
            .I(N__31830));
    InMux I__7208 (
            .O(N__31839),
            .I(N__31830));
    LocalMux I__7207 (
            .O(N__31836),
            .I(N__31824));
    InMux I__7206 (
            .O(N__31835),
            .I(N__31819));
    LocalMux I__7205 (
            .O(N__31830),
            .I(N__31815));
    InMux I__7204 (
            .O(N__31829),
            .I(N__31812));
    InMux I__7203 (
            .O(N__31828),
            .I(N__31809));
    InMux I__7202 (
            .O(N__31827),
            .I(N__31806));
    Span4Mux_h I__7201 (
            .O(N__31824),
            .I(N__31803));
    InMux I__7200 (
            .O(N__31823),
            .I(N__31799));
    InMux I__7199 (
            .O(N__31822),
            .I(N__31796));
    LocalMux I__7198 (
            .O(N__31819),
            .I(N__31793));
    InMux I__7197 (
            .O(N__31818),
            .I(N__31790));
    Span4Mux_h I__7196 (
            .O(N__31815),
            .I(N__31787));
    LocalMux I__7195 (
            .O(N__31812),
            .I(N__31783));
    LocalMux I__7194 (
            .O(N__31809),
            .I(N__31778));
    LocalMux I__7193 (
            .O(N__31806),
            .I(N__31778));
    Sp12to4 I__7192 (
            .O(N__31803),
            .I(N__31775));
    InMux I__7191 (
            .O(N__31802),
            .I(N__31772));
    LocalMux I__7190 (
            .O(N__31799),
            .I(N__31769));
    LocalMux I__7189 (
            .O(N__31796),
            .I(N__31764));
    Span4Mux_v I__7188 (
            .O(N__31793),
            .I(N__31764));
    LocalMux I__7187 (
            .O(N__31790),
            .I(N__31761));
    Span4Mux_v I__7186 (
            .O(N__31787),
            .I(N__31758));
    InMux I__7185 (
            .O(N__31786),
            .I(N__31755));
    Span12Mux_s9_h I__7184 (
            .O(N__31783),
            .I(N__31752));
    Span12Mux_v I__7183 (
            .O(N__31778),
            .I(N__31747));
    Span12Mux_v I__7182 (
            .O(N__31775),
            .I(N__31747));
    LocalMux I__7181 (
            .O(N__31772),
            .I(N__31736));
    Span4Mux_v I__7180 (
            .O(N__31769),
            .I(N__31736));
    Span4Mux_h I__7179 (
            .O(N__31764),
            .I(N__31736));
    Span4Mux_v I__7178 (
            .O(N__31761),
            .I(N__31736));
    Span4Mux_h I__7177 (
            .O(N__31758),
            .I(N__31736));
    LocalMux I__7176 (
            .O(N__31755),
            .I(uart_pc_data_1));
    Odrv12 I__7175 (
            .O(N__31752),
            .I(uart_pc_data_1));
    Odrv12 I__7174 (
            .O(N__31747),
            .I(uart_pc_data_1));
    Odrv4 I__7173 (
            .O(N__31736),
            .I(uart_pc_data_1));
    InMux I__7172 (
            .O(N__31727),
            .I(N__31716));
    InMux I__7171 (
            .O(N__31726),
            .I(N__31716));
    InMux I__7170 (
            .O(N__31725),
            .I(N__31711));
    InMux I__7169 (
            .O(N__31724),
            .I(N__31711));
    InMux I__7168 (
            .O(N__31723),
            .I(N__31704));
    InMux I__7167 (
            .O(N__31722),
            .I(N__31704));
    InMux I__7166 (
            .O(N__31721),
            .I(N__31704));
    LocalMux I__7165 (
            .O(N__31716),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__7164 (
            .O(N__31711),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__7163 (
            .O(N__31704),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    InMux I__7162 (
            .O(N__31697),
            .I(N__31692));
    InMux I__7161 (
            .O(N__31696),
            .I(N__31686));
    InMux I__7160 (
            .O(N__31695),
            .I(N__31683));
    LocalMux I__7159 (
            .O(N__31692),
            .I(N__31680));
    InMux I__7158 (
            .O(N__31691),
            .I(N__31677));
    InMux I__7157 (
            .O(N__31690),
            .I(N__31674));
    InMux I__7156 (
            .O(N__31689),
            .I(N__31671));
    LocalMux I__7155 (
            .O(N__31686),
            .I(N__31667));
    LocalMux I__7154 (
            .O(N__31683),
            .I(N__31660));
    Span4Mux_h I__7153 (
            .O(N__31680),
            .I(N__31660));
    LocalMux I__7152 (
            .O(N__31677),
            .I(N__31660));
    LocalMux I__7151 (
            .O(N__31674),
            .I(N__31655));
    LocalMux I__7150 (
            .O(N__31671),
            .I(N__31655));
    InMux I__7149 (
            .O(N__31670),
            .I(N__31648));
    Span4Mux_v I__7148 (
            .O(N__31667),
            .I(N__31643));
    Span4Mux_v I__7147 (
            .O(N__31660),
            .I(N__31643));
    Span4Mux_h I__7146 (
            .O(N__31655),
            .I(N__31640));
    InMux I__7145 (
            .O(N__31654),
            .I(N__31637));
    CascadeMux I__7144 (
            .O(N__31653),
            .I(N__31633));
    InMux I__7143 (
            .O(N__31652),
            .I(N__31630));
    InMux I__7142 (
            .O(N__31651),
            .I(N__31627));
    LocalMux I__7141 (
            .O(N__31648),
            .I(N__31624));
    Span4Mux_h I__7140 (
            .O(N__31643),
            .I(N__31619));
    Span4Mux_h I__7139 (
            .O(N__31640),
            .I(N__31619));
    LocalMux I__7138 (
            .O(N__31637),
            .I(N__31616));
    InMux I__7137 (
            .O(N__31636),
            .I(N__31613));
    InMux I__7136 (
            .O(N__31633),
            .I(N__31610));
    LocalMux I__7135 (
            .O(N__31630),
            .I(N__31607));
    LocalMux I__7134 (
            .O(N__31627),
            .I(N__31602));
    Span4Mux_h I__7133 (
            .O(N__31624),
            .I(N__31602));
    Sp12to4 I__7132 (
            .O(N__31619),
            .I(N__31595));
    Span12Mux_s9_h I__7131 (
            .O(N__31616),
            .I(N__31595));
    LocalMux I__7130 (
            .O(N__31613),
            .I(N__31595));
    LocalMux I__7129 (
            .O(N__31610),
            .I(uart_pc_data_4));
    Odrv4 I__7128 (
            .O(N__31607),
            .I(uart_pc_data_4));
    Odrv4 I__7127 (
            .O(N__31602),
            .I(uart_pc_data_4));
    Odrv12 I__7126 (
            .O(N__31595),
            .I(uart_pc_data_4));
    InMux I__7125 (
            .O(N__31586),
            .I(N__31583));
    LocalMux I__7124 (
            .O(N__31583),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__7123 (
            .O(N__31580),
            .I(N__31577));
    LocalMux I__7122 (
            .O(N__31577),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__7121 (
            .O(N__31574),
            .I(N__31571));
    LocalMux I__7120 (
            .O(N__31571),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__7119 (
            .O(N__31568),
            .I(N__31565));
    LocalMux I__7118 (
            .O(N__31565),
            .I(\uart_drone.data_Auxce_0_3 ));
    SRMux I__7117 (
            .O(N__31562),
            .I(N__31559));
    LocalMux I__7116 (
            .O(N__31559),
            .I(N__31556));
    Span4Mux_h I__7115 (
            .O(N__31556),
            .I(N__31552));
    InMux I__7114 (
            .O(N__31555),
            .I(N__31549));
    Odrv4 I__7113 (
            .O(N__31552),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    LocalMux I__7112 (
            .O(N__31549),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    InMux I__7111 (
            .O(N__31544),
            .I(N__31541));
    LocalMux I__7110 (
            .O(N__31541),
            .I(N__31536));
    InMux I__7109 (
            .O(N__31540),
            .I(N__31533));
    InMux I__7108 (
            .O(N__31539),
            .I(N__31530));
    Span4Mux_v I__7107 (
            .O(N__31536),
            .I(N__31523));
    LocalMux I__7106 (
            .O(N__31533),
            .I(N__31523));
    LocalMux I__7105 (
            .O(N__31530),
            .I(N__31523));
    Odrv4 I__7104 (
            .O(N__31523),
            .I(\uart_drone.data_rdyc_1 ));
    CEMux I__7103 (
            .O(N__31520),
            .I(N__31517));
    LocalMux I__7102 (
            .O(N__31517),
            .I(N__31514));
    Odrv12 I__7101 (
            .O(N__31514),
            .I(\uart_drone.data_rdyc_1_0 ));
    InMux I__7100 (
            .O(N__31511),
            .I(N__31507));
    InMux I__7099 (
            .O(N__31510),
            .I(N__31504));
    LocalMux I__7098 (
            .O(N__31507),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__7097 (
            .O(N__31504),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__7096 (
            .O(N__31499),
            .I(N__31495));
    InMux I__7095 (
            .O(N__31498),
            .I(N__31487));
    LocalMux I__7094 (
            .O(N__31495),
            .I(N__31484));
    InMux I__7093 (
            .O(N__31494),
            .I(N__31481));
    InMux I__7092 (
            .O(N__31493),
            .I(N__31478));
    InMux I__7091 (
            .O(N__31492),
            .I(N__31471));
    InMux I__7090 (
            .O(N__31491),
            .I(N__31468));
    InMux I__7089 (
            .O(N__31490),
            .I(N__31465));
    LocalMux I__7088 (
            .O(N__31487),
            .I(N__31462));
    Span4Mux_h I__7087 (
            .O(N__31484),
            .I(N__31459));
    LocalMux I__7086 (
            .O(N__31481),
            .I(N__31456));
    LocalMux I__7085 (
            .O(N__31478),
            .I(N__31453));
    CascadeMux I__7084 (
            .O(N__31477),
            .I(N__31450));
    CascadeMux I__7083 (
            .O(N__31476),
            .I(N__31446));
    InMux I__7082 (
            .O(N__31475),
            .I(N__31442));
    InMux I__7081 (
            .O(N__31474),
            .I(N__31439));
    LocalMux I__7080 (
            .O(N__31471),
            .I(N__31432));
    LocalMux I__7079 (
            .O(N__31468),
            .I(N__31432));
    LocalMux I__7078 (
            .O(N__31465),
            .I(N__31432));
    Span4Mux_h I__7077 (
            .O(N__31462),
            .I(N__31427));
    Span4Mux_v I__7076 (
            .O(N__31459),
            .I(N__31427));
    Span4Mux_h I__7075 (
            .O(N__31456),
            .I(N__31422));
    Span4Mux_h I__7074 (
            .O(N__31453),
            .I(N__31422));
    InMux I__7073 (
            .O(N__31450),
            .I(N__31419));
    InMux I__7072 (
            .O(N__31449),
            .I(N__31416));
    InMux I__7071 (
            .O(N__31446),
            .I(N__31410));
    InMux I__7070 (
            .O(N__31445),
            .I(N__31410));
    LocalMux I__7069 (
            .O(N__31442),
            .I(N__31399));
    LocalMux I__7068 (
            .O(N__31439),
            .I(N__31399));
    Span4Mux_v I__7067 (
            .O(N__31432),
            .I(N__31399));
    Span4Mux_v I__7066 (
            .O(N__31427),
            .I(N__31399));
    Span4Mux_v I__7065 (
            .O(N__31422),
            .I(N__31399));
    LocalMux I__7064 (
            .O(N__31419),
            .I(N__31396));
    LocalMux I__7063 (
            .O(N__31416),
            .I(N__31393));
    InMux I__7062 (
            .O(N__31415),
            .I(N__31390));
    LocalMux I__7061 (
            .O(N__31410),
            .I(N__31387));
    Span4Mux_h I__7060 (
            .O(N__31399),
            .I(N__31380));
    Span4Mux_v I__7059 (
            .O(N__31396),
            .I(N__31380));
    Span4Mux_v I__7058 (
            .O(N__31393),
            .I(N__31380));
    LocalMux I__7057 (
            .O(N__31390),
            .I(uart_pc_data_0));
    Odrv4 I__7056 (
            .O(N__31387),
            .I(uart_pc_data_0));
    Odrv4 I__7055 (
            .O(N__31380),
            .I(uart_pc_data_0));
    InMux I__7054 (
            .O(N__31373),
            .I(N__31370));
    LocalMux I__7053 (
            .O(N__31370),
            .I(N__31366));
    InMux I__7052 (
            .O(N__31369),
            .I(N__31363));
    Span4Mux_h I__7051 (
            .O(N__31366),
            .I(N__31353));
    LocalMux I__7050 (
            .O(N__31363),
            .I(N__31350));
    InMux I__7049 (
            .O(N__31362),
            .I(N__31347));
    InMux I__7048 (
            .O(N__31361),
            .I(N__31344));
    InMux I__7047 (
            .O(N__31360),
            .I(N__31340));
    InMux I__7046 (
            .O(N__31359),
            .I(N__31337));
    InMux I__7045 (
            .O(N__31358),
            .I(N__31334));
    InMux I__7044 (
            .O(N__31357),
            .I(N__31331));
    InMux I__7043 (
            .O(N__31356),
            .I(N__31328));
    Span4Mux_v I__7042 (
            .O(N__31353),
            .I(N__31323));
    Span4Mux_h I__7041 (
            .O(N__31350),
            .I(N__31323));
    LocalMux I__7040 (
            .O(N__31347),
            .I(N__31318));
    LocalMux I__7039 (
            .O(N__31344),
            .I(N__31318));
    InMux I__7038 (
            .O(N__31343),
            .I(N__31315));
    LocalMux I__7037 (
            .O(N__31340),
            .I(N__31312));
    LocalMux I__7036 (
            .O(N__31337),
            .I(N__31308));
    LocalMux I__7035 (
            .O(N__31334),
            .I(N__31304));
    LocalMux I__7034 (
            .O(N__31331),
            .I(N__31299));
    LocalMux I__7033 (
            .O(N__31328),
            .I(N__31299));
    Span4Mux_v I__7032 (
            .O(N__31323),
            .I(N__31296));
    Span4Mux_v I__7031 (
            .O(N__31318),
            .I(N__31291));
    LocalMux I__7030 (
            .O(N__31315),
            .I(N__31291));
    Span4Mux_h I__7029 (
            .O(N__31312),
            .I(N__31288));
    InMux I__7028 (
            .O(N__31311),
            .I(N__31285));
    Span12Mux_s9_h I__7027 (
            .O(N__31308),
            .I(N__31282));
    InMux I__7026 (
            .O(N__31307),
            .I(N__31279));
    Span4Mux_h I__7025 (
            .O(N__31304),
            .I(N__31272));
    Span4Mux_v I__7024 (
            .O(N__31299),
            .I(N__31272));
    Span4Mux_h I__7023 (
            .O(N__31296),
            .I(N__31272));
    Span4Mux_h I__7022 (
            .O(N__31291),
            .I(N__31265));
    Span4Mux_h I__7021 (
            .O(N__31288),
            .I(N__31265));
    LocalMux I__7020 (
            .O(N__31285),
            .I(N__31265));
    Odrv12 I__7019 (
            .O(N__31282),
            .I(uart_pc_data_6));
    LocalMux I__7018 (
            .O(N__31279),
            .I(uart_pc_data_6));
    Odrv4 I__7017 (
            .O(N__31272),
            .I(uart_pc_data_6));
    Odrv4 I__7016 (
            .O(N__31265),
            .I(uart_pc_data_6));
    CascadeMux I__7015 (
            .O(N__31256),
            .I(N__31251));
    InMux I__7014 (
            .O(N__31255),
            .I(N__31248));
    InMux I__7013 (
            .O(N__31254),
            .I(N__31243));
    InMux I__7012 (
            .O(N__31251),
            .I(N__31243));
    LocalMux I__7011 (
            .O(N__31248),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__7010 (
            .O(N__31243),
            .I(\uart_drone.stateZ0Z_1 ));
    CascadeMux I__7009 (
            .O(N__31238),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__7008 (
            .O(N__31235),
            .I(N__31232));
    LocalMux I__7007 (
            .O(N__31232),
            .I(N__31229));
    Span4Mux_v I__7006 (
            .O(N__31229),
            .I(N__31226));
    Odrv4 I__7005 (
            .O(N__31226),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    InMux I__7004 (
            .O(N__31223),
            .I(N__31217));
    InMux I__7003 (
            .O(N__31222),
            .I(N__31214));
    CascadeMux I__7002 (
            .O(N__31221),
            .I(N__31211));
    InMux I__7001 (
            .O(N__31220),
            .I(N__31206));
    LocalMux I__7000 (
            .O(N__31217),
            .I(N__31203));
    LocalMux I__6999 (
            .O(N__31214),
            .I(N__31196));
    InMux I__6998 (
            .O(N__31211),
            .I(N__31191));
    InMux I__6997 (
            .O(N__31210),
            .I(N__31191));
    InMux I__6996 (
            .O(N__31209),
            .I(N__31188));
    LocalMux I__6995 (
            .O(N__31206),
            .I(N__31185));
    Span4Mux_v I__6994 (
            .O(N__31203),
            .I(N__31182));
    InMux I__6993 (
            .O(N__31202),
            .I(N__31179));
    InMux I__6992 (
            .O(N__31201),
            .I(N__31176));
    InMux I__6991 (
            .O(N__31200),
            .I(N__31173));
    InMux I__6990 (
            .O(N__31199),
            .I(N__31170));
    Span4Mux_v I__6989 (
            .O(N__31196),
            .I(N__31165));
    LocalMux I__6988 (
            .O(N__31191),
            .I(N__31165));
    LocalMux I__6987 (
            .O(N__31188),
            .I(N__31162));
    Span4Mux_h I__6986 (
            .O(N__31185),
            .I(N__31159));
    Span4Mux_v I__6985 (
            .O(N__31182),
            .I(N__31149));
    LocalMux I__6984 (
            .O(N__31179),
            .I(N__31149));
    LocalMux I__6983 (
            .O(N__31176),
            .I(N__31149));
    LocalMux I__6982 (
            .O(N__31173),
            .I(N__31149));
    LocalMux I__6981 (
            .O(N__31170),
            .I(N__31144));
    Span4Mux_v I__6980 (
            .O(N__31165),
            .I(N__31144));
    Span4Mux_v I__6979 (
            .O(N__31162),
            .I(N__31138));
    Span4Mux_v I__6978 (
            .O(N__31159),
            .I(N__31138));
    InMux I__6977 (
            .O(N__31158),
            .I(N__31135));
    Span4Mux_v I__6976 (
            .O(N__31149),
            .I(N__31130));
    Span4Mux_v I__6975 (
            .O(N__31144),
            .I(N__31130));
    InMux I__6974 (
            .O(N__31143),
            .I(N__31127));
    Span4Mux_h I__6973 (
            .O(N__31138),
            .I(N__31124));
    LocalMux I__6972 (
            .O(N__31135),
            .I(N__31121));
    Sp12to4 I__6971 (
            .O(N__31130),
            .I(N__31118));
    LocalMux I__6970 (
            .O(N__31127),
            .I(uart_pc_data_3));
    Odrv4 I__6969 (
            .O(N__31124),
            .I(uart_pc_data_3));
    Odrv12 I__6968 (
            .O(N__31121),
            .I(uart_pc_data_3));
    Odrv12 I__6967 (
            .O(N__31118),
            .I(uart_pc_data_3));
    CascadeMux I__6966 (
            .O(N__31109),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ));
    InMux I__6965 (
            .O(N__31106),
            .I(N__31103));
    LocalMux I__6964 (
            .O(N__31103),
            .I(N__31098));
    InMux I__6963 (
            .O(N__31102),
            .I(N__31093));
    InMux I__6962 (
            .O(N__31101),
            .I(N__31093));
    Odrv4 I__6961 (
            .O(N__31098),
            .I(\Commands_frame_decoder.N_342 ));
    LocalMux I__6960 (
            .O(N__31093),
            .I(\Commands_frame_decoder.N_342 ));
    InMux I__6959 (
            .O(N__31088),
            .I(N__31085));
    LocalMux I__6958 (
            .O(N__31085),
            .I(N__31080));
    InMux I__6957 (
            .O(N__31084),
            .I(N__31073));
    InMux I__6956 (
            .O(N__31083),
            .I(N__31073));
    Span4Mux_h I__6955 (
            .O(N__31080),
            .I(N__31070));
    InMux I__6954 (
            .O(N__31079),
            .I(N__31067));
    InMux I__6953 (
            .O(N__31078),
            .I(N__31064));
    LocalMux I__6952 (
            .O(N__31073),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    Odrv4 I__6951 (
            .O(N__31070),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__6950 (
            .O(N__31067),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__6949 (
            .O(N__31064),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    InMux I__6948 (
            .O(N__31055),
            .I(N__31052));
    LocalMux I__6947 (
            .O(N__31052),
            .I(N__31049));
    Odrv4 I__6946 (
            .O(N__31049),
            .I(\Commands_frame_decoder.N_308_2 ));
    InMux I__6945 (
            .O(N__31046),
            .I(N__31042));
    InMux I__6944 (
            .O(N__31045),
            .I(N__31039));
    LocalMux I__6943 (
            .O(N__31042),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    LocalMux I__6942 (
            .O(N__31039),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    CascadeMux I__6941 (
            .O(N__31034),
            .I(\Commands_frame_decoder.N_308_2_cascade_ ));
    InMux I__6940 (
            .O(N__31031),
            .I(N__31028));
    LocalMux I__6939 (
            .O(N__31028),
            .I(\Commands_frame_decoder.state_ns_i_1_0 ));
    CascadeMux I__6938 (
            .O(N__31025),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__6937 (
            .O(N__31022),
            .I(N__31019));
    LocalMux I__6936 (
            .O(N__31019),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__6935 (
            .O(N__31016),
            .I(N__31013));
    LocalMux I__6934 (
            .O(N__31013),
            .I(N__31010));
    Odrv4 I__6933 (
            .O(N__31010),
            .I(uart_input_pc_c));
    InMux I__6932 (
            .O(N__31007),
            .I(N__31004));
    LocalMux I__6931 (
            .O(N__31004),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    CascadeMux I__6930 (
            .O(N__31001),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ));
    InMux I__6929 (
            .O(N__30998),
            .I(N__30995));
    LocalMux I__6928 (
            .O(N__30995),
            .I(\Commands_frame_decoder.N_338 ));
    CascadeMux I__6927 (
            .O(N__30992),
            .I(\Commands_frame_decoder.N_309_cascade_ ));
    InMux I__6926 (
            .O(N__30989),
            .I(N__30984));
    InMux I__6925 (
            .O(N__30988),
            .I(N__30978));
    InMux I__6924 (
            .O(N__30987),
            .I(N__30975));
    LocalMux I__6923 (
            .O(N__30984),
            .I(N__30970));
    InMux I__6922 (
            .O(N__30983),
            .I(N__30966));
    InMux I__6921 (
            .O(N__30982),
            .I(N__30963));
    InMux I__6920 (
            .O(N__30981),
            .I(N__30960));
    LocalMux I__6919 (
            .O(N__30978),
            .I(N__30954));
    LocalMux I__6918 (
            .O(N__30975),
            .I(N__30951));
    InMux I__6917 (
            .O(N__30974),
            .I(N__30946));
    InMux I__6916 (
            .O(N__30973),
            .I(N__30946));
    Span4Mux_v I__6915 (
            .O(N__30970),
            .I(N__30942));
    InMux I__6914 (
            .O(N__30969),
            .I(N__30939));
    LocalMux I__6913 (
            .O(N__30966),
            .I(N__30934));
    LocalMux I__6912 (
            .O(N__30963),
            .I(N__30934));
    LocalMux I__6911 (
            .O(N__30960),
            .I(N__30931));
    InMux I__6910 (
            .O(N__30959),
            .I(N__30928));
    InMux I__6909 (
            .O(N__30958),
            .I(N__30925));
    InMux I__6908 (
            .O(N__30957),
            .I(N__30922));
    Span4Mux_v I__6907 (
            .O(N__30954),
            .I(N__30916));
    Span4Mux_v I__6906 (
            .O(N__30951),
            .I(N__30916));
    LocalMux I__6905 (
            .O(N__30946),
            .I(N__30913));
    InMux I__6904 (
            .O(N__30945),
            .I(N__30910));
    Span4Mux_v I__6903 (
            .O(N__30942),
            .I(N__30905));
    LocalMux I__6902 (
            .O(N__30939),
            .I(N__30905));
    Span4Mux_v I__6901 (
            .O(N__30934),
            .I(N__30902));
    Span4Mux_v I__6900 (
            .O(N__30931),
            .I(N__30897));
    LocalMux I__6899 (
            .O(N__30928),
            .I(N__30897));
    LocalMux I__6898 (
            .O(N__30925),
            .I(N__30892));
    LocalMux I__6897 (
            .O(N__30922),
            .I(N__30892));
    InMux I__6896 (
            .O(N__30921),
            .I(N__30889));
    Span4Mux_h I__6895 (
            .O(N__30916),
            .I(N__30880));
    Span4Mux_h I__6894 (
            .O(N__30913),
            .I(N__30880));
    LocalMux I__6893 (
            .O(N__30910),
            .I(N__30880));
    Span4Mux_h I__6892 (
            .O(N__30905),
            .I(N__30880));
    Odrv4 I__6891 (
            .O(N__30902),
            .I(uart_pc_data_7));
    Odrv4 I__6890 (
            .O(N__30897),
            .I(uart_pc_data_7));
    Odrv12 I__6889 (
            .O(N__30892),
            .I(uart_pc_data_7));
    LocalMux I__6888 (
            .O(N__30889),
            .I(uart_pc_data_7));
    Odrv4 I__6887 (
            .O(N__30880),
            .I(uart_pc_data_7));
    InMux I__6886 (
            .O(N__30869),
            .I(N__30864));
    InMux I__6885 (
            .O(N__30868),
            .I(N__30861));
    InMux I__6884 (
            .O(N__30867),
            .I(N__30858));
    LocalMux I__6883 (
            .O(N__30864),
            .I(N__30847));
    LocalMux I__6882 (
            .O(N__30861),
            .I(N__30847));
    LocalMux I__6881 (
            .O(N__30858),
            .I(N__30841));
    InMux I__6880 (
            .O(N__30857),
            .I(N__30838));
    InMux I__6879 (
            .O(N__30856),
            .I(N__30835));
    InMux I__6878 (
            .O(N__30855),
            .I(N__30829));
    InMux I__6877 (
            .O(N__30854),
            .I(N__30829));
    InMux I__6876 (
            .O(N__30853),
            .I(N__30825));
    InMux I__6875 (
            .O(N__30852),
            .I(N__30822));
    Span4Mux_v I__6874 (
            .O(N__30847),
            .I(N__30818));
    InMux I__6873 (
            .O(N__30846),
            .I(N__30813));
    InMux I__6872 (
            .O(N__30845),
            .I(N__30813));
    InMux I__6871 (
            .O(N__30844),
            .I(N__30810));
    Span4Mux_h I__6870 (
            .O(N__30841),
            .I(N__30805));
    LocalMux I__6869 (
            .O(N__30838),
            .I(N__30805));
    LocalMux I__6868 (
            .O(N__30835),
            .I(N__30802));
    InMux I__6867 (
            .O(N__30834),
            .I(N__30799));
    LocalMux I__6866 (
            .O(N__30829),
            .I(N__30796));
    InMux I__6865 (
            .O(N__30828),
            .I(N__30793));
    LocalMux I__6864 (
            .O(N__30825),
            .I(N__30788));
    LocalMux I__6863 (
            .O(N__30822),
            .I(N__30788));
    InMux I__6862 (
            .O(N__30821),
            .I(N__30785));
    Sp12to4 I__6861 (
            .O(N__30818),
            .I(N__30780));
    LocalMux I__6860 (
            .O(N__30813),
            .I(N__30780));
    LocalMux I__6859 (
            .O(N__30810),
            .I(N__30777));
    Span4Mux_h I__6858 (
            .O(N__30805),
            .I(N__30768));
    Span4Mux_h I__6857 (
            .O(N__30802),
            .I(N__30768));
    LocalMux I__6856 (
            .O(N__30799),
            .I(N__30768));
    Span4Mux_v I__6855 (
            .O(N__30796),
            .I(N__30768));
    LocalMux I__6854 (
            .O(N__30793),
            .I(N__30759));
    Sp12to4 I__6853 (
            .O(N__30788),
            .I(N__30759));
    LocalMux I__6852 (
            .O(N__30785),
            .I(N__30759));
    Span12Mux_s8_h I__6851 (
            .O(N__30780),
            .I(N__30759));
    Odrv4 I__6850 (
            .O(N__30777),
            .I(uart_pc_data_2));
    Odrv4 I__6849 (
            .O(N__30768),
            .I(uart_pc_data_2));
    Odrv12 I__6848 (
            .O(N__30759),
            .I(uart_pc_data_2));
    CascadeMux I__6847 (
            .O(N__30752),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ));
    InMux I__6846 (
            .O(N__30749),
            .I(N__30746));
    LocalMux I__6845 (
            .O(N__30746),
            .I(N__30742));
    InMux I__6844 (
            .O(N__30745),
            .I(N__30739));
    Span4Mux_v I__6843 (
            .O(N__30742),
            .I(N__30731));
    LocalMux I__6842 (
            .O(N__30739),
            .I(N__30731));
    InMux I__6841 (
            .O(N__30738),
            .I(N__30725));
    InMux I__6840 (
            .O(N__30737),
            .I(N__30721));
    InMux I__6839 (
            .O(N__30736),
            .I(N__30718));
    Span4Mux_v I__6838 (
            .O(N__30731),
            .I(N__30712));
    InMux I__6837 (
            .O(N__30730),
            .I(N__30706));
    InMux I__6836 (
            .O(N__30729),
            .I(N__30706));
    InMux I__6835 (
            .O(N__30728),
            .I(N__30703));
    LocalMux I__6834 (
            .O(N__30725),
            .I(N__30700));
    InMux I__6833 (
            .O(N__30724),
            .I(N__30697));
    LocalMux I__6832 (
            .O(N__30721),
            .I(N__30692));
    LocalMux I__6831 (
            .O(N__30718),
            .I(N__30692));
    InMux I__6830 (
            .O(N__30717),
            .I(N__30689));
    InMux I__6829 (
            .O(N__30716),
            .I(N__30686));
    InMux I__6828 (
            .O(N__30715),
            .I(N__30683));
    Span4Mux_v I__6827 (
            .O(N__30712),
            .I(N__30679));
    InMux I__6826 (
            .O(N__30711),
            .I(N__30676));
    LocalMux I__6825 (
            .O(N__30706),
            .I(N__30673));
    LocalMux I__6824 (
            .O(N__30703),
            .I(N__30670));
    Span4Mux_h I__6823 (
            .O(N__30700),
            .I(N__30667));
    LocalMux I__6822 (
            .O(N__30697),
            .I(N__30664));
    Span4Mux_h I__6821 (
            .O(N__30692),
            .I(N__30655));
    LocalMux I__6820 (
            .O(N__30689),
            .I(N__30655));
    LocalMux I__6819 (
            .O(N__30686),
            .I(N__30655));
    LocalMux I__6818 (
            .O(N__30683),
            .I(N__30655));
    InMux I__6817 (
            .O(N__30682),
            .I(N__30652));
    Span4Mux_h I__6816 (
            .O(N__30679),
            .I(N__30649));
    LocalMux I__6815 (
            .O(N__30676),
            .I(N__30642));
    Span4Mux_h I__6814 (
            .O(N__30673),
            .I(N__30642));
    Span4Mux_h I__6813 (
            .O(N__30670),
            .I(N__30642));
    Odrv4 I__6812 (
            .O(N__30667),
            .I(uart_pc_data_5));
    Odrv12 I__6811 (
            .O(N__30664),
            .I(uart_pc_data_5));
    Odrv4 I__6810 (
            .O(N__30655),
            .I(uart_pc_data_5));
    LocalMux I__6809 (
            .O(N__30652),
            .I(uart_pc_data_5));
    Odrv4 I__6808 (
            .O(N__30649),
            .I(uart_pc_data_5));
    Odrv4 I__6807 (
            .O(N__30642),
            .I(uart_pc_data_5));
    CascadeMux I__6806 (
            .O(N__30629),
            .I(\Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ));
    CascadeMux I__6805 (
            .O(N__30626),
            .I(N__30622));
    InMux I__6804 (
            .O(N__30625),
            .I(N__30619));
    InMux I__6803 (
            .O(N__30622),
            .I(N__30615));
    LocalMux I__6802 (
            .O(N__30619),
            .I(N__30612));
    CascadeMux I__6801 (
            .O(N__30618),
            .I(N__30609));
    LocalMux I__6800 (
            .O(N__30615),
            .I(N__30602));
    Span4Mux_h I__6799 (
            .O(N__30612),
            .I(N__30602));
    InMux I__6798 (
            .O(N__30609),
            .I(N__30599));
    InMux I__6797 (
            .O(N__30608),
            .I(N__30594));
    InMux I__6796 (
            .O(N__30607),
            .I(N__30594));
    Span4Mux_v I__6795 (
            .O(N__30602),
            .I(N__30591));
    LocalMux I__6794 (
            .O(N__30599),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    LocalMux I__6793 (
            .O(N__30594),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__6792 (
            .O(N__30591),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    CascadeMux I__6791 (
            .O(N__30584),
            .I(N__30580));
    CascadeMux I__6790 (
            .O(N__30583),
            .I(N__30576));
    InMux I__6789 (
            .O(N__30580),
            .I(N__30572));
    CascadeMux I__6788 (
            .O(N__30579),
            .I(N__30564));
    InMux I__6787 (
            .O(N__30576),
            .I(N__30559));
    InMux I__6786 (
            .O(N__30575),
            .I(N__30559));
    LocalMux I__6785 (
            .O(N__30572),
            .I(N__30554));
    InMux I__6784 (
            .O(N__30571),
            .I(N__30551));
    InMux I__6783 (
            .O(N__30570),
            .I(N__30546));
    InMux I__6782 (
            .O(N__30569),
            .I(N__30546));
    InMux I__6781 (
            .O(N__30568),
            .I(N__30540));
    InMux I__6780 (
            .O(N__30567),
            .I(N__30540));
    InMux I__6779 (
            .O(N__30564),
            .I(N__30537));
    LocalMux I__6778 (
            .O(N__30559),
            .I(N__30534));
    InMux I__6777 (
            .O(N__30558),
            .I(N__30526));
    InMux I__6776 (
            .O(N__30557),
            .I(N__30526));
    Span4Mux_s2_v I__6775 (
            .O(N__30554),
            .I(N__30523));
    LocalMux I__6774 (
            .O(N__30551),
            .I(N__30520));
    LocalMux I__6773 (
            .O(N__30546),
            .I(N__30517));
    InMux I__6772 (
            .O(N__30545),
            .I(N__30514));
    LocalMux I__6771 (
            .O(N__30540),
            .I(N__30511));
    LocalMux I__6770 (
            .O(N__30537),
            .I(N__30506));
    Span4Mux_s2_h I__6769 (
            .O(N__30534),
            .I(N__30506));
    InMux I__6768 (
            .O(N__30533),
            .I(N__30501));
    InMux I__6767 (
            .O(N__30532),
            .I(N__30501));
    InMux I__6766 (
            .O(N__30531),
            .I(N__30498));
    LocalMux I__6765 (
            .O(N__30526),
            .I(N__30495));
    Sp12to4 I__6764 (
            .O(N__30523),
            .I(N__30490));
    Span12Mux_v I__6763 (
            .O(N__30520),
            .I(N__30490));
    Span4Mux_h I__6762 (
            .O(N__30517),
            .I(N__30487));
    LocalMux I__6761 (
            .O(N__30514),
            .I(N__30482));
    Span4Mux_v I__6760 (
            .O(N__30511),
            .I(N__30482));
    Span4Mux_h I__6759 (
            .O(N__30506),
            .I(N__30479));
    LocalMux I__6758 (
            .O(N__30501),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__6757 (
            .O(N__30498),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv12 I__6756 (
            .O(N__30495),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv12 I__6755 (
            .O(N__30490),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__6754 (
            .O(N__30487),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__6753 (
            .O(N__30482),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__6752 (
            .O(N__30479),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    InMux I__6751 (
            .O(N__30464),
            .I(N__30461));
    LocalMux I__6750 (
            .O(N__30461),
            .I(N__30458));
    Span4Mux_h I__6749 (
            .O(N__30458),
            .I(N__30455));
    Odrv4 I__6748 (
            .O(N__30455),
            .I(\ppm_encoder_1.N_320 ));
    InMux I__6747 (
            .O(N__30452),
            .I(N__30449));
    LocalMux I__6746 (
            .O(N__30449),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    InMux I__6745 (
            .O(N__30446),
            .I(N__30443));
    LocalMux I__6744 (
            .O(N__30443),
            .I(N__30440));
    Odrv4 I__6743 (
            .O(N__30440),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    InMux I__6742 (
            .O(N__30437),
            .I(N__30434));
    LocalMux I__6741 (
            .O(N__30434),
            .I(N__30430));
    InMux I__6740 (
            .O(N__30433),
            .I(N__30426));
    Span4Mux_h I__6739 (
            .O(N__30430),
            .I(N__30423));
    InMux I__6738 (
            .O(N__30429),
            .I(N__30420));
    LocalMux I__6737 (
            .O(N__30426),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__6736 (
            .O(N__30423),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__6735 (
            .O(N__30420),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    CascadeMux I__6734 (
            .O(N__30413),
            .I(N__30410));
    InMux I__6733 (
            .O(N__30410),
            .I(N__30407));
    LocalMux I__6732 (
            .O(N__30407),
            .I(N__30404));
    Odrv12 I__6731 (
            .O(N__30404),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__6730 (
            .O(N__30401),
            .I(N__30398));
    LocalMux I__6729 (
            .O(N__30398),
            .I(N__30395));
    Span4Mux_h I__6728 (
            .O(N__30395),
            .I(N__30391));
    InMux I__6727 (
            .O(N__30394),
            .I(N__30387));
    Span4Mux_h I__6726 (
            .O(N__30391),
            .I(N__30384));
    InMux I__6725 (
            .O(N__30390),
            .I(N__30381));
    LocalMux I__6724 (
            .O(N__30387),
            .I(N__30378));
    Odrv4 I__6723 (
            .O(N__30384),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__6722 (
            .O(N__30381),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__6721 (
            .O(N__30378),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__6720 (
            .O(N__30371),
            .I(N__30368));
    LocalMux I__6719 (
            .O(N__30368),
            .I(N__30364));
    InMux I__6718 (
            .O(N__30367),
            .I(N__30361));
    Span4Mux_h I__6717 (
            .O(N__30364),
            .I(N__30358));
    LocalMux I__6716 (
            .O(N__30361),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    Odrv4 I__6715 (
            .O(N__30358),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    InMux I__6714 (
            .O(N__30353),
            .I(N__30350));
    LocalMux I__6713 (
            .O(N__30350),
            .I(N__30347));
    Span4Mux_h I__6712 (
            .O(N__30347),
            .I(N__30344));
    Span4Mux_h I__6711 (
            .O(N__30344),
            .I(N__30339));
    InMux I__6710 (
            .O(N__30343),
            .I(N__30334));
    InMux I__6709 (
            .O(N__30342),
            .I(N__30334));
    Odrv4 I__6708 (
            .O(N__30339),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__6707 (
            .O(N__30334),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__6706 (
            .O(N__30329),
            .I(N__30326));
    InMux I__6705 (
            .O(N__30326),
            .I(N__30323));
    LocalMux I__6704 (
            .O(N__30323),
            .I(N__30319));
    InMux I__6703 (
            .O(N__30322),
            .I(N__30316));
    Span4Mux_s3_v I__6702 (
            .O(N__30319),
            .I(N__30313));
    LocalMux I__6701 (
            .O(N__30316),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    Odrv4 I__6700 (
            .O(N__30313),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__6699 (
            .O(N__30308),
            .I(N__30305));
    LocalMux I__6698 (
            .O(N__30305),
            .I(N__30301));
    InMux I__6697 (
            .O(N__30304),
            .I(N__30298));
    Span4Mux_v I__6696 (
            .O(N__30301),
            .I(N__30295));
    LocalMux I__6695 (
            .O(N__30298),
            .I(N__30291));
    Span4Mux_h I__6694 (
            .O(N__30295),
            .I(N__30288));
    InMux I__6693 (
            .O(N__30294),
            .I(N__30285));
    Span4Mux_v I__6692 (
            .O(N__30291),
            .I(N__30282));
    Odrv4 I__6691 (
            .O(N__30288),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__6690 (
            .O(N__30285),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__6689 (
            .O(N__30282),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    CascadeMux I__6688 (
            .O(N__30275),
            .I(N__30272));
    InMux I__6687 (
            .O(N__30272),
            .I(N__30266));
    InMux I__6686 (
            .O(N__30271),
            .I(N__30266));
    LocalMux I__6685 (
            .O(N__30266),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__6684 (
            .O(N__30263),
            .I(N__30260));
    LocalMux I__6683 (
            .O(N__30260),
            .I(N__30257));
    Span4Mux_h I__6682 (
            .O(N__30257),
            .I(N__30254));
    Odrv4 I__6681 (
            .O(N__30254),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__6680 (
            .O(N__30251),
            .I(N__30246));
    InMux I__6679 (
            .O(N__30250),
            .I(N__30241));
    InMux I__6678 (
            .O(N__30249),
            .I(N__30241));
    LocalMux I__6677 (
            .O(N__30246),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__6676 (
            .O(N__30241),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__6675 (
            .O(N__30236),
            .I(N__30231));
    InMux I__6674 (
            .O(N__30235),
            .I(N__30228));
    InMux I__6673 (
            .O(N__30234),
            .I(N__30225));
    LocalMux I__6672 (
            .O(N__30231),
            .I(N__30222));
    LocalMux I__6671 (
            .O(N__30228),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__6670 (
            .O(N__30225),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__6669 (
            .O(N__30222),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    CascadeMux I__6668 (
            .O(N__30215),
            .I(N__30210));
    InMux I__6667 (
            .O(N__30214),
            .I(N__30207));
    InMux I__6666 (
            .O(N__30213),
            .I(N__30204));
    InMux I__6665 (
            .O(N__30210),
            .I(N__30201));
    LocalMux I__6664 (
            .O(N__30207),
            .I(N__30198));
    LocalMux I__6663 (
            .O(N__30204),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__6662 (
            .O(N__30201),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__6661 (
            .O(N__30198),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__6660 (
            .O(N__30191),
            .I(N__30186));
    InMux I__6659 (
            .O(N__30190),
            .I(N__30181));
    InMux I__6658 (
            .O(N__30189),
            .I(N__30181));
    LocalMux I__6657 (
            .O(N__30186),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__6656 (
            .O(N__30181),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__6655 (
            .O(N__30176),
            .I(N__30170));
    InMux I__6654 (
            .O(N__30175),
            .I(N__30170));
    LocalMux I__6653 (
            .O(N__30170),
            .I(N__30167));
    Span4Mux_v I__6652 (
            .O(N__30167),
            .I(N__30164));
    Odrv4 I__6651 (
            .O(N__30164),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    InMux I__6650 (
            .O(N__30161),
            .I(N__30158));
    LocalMux I__6649 (
            .O(N__30158),
            .I(N__30155));
    Span12Mux_h I__6648 (
            .O(N__30155),
            .I(N__30150));
    InMux I__6647 (
            .O(N__30154),
            .I(N__30145));
    InMux I__6646 (
            .O(N__30153),
            .I(N__30145));
    Odrv12 I__6645 (
            .O(N__30150),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__6644 (
            .O(N__30145),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    CascadeMux I__6643 (
            .O(N__30140),
            .I(N__30134));
    CascadeMux I__6642 (
            .O(N__30139),
            .I(N__30131));
    CascadeMux I__6641 (
            .O(N__30138),
            .I(N__30128));
    InMux I__6640 (
            .O(N__30137),
            .I(N__30121));
    InMux I__6639 (
            .O(N__30134),
            .I(N__30121));
    InMux I__6638 (
            .O(N__30131),
            .I(N__30121));
    InMux I__6637 (
            .O(N__30128),
            .I(N__30118));
    LocalMux I__6636 (
            .O(N__30121),
            .I(N__30113));
    LocalMux I__6635 (
            .O(N__30118),
            .I(N__30113));
    Span12Mux_v I__6634 (
            .O(N__30113),
            .I(N__30109));
    InMux I__6633 (
            .O(N__30112),
            .I(N__30106));
    Odrv12 I__6632 (
            .O(N__30109),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ));
    LocalMux I__6631 (
            .O(N__30106),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ));
    CascadeMux I__6630 (
            .O(N__30101),
            .I(N__30093));
    CascadeMux I__6629 (
            .O(N__30100),
            .I(N__30080));
    InMux I__6628 (
            .O(N__30099),
            .I(N__30077));
    CascadeMux I__6627 (
            .O(N__30098),
            .I(N__30073));
    CascadeMux I__6626 (
            .O(N__30097),
            .I(N__30069));
    CascadeMux I__6625 (
            .O(N__30096),
            .I(N__30066));
    InMux I__6624 (
            .O(N__30093),
            .I(N__30056));
    InMux I__6623 (
            .O(N__30092),
            .I(N__30056));
    InMux I__6622 (
            .O(N__30091),
            .I(N__30056));
    InMux I__6621 (
            .O(N__30090),
            .I(N__30056));
    CascadeMux I__6620 (
            .O(N__30089),
            .I(N__30053));
    CascadeMux I__6619 (
            .O(N__30088),
            .I(N__30032));
    CascadeMux I__6618 (
            .O(N__30087),
            .I(N__30029));
    InMux I__6617 (
            .O(N__30086),
            .I(N__30017));
    InMux I__6616 (
            .O(N__30085),
            .I(N__30017));
    InMux I__6615 (
            .O(N__30084),
            .I(N__30017));
    InMux I__6614 (
            .O(N__30083),
            .I(N__30014));
    InMux I__6613 (
            .O(N__30080),
            .I(N__30011));
    LocalMux I__6612 (
            .O(N__30077),
            .I(N__30008));
    InMux I__6611 (
            .O(N__30076),
            .I(N__30005));
    InMux I__6610 (
            .O(N__30073),
            .I(N__29994));
    InMux I__6609 (
            .O(N__30072),
            .I(N__29994));
    InMux I__6608 (
            .O(N__30069),
            .I(N__29994));
    InMux I__6607 (
            .O(N__30066),
            .I(N__29994));
    InMux I__6606 (
            .O(N__30065),
            .I(N__29994));
    LocalMux I__6605 (
            .O(N__30056),
            .I(N__29991));
    InMux I__6604 (
            .O(N__30053),
            .I(N__29982));
    InMux I__6603 (
            .O(N__30052),
            .I(N__29982));
    InMux I__6602 (
            .O(N__30051),
            .I(N__29982));
    InMux I__6601 (
            .O(N__30050),
            .I(N__29982));
    InMux I__6600 (
            .O(N__30049),
            .I(N__29973));
    InMux I__6599 (
            .O(N__30048),
            .I(N__29973));
    InMux I__6598 (
            .O(N__30047),
            .I(N__29973));
    InMux I__6597 (
            .O(N__30046),
            .I(N__29973));
    InMux I__6596 (
            .O(N__30045),
            .I(N__29968));
    InMux I__6595 (
            .O(N__30044),
            .I(N__29968));
    InMux I__6594 (
            .O(N__30043),
            .I(N__29959));
    InMux I__6593 (
            .O(N__30042),
            .I(N__29952));
    InMux I__6592 (
            .O(N__30041),
            .I(N__29952));
    InMux I__6591 (
            .O(N__30040),
            .I(N__29952));
    InMux I__6590 (
            .O(N__30039),
            .I(N__29945));
    InMux I__6589 (
            .O(N__30038),
            .I(N__29945));
    InMux I__6588 (
            .O(N__30037),
            .I(N__29945));
    InMux I__6587 (
            .O(N__30036),
            .I(N__29940));
    InMux I__6586 (
            .O(N__30035),
            .I(N__29940));
    InMux I__6585 (
            .O(N__30032),
            .I(N__29929));
    InMux I__6584 (
            .O(N__30029),
            .I(N__29929));
    InMux I__6583 (
            .O(N__30028),
            .I(N__29929));
    InMux I__6582 (
            .O(N__30027),
            .I(N__29929));
    InMux I__6581 (
            .O(N__30026),
            .I(N__29929));
    CascadeMux I__6580 (
            .O(N__30025),
            .I(N__29924));
    InMux I__6579 (
            .O(N__30024),
            .I(N__29921));
    LocalMux I__6578 (
            .O(N__30017),
            .I(N__29918));
    LocalMux I__6577 (
            .O(N__30014),
            .I(N__29915));
    LocalMux I__6576 (
            .O(N__30011),
            .I(N__29905));
    Span4Mux_v I__6575 (
            .O(N__30008),
            .I(N__29902));
    LocalMux I__6574 (
            .O(N__30005),
            .I(N__29889));
    LocalMux I__6573 (
            .O(N__29994),
            .I(N__29889));
    Span4Mux_s2_h I__6572 (
            .O(N__29991),
            .I(N__29889));
    LocalMux I__6571 (
            .O(N__29982),
            .I(N__29889));
    LocalMux I__6570 (
            .O(N__29973),
            .I(N__29889));
    LocalMux I__6569 (
            .O(N__29968),
            .I(N__29889));
    InMux I__6568 (
            .O(N__29967),
            .I(N__29866));
    InMux I__6567 (
            .O(N__29966),
            .I(N__29866));
    InMux I__6566 (
            .O(N__29965),
            .I(N__29866));
    InMux I__6565 (
            .O(N__29964),
            .I(N__29866));
    InMux I__6564 (
            .O(N__29963),
            .I(N__29866));
    InMux I__6563 (
            .O(N__29962),
            .I(N__29866));
    LocalMux I__6562 (
            .O(N__29959),
            .I(N__29855));
    LocalMux I__6561 (
            .O(N__29952),
            .I(N__29855));
    LocalMux I__6560 (
            .O(N__29945),
            .I(N__29855));
    LocalMux I__6559 (
            .O(N__29940),
            .I(N__29855));
    LocalMux I__6558 (
            .O(N__29929),
            .I(N__29855));
    InMux I__6557 (
            .O(N__29928),
            .I(N__29848));
    InMux I__6556 (
            .O(N__29927),
            .I(N__29848));
    InMux I__6555 (
            .O(N__29924),
            .I(N__29848));
    LocalMux I__6554 (
            .O(N__29921),
            .I(N__29845));
    Span4Mux_h I__6553 (
            .O(N__29918),
            .I(N__29842));
    Span4Mux_h I__6552 (
            .O(N__29915),
            .I(N__29839));
    InMux I__6551 (
            .O(N__29914),
            .I(N__29832));
    InMux I__6550 (
            .O(N__29913),
            .I(N__29832));
    InMux I__6549 (
            .O(N__29912),
            .I(N__29832));
    InMux I__6548 (
            .O(N__29911),
            .I(N__29823));
    InMux I__6547 (
            .O(N__29910),
            .I(N__29823));
    InMux I__6546 (
            .O(N__29909),
            .I(N__29823));
    InMux I__6545 (
            .O(N__29908),
            .I(N__29823));
    Span4Mux_v I__6544 (
            .O(N__29905),
            .I(N__29816));
    Span4Mux_v I__6543 (
            .O(N__29902),
            .I(N__29816));
    Span4Mux_v I__6542 (
            .O(N__29889),
            .I(N__29816));
    InMux I__6541 (
            .O(N__29888),
            .I(N__29803));
    InMux I__6540 (
            .O(N__29887),
            .I(N__29803));
    InMux I__6539 (
            .O(N__29886),
            .I(N__29803));
    InMux I__6538 (
            .O(N__29885),
            .I(N__29803));
    InMux I__6537 (
            .O(N__29884),
            .I(N__29803));
    InMux I__6536 (
            .O(N__29883),
            .I(N__29803));
    InMux I__6535 (
            .O(N__29882),
            .I(N__29794));
    InMux I__6534 (
            .O(N__29881),
            .I(N__29794));
    InMux I__6533 (
            .O(N__29880),
            .I(N__29794));
    InMux I__6532 (
            .O(N__29879),
            .I(N__29794));
    LocalMux I__6531 (
            .O(N__29866),
            .I(N__29785));
    Span4Mux_s3_v I__6530 (
            .O(N__29855),
            .I(N__29785));
    LocalMux I__6529 (
            .O(N__29848),
            .I(N__29785));
    Span4Mux_h I__6528 (
            .O(N__29845),
            .I(N__29785));
    Odrv4 I__6527 (
            .O(N__29842),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__6526 (
            .O(N__29839),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__6525 (
            .O(N__29832),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__6524 (
            .O(N__29823),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__6523 (
            .O(N__29816),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__6522 (
            .O(N__29803),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__6521 (
            .O(N__29794),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__6520 (
            .O(N__29785),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    CascadeMux I__6519 (
            .O(N__29768),
            .I(N__29764));
    InMux I__6518 (
            .O(N__29767),
            .I(N__29761));
    InMux I__6517 (
            .O(N__29764),
            .I(N__29758));
    LocalMux I__6516 (
            .O(N__29761),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    LocalMux I__6515 (
            .O(N__29758),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    CascadeMux I__6514 (
            .O(N__29753),
            .I(N__29750));
    InMux I__6513 (
            .O(N__29750),
            .I(N__29744));
    InMux I__6512 (
            .O(N__29749),
            .I(N__29744));
    LocalMux I__6511 (
            .O(N__29744),
            .I(N__29741));
    Odrv4 I__6510 (
            .O(N__29741),
            .I(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ));
    InMux I__6509 (
            .O(N__29738),
            .I(N__29734));
    InMux I__6508 (
            .O(N__29737),
            .I(N__29731));
    LocalMux I__6507 (
            .O(N__29734),
            .I(N__29726));
    LocalMux I__6506 (
            .O(N__29731),
            .I(N__29726));
    Odrv12 I__6505 (
            .O(N__29726),
            .I(scaler_3_data_11));
    InMux I__6504 (
            .O(N__29723),
            .I(\scaler_3.un2_source_data_0_cry_6 ));
    CascadeMux I__6503 (
            .O(N__29720),
            .I(N__29717));
    InMux I__6502 (
            .O(N__29717),
            .I(N__29711));
    InMux I__6501 (
            .O(N__29716),
            .I(N__29711));
    LocalMux I__6500 (
            .O(N__29711),
            .I(N__29708));
    Odrv12 I__6499 (
            .O(N__29708),
            .I(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ));
    InMux I__6498 (
            .O(N__29705),
            .I(N__29701));
    InMux I__6497 (
            .O(N__29704),
            .I(N__29698));
    LocalMux I__6496 (
            .O(N__29701),
            .I(N__29695));
    LocalMux I__6495 (
            .O(N__29698),
            .I(N__29692));
    Odrv12 I__6494 (
            .O(N__29695),
            .I(scaler_3_data_12));
    Odrv12 I__6493 (
            .O(N__29692),
            .I(scaler_3_data_12));
    InMux I__6492 (
            .O(N__29687),
            .I(\scaler_3.un2_source_data_0_cry_7 ));
    InMux I__6491 (
            .O(N__29684),
            .I(N__29681));
    LocalMux I__6490 (
            .O(N__29681),
            .I(N__29677));
    InMux I__6489 (
            .O(N__29680),
            .I(N__29674));
    Odrv4 I__6488 (
            .O(N__29677),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    LocalMux I__6487 (
            .O(N__29674),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    CascadeMux I__6486 (
            .O(N__29669),
            .I(N__29666));
    InMux I__6485 (
            .O(N__29666),
            .I(N__29663));
    LocalMux I__6484 (
            .O(N__29663),
            .I(N__29660));
    Odrv4 I__6483 (
            .O(N__29660),
            .I(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ));
    InMux I__6482 (
            .O(N__29657),
            .I(N__29653));
    InMux I__6481 (
            .O(N__29656),
            .I(N__29650));
    LocalMux I__6480 (
            .O(N__29653),
            .I(N__29647));
    LocalMux I__6479 (
            .O(N__29650),
            .I(N__29644));
    Span4Mux_h I__6478 (
            .O(N__29647),
            .I(N__29641));
    Span4Mux_v I__6477 (
            .O(N__29644),
            .I(N__29638));
    Odrv4 I__6476 (
            .O(N__29641),
            .I(scaler_3_data_13));
    Odrv4 I__6475 (
            .O(N__29638),
            .I(scaler_3_data_13));
    InMux I__6474 (
            .O(N__29633),
            .I(bfn_8_23_0_));
    InMux I__6473 (
            .O(N__29630),
            .I(\scaler_3.un2_source_data_0_cry_9 ));
    InMux I__6472 (
            .O(N__29627),
            .I(N__29624));
    LocalMux I__6471 (
            .O(N__29624),
            .I(N__29621));
    Odrv12 I__6470 (
            .O(N__29621),
            .I(scaler_3_data_14));
    InMux I__6469 (
            .O(N__29618),
            .I(N__29614));
    CascadeMux I__6468 (
            .O(N__29617),
            .I(N__29611));
    LocalMux I__6467 (
            .O(N__29614),
            .I(N__29606));
    InMux I__6466 (
            .O(N__29611),
            .I(N__29601));
    InMux I__6465 (
            .O(N__29610),
            .I(N__29601));
    InMux I__6464 (
            .O(N__29609),
            .I(N__29598));
    Span4Mux_v I__6463 (
            .O(N__29606),
            .I(N__29593));
    LocalMux I__6462 (
            .O(N__29601),
            .I(N__29593));
    LocalMux I__6461 (
            .O(N__29598),
            .I(\scaler_3.un2_source_data_0 ));
    Odrv4 I__6460 (
            .O(N__29593),
            .I(\scaler_3.un2_source_data_0 ));
    InMux I__6459 (
            .O(N__29588),
            .I(N__29585));
    LocalMux I__6458 (
            .O(N__29585),
            .I(N__29582));
    Span4Mux_v I__6457 (
            .O(N__29582),
            .I(N__29579));
    Span4Mux_h I__6456 (
            .O(N__29579),
            .I(N__29576));
    Odrv4 I__6455 (
            .O(N__29576),
            .I(scaler_3_data_5));
    CEMux I__6454 (
            .O(N__29573),
            .I(N__29552));
    CEMux I__6453 (
            .O(N__29572),
            .I(N__29552));
    CEMux I__6452 (
            .O(N__29571),
            .I(N__29552));
    CEMux I__6451 (
            .O(N__29570),
            .I(N__29552));
    CEMux I__6450 (
            .O(N__29569),
            .I(N__29552));
    CEMux I__6449 (
            .O(N__29568),
            .I(N__29552));
    CEMux I__6448 (
            .O(N__29567),
            .I(N__29552));
    GlobalMux I__6447 (
            .O(N__29552),
            .I(N__29549));
    gio2CtrlBuf I__6446 (
            .O(N__29549),
            .I(debug_CH3_20A_c_0_g));
    InMux I__6445 (
            .O(N__29546),
            .I(N__29543));
    LocalMux I__6444 (
            .O(N__29543),
            .I(N__29540));
    Span4Mux_v I__6443 (
            .O(N__29540),
            .I(N__29537));
    Odrv4 I__6442 (
            .O(N__29537),
            .I(\ppm_encoder_1.N_305 ));
    CascadeMux I__6441 (
            .O(N__29534),
            .I(N__29530));
    InMux I__6440 (
            .O(N__29533),
            .I(N__29527));
    InMux I__6439 (
            .O(N__29530),
            .I(N__29524));
    LocalMux I__6438 (
            .O(N__29527),
            .I(N__29520));
    LocalMux I__6437 (
            .O(N__29524),
            .I(N__29517));
    InMux I__6436 (
            .O(N__29523),
            .I(N__29514));
    Span4Mux_h I__6435 (
            .O(N__29520),
            .I(N__29509));
    Span4Mux_h I__6434 (
            .O(N__29517),
            .I(N__29509));
    LocalMux I__6433 (
            .O(N__29514),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    Odrv4 I__6432 (
            .O(N__29509),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__6431 (
            .O(N__29504),
            .I(N__29501));
    LocalMux I__6430 (
            .O(N__29501),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__6429 (
            .O(N__29498),
            .I(N__29495));
    LocalMux I__6428 (
            .O(N__29495),
            .I(N__29491));
    InMux I__6427 (
            .O(N__29494),
            .I(N__29486));
    Span4Mux_v I__6426 (
            .O(N__29491),
            .I(N__29477));
    InMux I__6425 (
            .O(N__29490),
            .I(N__29474));
    InMux I__6424 (
            .O(N__29489),
            .I(N__29471));
    LocalMux I__6423 (
            .O(N__29486),
            .I(N__29468));
    InMux I__6422 (
            .O(N__29485),
            .I(N__29463));
    CascadeMux I__6421 (
            .O(N__29484),
            .I(N__29457));
    InMux I__6420 (
            .O(N__29483),
            .I(N__29454));
    InMux I__6419 (
            .O(N__29482),
            .I(N__29449));
    InMux I__6418 (
            .O(N__29481),
            .I(N__29449));
    InMux I__6417 (
            .O(N__29480),
            .I(N__29446));
    Span4Mux_h I__6416 (
            .O(N__29477),
            .I(N__29441));
    LocalMux I__6415 (
            .O(N__29474),
            .I(N__29441));
    LocalMux I__6414 (
            .O(N__29471),
            .I(N__29436));
    Span4Mux_v I__6413 (
            .O(N__29468),
            .I(N__29436));
    InMux I__6412 (
            .O(N__29467),
            .I(N__29431));
    InMux I__6411 (
            .O(N__29466),
            .I(N__29431));
    LocalMux I__6410 (
            .O(N__29463),
            .I(N__29428));
    InMux I__6409 (
            .O(N__29462),
            .I(N__29423));
    InMux I__6408 (
            .O(N__29461),
            .I(N__29420));
    InMux I__6407 (
            .O(N__29460),
            .I(N__29415));
    InMux I__6406 (
            .O(N__29457),
            .I(N__29415));
    LocalMux I__6405 (
            .O(N__29454),
            .I(N__29412));
    LocalMux I__6404 (
            .O(N__29449),
            .I(N__29409));
    LocalMux I__6403 (
            .O(N__29446),
            .I(N__29402));
    Span4Mux_h I__6402 (
            .O(N__29441),
            .I(N__29402));
    Span4Mux_v I__6401 (
            .O(N__29436),
            .I(N__29402));
    LocalMux I__6400 (
            .O(N__29431),
            .I(N__29399));
    Span4Mux_v I__6399 (
            .O(N__29428),
            .I(N__29396));
    InMux I__6398 (
            .O(N__29427),
            .I(N__29393));
    InMux I__6397 (
            .O(N__29426),
            .I(N__29389));
    LocalMux I__6396 (
            .O(N__29423),
            .I(N__29385));
    LocalMux I__6395 (
            .O(N__29420),
            .I(N__29374));
    LocalMux I__6394 (
            .O(N__29415),
            .I(N__29374));
    Span4Mux_h I__6393 (
            .O(N__29412),
            .I(N__29374));
    Span4Mux_v I__6392 (
            .O(N__29409),
            .I(N__29374));
    Span4Mux_v I__6391 (
            .O(N__29402),
            .I(N__29374));
    Span4Mux_v I__6390 (
            .O(N__29399),
            .I(N__29367));
    Span4Mux_v I__6389 (
            .O(N__29396),
            .I(N__29367));
    LocalMux I__6388 (
            .O(N__29393),
            .I(N__29367));
    InMux I__6387 (
            .O(N__29392),
            .I(N__29364));
    LocalMux I__6386 (
            .O(N__29389),
            .I(N__29361));
    InMux I__6385 (
            .O(N__29388),
            .I(N__29358));
    Span12Mux_v I__6384 (
            .O(N__29385),
            .I(N__29355));
    Span4Mux_v I__6383 (
            .O(N__29374),
            .I(N__29352));
    Span4Mux_v I__6382 (
            .O(N__29367),
            .I(N__29349));
    LocalMux I__6381 (
            .O(N__29364),
            .I(N__29344));
    Span12Mux_v I__6380 (
            .O(N__29361),
            .I(N__29344));
    LocalMux I__6379 (
            .O(N__29358),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv12 I__6378 (
            .O(N__29355),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__6377 (
            .O(N__29352),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__6376 (
            .O(N__29349),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv12 I__6375 (
            .O(N__29344),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__6374 (
            .O(N__29333),
            .I(N__29330));
    LocalMux I__6373 (
            .O(N__29330),
            .I(N__29326));
    CascadeMux I__6372 (
            .O(N__29329),
            .I(N__29322));
    Span4Mux_h I__6371 (
            .O(N__29326),
            .I(N__29319));
    InMux I__6370 (
            .O(N__29325),
            .I(N__29316));
    InMux I__6369 (
            .O(N__29322),
            .I(N__29313));
    Span4Mux_h I__6368 (
            .O(N__29319),
            .I(N__29308));
    LocalMux I__6367 (
            .O(N__29316),
            .I(N__29308));
    LocalMux I__6366 (
            .O(N__29313),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__6365 (
            .O(N__29308),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    InMux I__6364 (
            .O(N__29303),
            .I(N__29298));
    InMux I__6363 (
            .O(N__29302),
            .I(N__29295));
    InMux I__6362 (
            .O(N__29301),
            .I(N__29292));
    LocalMux I__6361 (
            .O(N__29298),
            .I(N__29289));
    LocalMux I__6360 (
            .O(N__29295),
            .I(N__29286));
    LocalMux I__6359 (
            .O(N__29292),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    Odrv4 I__6358 (
            .O(N__29289),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    Odrv4 I__6357 (
            .O(N__29286),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    CascadeMux I__6356 (
            .O(N__29279),
            .I(N__29276));
    InMux I__6355 (
            .O(N__29276),
            .I(N__29269));
    InMux I__6354 (
            .O(N__29275),
            .I(N__29263));
    InMux I__6353 (
            .O(N__29274),
            .I(N__29263));
    InMux I__6352 (
            .O(N__29273),
            .I(N__29254));
    InMux I__6351 (
            .O(N__29272),
            .I(N__29254));
    LocalMux I__6350 (
            .O(N__29269),
            .I(N__29249));
    InMux I__6349 (
            .O(N__29268),
            .I(N__29246));
    LocalMux I__6348 (
            .O(N__29263),
            .I(N__29241));
    InMux I__6347 (
            .O(N__29262),
            .I(N__29238));
    InMux I__6346 (
            .O(N__29261),
            .I(N__29230));
    InMux I__6345 (
            .O(N__29260),
            .I(N__29230));
    InMux I__6344 (
            .O(N__29259),
            .I(N__29230));
    LocalMux I__6343 (
            .O(N__29254),
            .I(N__29227));
    InMux I__6342 (
            .O(N__29253),
            .I(N__29224));
    CascadeMux I__6341 (
            .O(N__29252),
            .I(N__29219));
    Span4Mux_s2_v I__6340 (
            .O(N__29249),
            .I(N__29214));
    LocalMux I__6339 (
            .O(N__29246),
            .I(N__29211));
    InMux I__6338 (
            .O(N__29245),
            .I(N__29206));
    InMux I__6337 (
            .O(N__29244),
            .I(N__29206));
    Span4Mux_v I__6336 (
            .O(N__29241),
            .I(N__29203));
    LocalMux I__6335 (
            .O(N__29238),
            .I(N__29200));
    InMux I__6334 (
            .O(N__29237),
            .I(N__29197));
    LocalMux I__6333 (
            .O(N__29230),
            .I(N__29188));
    Span4Mux_s2_v I__6332 (
            .O(N__29227),
            .I(N__29188));
    LocalMux I__6331 (
            .O(N__29224),
            .I(N__29188));
    InMux I__6330 (
            .O(N__29223),
            .I(N__29185));
    CascadeMux I__6329 (
            .O(N__29222),
            .I(N__29182));
    InMux I__6328 (
            .O(N__29219),
            .I(N__29174));
    InMux I__6327 (
            .O(N__29218),
            .I(N__29174));
    InMux I__6326 (
            .O(N__29217),
            .I(N__29174));
    Span4Mux_v I__6325 (
            .O(N__29214),
            .I(N__29169));
    Span4Mux_v I__6324 (
            .O(N__29211),
            .I(N__29169));
    LocalMux I__6323 (
            .O(N__29206),
            .I(N__29166));
    Span4Mux_v I__6322 (
            .O(N__29203),
            .I(N__29161));
    Span4Mux_h I__6321 (
            .O(N__29200),
            .I(N__29161));
    LocalMux I__6320 (
            .O(N__29197),
            .I(N__29158));
    InMux I__6319 (
            .O(N__29196),
            .I(N__29153));
    InMux I__6318 (
            .O(N__29195),
            .I(N__29153));
    Span4Mux_v I__6317 (
            .O(N__29188),
            .I(N__29148));
    LocalMux I__6316 (
            .O(N__29185),
            .I(N__29148));
    InMux I__6315 (
            .O(N__29182),
            .I(N__29143));
    InMux I__6314 (
            .O(N__29181),
            .I(N__29143));
    LocalMux I__6313 (
            .O(N__29174),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6312 (
            .O(N__29169),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv12 I__6311 (
            .O(N__29166),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6310 (
            .O(N__29161),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6309 (
            .O(N__29158),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__6308 (
            .O(N__29153),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6307 (
            .O(N__29148),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__6306 (
            .O(N__29143),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    CascadeMux I__6305 (
            .O(N__29126),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    CascadeMux I__6304 (
            .O(N__29123),
            .I(N__29119));
    InMux I__6303 (
            .O(N__29122),
            .I(N__29116));
    InMux I__6302 (
            .O(N__29119),
            .I(N__29113));
    LocalMux I__6301 (
            .O(N__29116),
            .I(N__29109));
    LocalMux I__6300 (
            .O(N__29113),
            .I(N__29106));
    InMux I__6299 (
            .O(N__29112),
            .I(N__29103));
    Span4Mux_h I__6298 (
            .O(N__29109),
            .I(N__29098));
    Span4Mux_s3_h I__6297 (
            .O(N__29106),
            .I(N__29098));
    LocalMux I__6296 (
            .O(N__29103),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv4 I__6295 (
            .O(N__29098),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__6294 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__6293 (
            .O(N__29090),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__6292 (
            .O(N__29087),
            .I(N__29083));
    InMux I__6291 (
            .O(N__29086),
            .I(N__29080));
    LocalMux I__6290 (
            .O(N__29083),
            .I(N__29077));
    LocalMux I__6289 (
            .O(N__29080),
            .I(N__29074));
    Span4Mux_h I__6288 (
            .O(N__29077),
            .I(N__29071));
    Odrv4 I__6287 (
            .O(N__29074),
            .I(frame_decoder_OFF3data_7));
    Odrv4 I__6286 (
            .O(N__29071),
            .I(frame_decoder_OFF3data_7));
    InMux I__6285 (
            .O(N__29066),
            .I(N__29063));
    LocalMux I__6284 (
            .O(N__29063),
            .I(N__29059));
    InMux I__6283 (
            .O(N__29062),
            .I(N__29056));
    Span4Mux_h I__6282 (
            .O(N__29059),
            .I(N__29053));
    LocalMux I__6281 (
            .O(N__29056),
            .I(N__29050));
    Span4Mux_v I__6280 (
            .O(N__29053),
            .I(N__29047));
    Odrv4 I__6279 (
            .O(N__29050),
            .I(frame_decoder_CH3data_7));
    Odrv4 I__6278 (
            .O(N__29047),
            .I(frame_decoder_CH3data_7));
    InMux I__6277 (
            .O(N__29042),
            .I(N__29039));
    LocalMux I__6276 (
            .O(N__29039),
            .I(\scaler_3.N_893_i_l_ofxZ0 ));
    CascadeMux I__6275 (
            .O(N__29036),
            .I(N__29033));
    InMux I__6274 (
            .O(N__29033),
            .I(N__29030));
    LocalMux I__6273 (
            .O(N__29030),
            .I(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ));
    InMux I__6272 (
            .O(N__29027),
            .I(N__29024));
    LocalMux I__6271 (
            .O(N__29024),
            .I(N__29020));
    InMux I__6270 (
            .O(N__29023),
            .I(N__29017));
    Span4Mux_h I__6269 (
            .O(N__29020),
            .I(N__29014));
    LocalMux I__6268 (
            .O(N__29017),
            .I(N__29011));
    Odrv4 I__6267 (
            .O(N__29014),
            .I(scaler_3_data_6));
    Odrv12 I__6266 (
            .O(N__29011),
            .I(scaler_3_data_6));
    InMux I__6265 (
            .O(N__29006),
            .I(\scaler_3.un2_source_data_0_cry_1 ));
    CascadeMux I__6264 (
            .O(N__29003),
            .I(N__29000));
    InMux I__6263 (
            .O(N__29000),
            .I(N__28994));
    InMux I__6262 (
            .O(N__28999),
            .I(N__28994));
    LocalMux I__6261 (
            .O(N__28994),
            .I(N__28991));
    Odrv4 I__6260 (
            .O(N__28991),
            .I(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ));
    CascadeMux I__6259 (
            .O(N__28988),
            .I(N__28985));
    InMux I__6258 (
            .O(N__28985),
            .I(N__28982));
    LocalMux I__6257 (
            .O(N__28982),
            .I(N__28979));
    Span4Mux_h I__6256 (
            .O(N__28979),
            .I(N__28975));
    InMux I__6255 (
            .O(N__28978),
            .I(N__28972));
    Span4Mux_h I__6254 (
            .O(N__28975),
            .I(N__28969));
    LocalMux I__6253 (
            .O(N__28972),
            .I(N__28966));
    Odrv4 I__6252 (
            .O(N__28969),
            .I(scaler_3_data_7));
    Odrv4 I__6251 (
            .O(N__28966),
            .I(scaler_3_data_7));
    InMux I__6250 (
            .O(N__28961),
            .I(\scaler_3.un2_source_data_0_cry_2 ));
    CascadeMux I__6249 (
            .O(N__28958),
            .I(N__28955));
    InMux I__6248 (
            .O(N__28955),
            .I(N__28949));
    InMux I__6247 (
            .O(N__28954),
            .I(N__28949));
    LocalMux I__6246 (
            .O(N__28949),
            .I(N__28946));
    Odrv4 I__6245 (
            .O(N__28946),
            .I(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ));
    InMux I__6244 (
            .O(N__28943),
            .I(N__28940));
    LocalMux I__6243 (
            .O(N__28940),
            .I(N__28936));
    InMux I__6242 (
            .O(N__28939),
            .I(N__28933));
    Span4Mux_v I__6241 (
            .O(N__28936),
            .I(N__28928));
    LocalMux I__6240 (
            .O(N__28933),
            .I(N__28928));
    Odrv4 I__6239 (
            .O(N__28928),
            .I(scaler_3_data_8));
    InMux I__6238 (
            .O(N__28925),
            .I(\scaler_3.un2_source_data_0_cry_3 ));
    CascadeMux I__6237 (
            .O(N__28922),
            .I(N__28919));
    InMux I__6236 (
            .O(N__28919),
            .I(N__28913));
    InMux I__6235 (
            .O(N__28918),
            .I(N__28913));
    LocalMux I__6234 (
            .O(N__28913),
            .I(N__28910));
    Odrv4 I__6233 (
            .O(N__28910),
            .I(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ));
    InMux I__6232 (
            .O(N__28907),
            .I(N__28904));
    LocalMux I__6231 (
            .O(N__28904),
            .I(N__28900));
    InMux I__6230 (
            .O(N__28903),
            .I(N__28897));
    Span12Mux_s8_h I__6229 (
            .O(N__28900),
            .I(N__28894));
    LocalMux I__6228 (
            .O(N__28897),
            .I(N__28891));
    Odrv12 I__6227 (
            .O(N__28894),
            .I(scaler_3_data_9));
    Odrv4 I__6226 (
            .O(N__28891),
            .I(scaler_3_data_9));
    InMux I__6225 (
            .O(N__28886),
            .I(\scaler_3.un2_source_data_0_cry_4 ));
    CascadeMux I__6224 (
            .O(N__28883),
            .I(N__28880));
    InMux I__6223 (
            .O(N__28880),
            .I(N__28874));
    InMux I__6222 (
            .O(N__28879),
            .I(N__28874));
    LocalMux I__6221 (
            .O(N__28874),
            .I(N__28871));
    Odrv12 I__6220 (
            .O(N__28871),
            .I(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ));
    InMux I__6219 (
            .O(N__28868),
            .I(N__28865));
    LocalMux I__6218 (
            .O(N__28865),
            .I(N__28861));
    InMux I__6217 (
            .O(N__28864),
            .I(N__28858));
    Span4Mux_v I__6216 (
            .O(N__28861),
            .I(N__28853));
    LocalMux I__6215 (
            .O(N__28858),
            .I(N__28853));
    Odrv4 I__6214 (
            .O(N__28853),
            .I(scaler_3_data_10));
    InMux I__6213 (
            .O(N__28850),
            .I(\scaler_3.un2_source_data_0_cry_5 ));
    InMux I__6212 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__6211 (
            .O(N__28844),
            .I(frame_decoder_CH3data_2));
    CascadeMux I__6210 (
            .O(N__28841),
            .I(N__28838));
    InMux I__6209 (
            .O(N__28838),
            .I(N__28835));
    LocalMux I__6208 (
            .O(N__28835),
            .I(N__28832));
    Odrv12 I__6207 (
            .O(N__28832),
            .I(frame_decoder_OFF3data_2));
    InMux I__6206 (
            .O(N__28829),
            .I(\scaler_3.un3_source_data_0_cry_1 ));
    InMux I__6205 (
            .O(N__28826),
            .I(N__28823));
    LocalMux I__6204 (
            .O(N__28823),
            .I(N__28820));
    Odrv4 I__6203 (
            .O(N__28820),
            .I(frame_decoder_OFF3data_3));
    CascadeMux I__6202 (
            .O(N__28817),
            .I(N__28814));
    InMux I__6201 (
            .O(N__28814),
            .I(N__28811));
    LocalMux I__6200 (
            .O(N__28811),
            .I(frame_decoder_CH3data_3));
    InMux I__6199 (
            .O(N__28808),
            .I(\scaler_3.un3_source_data_0_cry_2 ));
    InMux I__6198 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__6197 (
            .O(N__28802),
            .I(N__28799));
    Span4Mux_v I__6196 (
            .O(N__28799),
            .I(N__28796));
    Odrv4 I__6195 (
            .O(N__28796),
            .I(frame_decoder_CH3data_4));
    CascadeMux I__6194 (
            .O(N__28793),
            .I(N__28790));
    InMux I__6193 (
            .O(N__28790),
            .I(N__28787));
    LocalMux I__6192 (
            .O(N__28787),
            .I(N__28784));
    Odrv4 I__6191 (
            .O(N__28784),
            .I(frame_decoder_OFF3data_4));
    InMux I__6190 (
            .O(N__28781),
            .I(\scaler_3.un3_source_data_0_cry_3 ));
    InMux I__6189 (
            .O(N__28778),
            .I(N__28775));
    LocalMux I__6188 (
            .O(N__28775),
            .I(frame_decoder_CH3data_5));
    CascadeMux I__6187 (
            .O(N__28772),
            .I(N__28769));
    InMux I__6186 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__6185 (
            .O(N__28766),
            .I(N__28763));
    Odrv12 I__6184 (
            .O(N__28763),
            .I(frame_decoder_OFF3data_5));
    InMux I__6183 (
            .O(N__28760),
            .I(\scaler_3.un3_source_data_0_cry_4 ));
    InMux I__6182 (
            .O(N__28757),
            .I(N__28754));
    LocalMux I__6181 (
            .O(N__28754),
            .I(frame_decoder_CH3data_6));
    CascadeMux I__6180 (
            .O(N__28751),
            .I(N__28748));
    InMux I__6179 (
            .O(N__28748),
            .I(N__28745));
    LocalMux I__6178 (
            .O(N__28745),
            .I(N__28742));
    Odrv4 I__6177 (
            .O(N__28742),
            .I(frame_decoder_OFF3data_6));
    InMux I__6176 (
            .O(N__28739),
            .I(\scaler_3.un3_source_data_0_cry_5 ));
    InMux I__6175 (
            .O(N__28736),
            .I(N__28733));
    LocalMux I__6174 (
            .O(N__28733),
            .I(N__28730));
    Span4Mux_v I__6173 (
            .O(N__28730),
            .I(N__28727));
    Span4Mux_h I__6172 (
            .O(N__28727),
            .I(N__28724));
    Odrv4 I__6171 (
            .O(N__28724),
            .I(\scaler_3.un3_source_data_0_axb_7 ));
    InMux I__6170 (
            .O(N__28721),
            .I(\scaler_3.un3_source_data_0_cry_6 ));
    InMux I__6169 (
            .O(N__28718),
            .I(N__28714));
    InMux I__6168 (
            .O(N__28717),
            .I(N__28711));
    LocalMux I__6167 (
            .O(N__28714),
            .I(N__28708));
    LocalMux I__6166 (
            .O(N__28711),
            .I(N__28705));
    Span4Mux_h I__6165 (
            .O(N__28708),
            .I(N__28694));
    Span4Mux_v I__6164 (
            .O(N__28705),
            .I(N__28694));
    InMux I__6163 (
            .O(N__28704),
            .I(N__28691));
    CascadeMux I__6162 (
            .O(N__28703),
            .I(N__28687));
    CascadeMux I__6161 (
            .O(N__28702),
            .I(N__28682));
    CascadeMux I__6160 (
            .O(N__28701),
            .I(N__28679));
    CascadeMux I__6159 (
            .O(N__28700),
            .I(N__28675));
    InMux I__6158 (
            .O(N__28699),
            .I(N__28668));
    Span4Mux_v I__6157 (
            .O(N__28694),
            .I(N__28663));
    LocalMux I__6156 (
            .O(N__28691),
            .I(N__28663));
    CascadeMux I__6155 (
            .O(N__28690),
            .I(N__28660));
    InMux I__6154 (
            .O(N__28687),
            .I(N__28654));
    InMux I__6153 (
            .O(N__28686),
            .I(N__28641));
    InMux I__6152 (
            .O(N__28685),
            .I(N__28641));
    InMux I__6151 (
            .O(N__28682),
            .I(N__28641));
    InMux I__6150 (
            .O(N__28679),
            .I(N__28641));
    InMux I__6149 (
            .O(N__28678),
            .I(N__28641));
    InMux I__6148 (
            .O(N__28675),
            .I(N__28641));
    CascadeMux I__6147 (
            .O(N__28674),
            .I(N__28638));
    CascadeMux I__6146 (
            .O(N__28673),
            .I(N__28635));
    CascadeMux I__6145 (
            .O(N__28672),
            .I(N__28632));
    CascadeMux I__6144 (
            .O(N__28671),
            .I(N__28629));
    LocalMux I__6143 (
            .O(N__28668),
            .I(N__28626));
    Span4Mux_h I__6142 (
            .O(N__28663),
            .I(N__28623));
    InMux I__6141 (
            .O(N__28660),
            .I(N__28620));
    InMux I__6140 (
            .O(N__28659),
            .I(N__28617));
    CascadeMux I__6139 (
            .O(N__28658),
            .I(N__28614));
    CascadeMux I__6138 (
            .O(N__28657),
            .I(N__28611));
    LocalMux I__6137 (
            .O(N__28654),
            .I(N__28606));
    LocalMux I__6136 (
            .O(N__28641),
            .I(N__28606));
    InMux I__6135 (
            .O(N__28638),
            .I(N__28603));
    InMux I__6134 (
            .O(N__28635),
            .I(N__28599));
    InMux I__6133 (
            .O(N__28632),
            .I(N__28596));
    InMux I__6132 (
            .O(N__28629),
            .I(N__28593));
    Span4Mux_v I__6131 (
            .O(N__28626),
            .I(N__28584));
    Span4Mux_v I__6130 (
            .O(N__28623),
            .I(N__28584));
    LocalMux I__6129 (
            .O(N__28620),
            .I(N__28584));
    LocalMux I__6128 (
            .O(N__28617),
            .I(N__28584));
    InMux I__6127 (
            .O(N__28614),
            .I(N__28581));
    InMux I__6126 (
            .O(N__28611),
            .I(N__28578));
    Span4Mux_v I__6125 (
            .O(N__28606),
            .I(N__28573));
    LocalMux I__6124 (
            .O(N__28603),
            .I(N__28573));
    CascadeMux I__6123 (
            .O(N__28602),
            .I(N__28570));
    LocalMux I__6122 (
            .O(N__28599),
            .I(N__28562));
    LocalMux I__6121 (
            .O(N__28596),
            .I(N__28562));
    LocalMux I__6120 (
            .O(N__28593),
            .I(N__28559));
    Span4Mux_h I__6119 (
            .O(N__28584),
            .I(N__28556));
    LocalMux I__6118 (
            .O(N__28581),
            .I(N__28553));
    LocalMux I__6117 (
            .O(N__28578),
            .I(N__28548));
    Span4Mux_v I__6116 (
            .O(N__28573),
            .I(N__28548));
    InMux I__6115 (
            .O(N__28570),
            .I(N__28545));
    CascadeMux I__6114 (
            .O(N__28569),
            .I(N__28542));
    CascadeMux I__6113 (
            .O(N__28568),
            .I(N__28539));
    CascadeMux I__6112 (
            .O(N__28567),
            .I(N__28536));
    Span4Mux_v I__6111 (
            .O(N__28562),
            .I(N__28532));
    Span4Mux_v I__6110 (
            .O(N__28559),
            .I(N__28529));
    Span4Mux_v I__6109 (
            .O(N__28556),
            .I(N__28526));
    Span4Mux_h I__6108 (
            .O(N__28553),
            .I(N__28523));
    Span4Mux_h I__6107 (
            .O(N__28548),
            .I(N__28518));
    LocalMux I__6106 (
            .O(N__28545),
            .I(N__28518));
    InMux I__6105 (
            .O(N__28542),
            .I(N__28515));
    InMux I__6104 (
            .O(N__28539),
            .I(N__28510));
    InMux I__6103 (
            .O(N__28536),
            .I(N__28510));
    CascadeMux I__6102 (
            .O(N__28535),
            .I(N__28507));
    Span4Mux_h I__6101 (
            .O(N__28532),
            .I(N__28504));
    Span4Mux_h I__6100 (
            .O(N__28529),
            .I(N__28497));
    Span4Mux_v I__6099 (
            .O(N__28526),
            .I(N__28497));
    Span4Mux_v I__6098 (
            .O(N__28523),
            .I(N__28497));
    Span4Mux_h I__6097 (
            .O(N__28518),
            .I(N__28490));
    LocalMux I__6096 (
            .O(N__28515),
            .I(N__28490));
    LocalMux I__6095 (
            .O(N__28510),
            .I(N__28490));
    InMux I__6094 (
            .O(N__28507),
            .I(N__28487));
    Odrv4 I__6093 (
            .O(N__28504),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6092 (
            .O(N__28497),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6091 (
            .O(N__28490),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6090 (
            .O(N__28487),
            .I(CONSTANT_ONE_NET));
    InMux I__6089 (
            .O(N__28478),
            .I(bfn_8_21_0_));
    InMux I__6088 (
            .O(N__28475),
            .I(\scaler_3.un3_source_data_0_cry_8 ));
    CEMux I__6087 (
            .O(N__28472),
            .I(N__28469));
    LocalMux I__6086 (
            .O(N__28469),
            .I(N__28465));
    CEMux I__6085 (
            .O(N__28468),
            .I(N__28461));
    Span4Mux_h I__6084 (
            .O(N__28465),
            .I(N__28458));
    CEMux I__6083 (
            .O(N__28464),
            .I(N__28455));
    LocalMux I__6082 (
            .O(N__28461),
            .I(N__28452));
    Span4Mux_v I__6081 (
            .O(N__28458),
            .I(N__28447));
    LocalMux I__6080 (
            .O(N__28455),
            .I(N__28447));
    Span4Mux_v I__6079 (
            .O(N__28452),
            .I(N__28444));
    Span4Mux_v I__6078 (
            .O(N__28447),
            .I(N__28441));
    Odrv4 I__6077 (
            .O(N__28444),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    Odrv4 I__6076 (
            .O(N__28441),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__6075 (
            .O(N__28436),
            .I(N__28433));
    LocalMux I__6074 (
            .O(N__28433),
            .I(frame_decoder_CH3data_1));
    CascadeMux I__6073 (
            .O(N__28430),
            .I(N__28427));
    InMux I__6072 (
            .O(N__28427),
            .I(N__28424));
    LocalMux I__6071 (
            .O(N__28424),
            .I(N__28421));
    Odrv4 I__6070 (
            .O(N__28421),
            .I(frame_decoder_OFF3data_1));
    InMux I__6069 (
            .O(N__28418),
            .I(\scaler_3.un3_source_data_0_cry_0 ));
    InMux I__6068 (
            .O(N__28415),
            .I(N__28411));
    InMux I__6067 (
            .O(N__28414),
            .I(N__28408));
    LocalMux I__6066 (
            .O(N__28411),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__6065 (
            .O(N__28408),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__6064 (
            .O(N__28403),
            .I(N__28399));
    InMux I__6063 (
            .O(N__28402),
            .I(N__28396));
    LocalMux I__6062 (
            .O(N__28399),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__6061 (
            .O(N__28396),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__6060 (
            .O(N__28391),
            .I(N__28387));
    InMux I__6059 (
            .O(N__28390),
            .I(N__28384));
    InMux I__6058 (
            .O(N__28387),
            .I(N__28381));
    LocalMux I__6057 (
            .O(N__28384),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__6056 (
            .O(N__28381),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__6055 (
            .O(N__28376),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ));
    InMux I__6054 (
            .O(N__28373),
            .I(N__28369));
    InMux I__6053 (
            .O(N__28372),
            .I(N__28366));
    LocalMux I__6052 (
            .O(N__28369),
            .I(N__28363));
    LocalMux I__6051 (
            .O(N__28366),
            .I(N__28360));
    Odrv4 I__6050 (
            .O(N__28363),
            .I(frame_decoder_OFF4data_7));
    Odrv4 I__6049 (
            .O(N__28360),
            .I(frame_decoder_OFF4data_7));
    InMux I__6048 (
            .O(N__28355),
            .I(N__28351));
    InMux I__6047 (
            .O(N__28354),
            .I(N__28348));
    LocalMux I__6046 (
            .O(N__28351),
            .I(N__28345));
    LocalMux I__6045 (
            .O(N__28348),
            .I(N__28342));
    Span4Mux_h I__6044 (
            .O(N__28345),
            .I(N__28339));
    Odrv4 I__6043 (
            .O(N__28342),
            .I(frame_decoder_CH4data_7));
    Odrv4 I__6042 (
            .O(N__28339),
            .I(frame_decoder_CH4data_7));
    InMux I__6041 (
            .O(N__28334),
            .I(N__28331));
    LocalMux I__6040 (
            .O(N__28331),
            .I(N__28328));
    Span4Mux_v I__6039 (
            .O(N__28328),
            .I(N__28325));
    Odrv4 I__6038 (
            .O(N__28325),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    CascadeMux I__6037 (
            .O(N__28322),
            .I(N__28318));
    InMux I__6036 (
            .O(N__28321),
            .I(N__28315));
    InMux I__6035 (
            .O(N__28318),
            .I(N__28312));
    LocalMux I__6034 (
            .O(N__28315),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__6033 (
            .O(N__28312),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    InMux I__6032 (
            .O(N__28307),
            .I(N__28303));
    InMux I__6031 (
            .O(N__28306),
            .I(N__28300));
    LocalMux I__6030 (
            .O(N__28303),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__6029 (
            .O(N__28300),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__6028 (
            .O(N__28295),
            .I(N__28292));
    InMux I__6027 (
            .O(N__28292),
            .I(N__28288));
    InMux I__6026 (
            .O(N__28291),
            .I(N__28285));
    LocalMux I__6025 (
            .O(N__28288),
            .I(N__28282));
    LocalMux I__6024 (
            .O(N__28285),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    Odrv4 I__6023 (
            .O(N__28282),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    InMux I__6022 (
            .O(N__28277),
            .I(N__28271));
    InMux I__6021 (
            .O(N__28276),
            .I(N__28271));
    LocalMux I__6020 (
            .O(N__28271),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    InMux I__6019 (
            .O(N__28268),
            .I(N__28265));
    LocalMux I__6018 (
            .O(N__28265),
            .I(N__28262));
    Span4Mux_h I__6017 (
            .O(N__28262),
            .I(N__28259));
    Odrv4 I__6016 (
            .O(N__28259),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa ));
    CascadeMux I__6015 (
            .O(N__28256),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ));
    InMux I__6014 (
            .O(N__28253),
            .I(N__28249));
    InMux I__6013 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__6012 (
            .O(N__28249),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    LocalMux I__6011 (
            .O(N__28246),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    InMux I__6010 (
            .O(N__28241),
            .I(N__28231));
    InMux I__6009 (
            .O(N__28240),
            .I(N__28231));
    InMux I__6008 (
            .O(N__28239),
            .I(N__28231));
    InMux I__6007 (
            .O(N__28238),
            .I(N__28228));
    LocalMux I__6006 (
            .O(N__28231),
            .I(N__28225));
    LocalMux I__6005 (
            .O(N__28228),
            .I(N__28220));
    Span4Mux_v I__6004 (
            .O(N__28225),
            .I(N__28220));
    Odrv4 I__6003 (
            .O(N__28220),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    InMux I__6002 (
            .O(N__28217),
            .I(N__28213));
    InMux I__6001 (
            .O(N__28216),
            .I(N__28210));
    LocalMux I__6000 (
            .O(N__28213),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    LocalMux I__5999 (
            .O(N__28210),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__5998 (
            .O(N__28205),
            .I(N__28201));
    InMux I__5997 (
            .O(N__28204),
            .I(N__28198));
    LocalMux I__5996 (
            .O(N__28201),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    LocalMux I__5995 (
            .O(N__28198),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__5994 (
            .O(N__28193),
            .I(N__28190));
    LocalMux I__5993 (
            .O(N__28190),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    CascadeMux I__5992 (
            .O(N__28187),
            .I(N__28184));
    InMux I__5991 (
            .O(N__28184),
            .I(N__28181));
    LocalMux I__5990 (
            .O(N__28181),
            .I(N__28178));
    Span4Mux_v I__5989 (
            .O(N__28178),
            .I(N__28173));
    InMux I__5988 (
            .O(N__28177),
            .I(N__28170));
    InMux I__5987 (
            .O(N__28176),
            .I(N__28166));
    Span4Mux_h I__5986 (
            .O(N__28173),
            .I(N__28161));
    LocalMux I__5985 (
            .O(N__28170),
            .I(N__28161));
    InMux I__5984 (
            .O(N__28169),
            .I(N__28158));
    LocalMux I__5983 (
            .O(N__28166),
            .I(N__28153));
    Sp12to4 I__5982 (
            .O(N__28161),
            .I(N__28153));
    LocalMux I__5981 (
            .O(N__28158),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv12 I__5980 (
            .O(N__28153),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__5979 (
            .O(N__28148),
            .I(N__28144));
    InMux I__5978 (
            .O(N__28147),
            .I(N__28141));
    LocalMux I__5977 (
            .O(N__28144),
            .I(N__28138));
    LocalMux I__5976 (
            .O(N__28141),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    Odrv12 I__5975 (
            .O(N__28138),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    InMux I__5974 (
            .O(N__28133),
            .I(N__28129));
    InMux I__5973 (
            .O(N__28132),
            .I(N__28126));
    LocalMux I__5972 (
            .O(N__28129),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    LocalMux I__5971 (
            .O(N__28126),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    CEMux I__5970 (
            .O(N__28121),
            .I(N__28118));
    LocalMux I__5969 (
            .O(N__28118),
            .I(N__28115));
    Span4Mux_v I__5968 (
            .O(N__28115),
            .I(N__28112));
    Span4Mux_h I__5967 (
            .O(N__28112),
            .I(N__28108));
    CEMux I__5966 (
            .O(N__28111),
            .I(N__28105));
    Odrv4 I__5965 (
            .O(N__28108),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    LocalMux I__5964 (
            .O(N__28105),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    CascadeMux I__5963 (
            .O(N__28100),
            .I(N__28096));
    CascadeMux I__5962 (
            .O(N__28099),
            .I(N__28093));
    InMux I__5961 (
            .O(N__28096),
            .I(N__28087));
    InMux I__5960 (
            .O(N__28093),
            .I(N__28087));
    InMux I__5959 (
            .O(N__28092),
            .I(N__28084));
    LocalMux I__5958 (
            .O(N__28087),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__5957 (
            .O(N__28084),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    InMux I__5956 (
            .O(N__28079),
            .I(N__28073));
    InMux I__5955 (
            .O(N__28078),
            .I(N__28073));
    LocalMux I__5954 (
            .O(N__28073),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ));
    InMux I__5953 (
            .O(N__28070),
            .I(N__28067));
    LocalMux I__5952 (
            .O(N__28067),
            .I(N__28063));
    InMux I__5951 (
            .O(N__28066),
            .I(N__28060));
    Span4Mux_v I__5950 (
            .O(N__28063),
            .I(N__28057));
    LocalMux I__5949 (
            .O(N__28060),
            .I(N__28054));
    Odrv4 I__5948 (
            .O(N__28057),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ));
    Odrv4 I__5947 (
            .O(N__28054),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ));
    CEMux I__5946 (
            .O(N__28049),
            .I(N__28046));
    LocalMux I__5945 (
            .O(N__28046),
            .I(N__28042));
    CEMux I__5944 (
            .O(N__28045),
            .I(N__28038));
    Span4Mux_v I__5943 (
            .O(N__28042),
            .I(N__28035));
    CEMux I__5942 (
            .O(N__28041),
            .I(N__28032));
    LocalMux I__5941 (
            .O(N__28038),
            .I(N__28029));
    Span4Mux_h I__5940 (
            .O(N__28035),
            .I(N__28024));
    LocalMux I__5939 (
            .O(N__28032),
            .I(N__28024));
    Span4Mux_h I__5938 (
            .O(N__28029),
            .I(N__28021));
    Span4Mux_v I__5937 (
            .O(N__28024),
            .I(N__28018));
    Span4Mux_h I__5936 (
            .O(N__28021),
            .I(N__28015));
    Span4Mux_v I__5935 (
            .O(N__28018),
            .I(N__28012));
    Span4Mux_h I__5934 (
            .O(N__28015),
            .I(N__28009));
    Odrv4 I__5933 (
            .O(N__28012),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    Odrv4 I__5932 (
            .O(N__28009),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__5931 (
            .O(N__28004),
            .I(N__28001));
    LocalMux I__5930 (
            .O(N__28001),
            .I(N__27997));
    InMux I__5929 (
            .O(N__28000),
            .I(N__27994));
    Odrv4 I__5928 (
            .O(N__27997),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    LocalMux I__5927 (
            .O(N__27994),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    InMux I__5926 (
            .O(N__27989),
            .I(N__27980));
    InMux I__5925 (
            .O(N__27988),
            .I(N__27980));
    InMux I__5924 (
            .O(N__27987),
            .I(N__27980));
    LocalMux I__5923 (
            .O(N__27980),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    InMux I__5922 (
            .O(N__27977),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__5921 (
            .O(N__27974),
            .I(N__27965));
    SRMux I__5920 (
            .O(N__27973),
            .I(N__27965));
    SRMux I__5919 (
            .O(N__27972),
            .I(N__27965));
    GlobalMux I__5918 (
            .O(N__27965),
            .I(N__27962));
    gio2CtrlBuf I__5917 (
            .O(N__27962),
            .I(\ppm_encoder_1.N_320_g ));
    InMux I__5916 (
            .O(N__27959),
            .I(N__27950));
    InMux I__5915 (
            .O(N__27958),
            .I(N__27950));
    InMux I__5914 (
            .O(N__27957),
            .I(N__27942));
    InMux I__5913 (
            .O(N__27956),
            .I(N__27942));
    InMux I__5912 (
            .O(N__27955),
            .I(N__27938));
    LocalMux I__5911 (
            .O(N__27950),
            .I(N__27935));
    InMux I__5910 (
            .O(N__27949),
            .I(N__27930));
    InMux I__5909 (
            .O(N__27948),
            .I(N__27930));
    InMux I__5908 (
            .O(N__27947),
            .I(N__27927));
    LocalMux I__5907 (
            .O(N__27942),
            .I(N__27919));
    InMux I__5906 (
            .O(N__27941),
            .I(N__27916));
    LocalMux I__5905 (
            .O(N__27938),
            .I(N__27907));
    Span4Mux_v I__5904 (
            .O(N__27935),
            .I(N__27907));
    LocalMux I__5903 (
            .O(N__27930),
            .I(N__27907));
    LocalMux I__5902 (
            .O(N__27927),
            .I(N__27907));
    InMux I__5901 (
            .O(N__27926),
            .I(N__27902));
    InMux I__5900 (
            .O(N__27925),
            .I(N__27902));
    InMux I__5899 (
            .O(N__27924),
            .I(N__27899));
    CascadeMux I__5898 (
            .O(N__27923),
            .I(N__27891));
    InMux I__5897 (
            .O(N__27922),
            .I(N__27888));
    Span4Mux_v I__5896 (
            .O(N__27919),
            .I(N__27885));
    LocalMux I__5895 (
            .O(N__27916),
            .I(N__27882));
    Span4Mux_v I__5894 (
            .O(N__27907),
            .I(N__27877));
    LocalMux I__5893 (
            .O(N__27902),
            .I(N__27877));
    LocalMux I__5892 (
            .O(N__27899),
            .I(N__27874));
    InMux I__5891 (
            .O(N__27898),
            .I(N__27867));
    InMux I__5890 (
            .O(N__27897),
            .I(N__27867));
    InMux I__5889 (
            .O(N__27896),
            .I(N__27867));
    InMux I__5888 (
            .O(N__27895),
            .I(N__27862));
    InMux I__5887 (
            .O(N__27894),
            .I(N__27862));
    InMux I__5886 (
            .O(N__27891),
            .I(N__27859));
    LocalMux I__5885 (
            .O(N__27888),
            .I(N__27856));
    Odrv4 I__5884 (
            .O(N__27885),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5883 (
            .O(N__27882),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5882 (
            .O(N__27877),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5881 (
            .O(N__27874),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5880 (
            .O(N__27867),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5879 (
            .O(N__27862),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5878 (
            .O(N__27859),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5877 (
            .O(N__27856),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    CascadeMux I__5876 (
            .O(N__27839),
            .I(N__27834));
    InMux I__5875 (
            .O(N__27838),
            .I(N__27831));
    InMux I__5874 (
            .O(N__27837),
            .I(N__27828));
    InMux I__5873 (
            .O(N__27834),
            .I(N__27825));
    LocalMux I__5872 (
            .O(N__27831),
            .I(N__27822));
    LocalMux I__5871 (
            .O(N__27828),
            .I(N__27819));
    LocalMux I__5870 (
            .O(N__27825),
            .I(N__27816));
    Span4Mux_h I__5869 (
            .O(N__27822),
            .I(N__27813));
    Span4Mux_h I__5868 (
            .O(N__27819),
            .I(N__27806));
    Span4Mux_s1_v I__5867 (
            .O(N__27816),
            .I(N__27806));
    Span4Mux_v I__5866 (
            .O(N__27813),
            .I(N__27806));
    Odrv4 I__5865 (
            .O(N__27806),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__5864 (
            .O(N__27803),
            .I(N__27800));
    LocalMux I__5863 (
            .O(N__27800),
            .I(N__27796));
    CascadeMux I__5862 (
            .O(N__27799),
            .I(N__27793));
    Span4Mux_v I__5861 (
            .O(N__27796),
            .I(N__27790));
    InMux I__5860 (
            .O(N__27793),
            .I(N__27786));
    Span4Mux_v I__5859 (
            .O(N__27790),
            .I(N__27783));
    InMux I__5858 (
            .O(N__27789),
            .I(N__27780));
    LocalMux I__5857 (
            .O(N__27786),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__5856 (
            .O(N__27783),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    LocalMux I__5855 (
            .O(N__27780),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    InMux I__5854 (
            .O(N__27773),
            .I(N__27770));
    LocalMux I__5853 (
            .O(N__27770),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__5852 (
            .O(N__27767),
            .I(N__27764));
    LocalMux I__5851 (
            .O(N__27764),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    InMux I__5850 (
            .O(N__27761),
            .I(N__27758));
    LocalMux I__5849 (
            .O(N__27758),
            .I(N__27755));
    Odrv12 I__5848 (
            .O(N__27755),
            .I(uart_input_drone_c));
    InMux I__5847 (
            .O(N__27752),
            .I(N__27749));
    LocalMux I__5846 (
            .O(N__27749),
            .I(N__27746));
    Odrv4 I__5845 (
            .O(N__27746),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__5844 (
            .O(N__27743),
            .I(N__27740));
    LocalMux I__5843 (
            .O(N__27740),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__5842 (
            .O(N__27737),
            .I(N__27734));
    LocalMux I__5841 (
            .O(N__27734),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__5840 (
            .O(N__27731),
            .I(N__27727));
    InMux I__5839 (
            .O(N__27730),
            .I(N__27724));
    LocalMux I__5838 (
            .O(N__27727),
            .I(N__27720));
    LocalMux I__5837 (
            .O(N__27724),
            .I(N__27717));
    InMux I__5836 (
            .O(N__27723),
            .I(N__27714));
    Span4Mux_v I__5835 (
            .O(N__27720),
            .I(N__27711));
    Span4Mux_h I__5834 (
            .O(N__27717),
            .I(N__27708));
    LocalMux I__5833 (
            .O(N__27714),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__5832 (
            .O(N__27711),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__5831 (
            .O(N__27708),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__5830 (
            .O(N__27701),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__5829 (
            .O(N__27698),
            .I(N__27695));
    LocalMux I__5828 (
            .O(N__27695),
            .I(N__27690));
    InMux I__5827 (
            .O(N__27694),
            .I(N__27687));
    InMux I__5826 (
            .O(N__27693),
            .I(N__27684));
    Span4Mux_h I__5825 (
            .O(N__27690),
            .I(N__27681));
    LocalMux I__5824 (
            .O(N__27687),
            .I(N__27678));
    LocalMux I__5823 (
            .O(N__27684),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__5822 (
            .O(N__27681),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__5821 (
            .O(N__27678),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__5820 (
            .O(N__27671),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    CascadeMux I__5819 (
            .O(N__27668),
            .I(N__27665));
    InMux I__5818 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__5817 (
            .O(N__27662),
            .I(N__27657));
    InMux I__5816 (
            .O(N__27661),
            .I(N__27654));
    InMux I__5815 (
            .O(N__27660),
            .I(N__27651));
    Span4Mux_h I__5814 (
            .O(N__27657),
            .I(N__27648));
    LocalMux I__5813 (
            .O(N__27654),
            .I(N__27645));
    LocalMux I__5812 (
            .O(N__27651),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__5811 (
            .O(N__27648),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__5810 (
            .O(N__27645),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__5809 (
            .O(N__27638),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__5808 (
            .O(N__27635),
            .I(N__27632));
    LocalMux I__5807 (
            .O(N__27632),
            .I(N__27627));
    InMux I__5806 (
            .O(N__27631),
            .I(N__27624));
    InMux I__5805 (
            .O(N__27630),
            .I(N__27621));
    Span4Mux_h I__5804 (
            .O(N__27627),
            .I(N__27618));
    LocalMux I__5803 (
            .O(N__27624),
            .I(N__27615));
    LocalMux I__5802 (
            .O(N__27621),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__5801 (
            .O(N__27618),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv12 I__5800 (
            .O(N__27615),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__5799 (
            .O(N__27608),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__5798 (
            .O(N__27605),
            .I(N__27602));
    LocalMux I__5797 (
            .O(N__27602),
            .I(N__27597));
    InMux I__5796 (
            .O(N__27601),
            .I(N__27594));
    InMux I__5795 (
            .O(N__27600),
            .I(N__27591));
    Span4Mux_h I__5794 (
            .O(N__27597),
            .I(N__27588));
    LocalMux I__5793 (
            .O(N__27594),
            .I(N__27585));
    LocalMux I__5792 (
            .O(N__27591),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__5791 (
            .O(N__27588),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__5790 (
            .O(N__27585),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__5789 (
            .O(N__27578),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__5788 (
            .O(N__27575),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__5787 (
            .O(N__27572),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__5786 (
            .O(N__27569),
            .I(bfn_7_28_0_));
    InMux I__5785 (
            .O(N__27566),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    CascadeMux I__5784 (
            .O(N__27563),
            .I(N__27559));
    InMux I__5783 (
            .O(N__27562),
            .I(N__27554));
    InMux I__5782 (
            .O(N__27559),
            .I(N__27549));
    InMux I__5781 (
            .O(N__27558),
            .I(N__27549));
    InMux I__5780 (
            .O(N__27557),
            .I(N__27546));
    LocalMux I__5779 (
            .O(N__27554),
            .I(N__27541));
    LocalMux I__5778 (
            .O(N__27549),
            .I(N__27541));
    LocalMux I__5777 (
            .O(N__27546),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__5776 (
            .O(N__27541),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__5775 (
            .O(N__27536),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    CascadeMux I__5774 (
            .O(N__27533),
            .I(N__27528));
    InMux I__5773 (
            .O(N__27532),
            .I(N__27520));
    InMux I__5772 (
            .O(N__27531),
            .I(N__27520));
    InMux I__5771 (
            .O(N__27528),
            .I(N__27520));
    InMux I__5770 (
            .O(N__27527),
            .I(N__27517));
    LocalMux I__5769 (
            .O(N__27520),
            .I(N__27514));
    LocalMux I__5768 (
            .O(N__27517),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    Odrv4 I__5767 (
            .O(N__27514),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__5766 (
            .O(N__27509),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__5765 (
            .O(N__27506),
            .I(N__27496));
    InMux I__5764 (
            .O(N__27505),
            .I(N__27496));
    InMux I__5763 (
            .O(N__27504),
            .I(N__27496));
    InMux I__5762 (
            .O(N__27503),
            .I(N__27493));
    LocalMux I__5761 (
            .O(N__27496),
            .I(N__27490));
    LocalMux I__5760 (
            .O(N__27493),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    Odrv4 I__5759 (
            .O(N__27490),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__5758 (
            .O(N__27485),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__5757 (
            .O(N__27482),
            .I(N__27478));
    InMux I__5756 (
            .O(N__27481),
            .I(N__27474));
    LocalMux I__5755 (
            .O(N__27478),
            .I(N__27471));
    InMux I__5754 (
            .O(N__27477),
            .I(N__27468));
    LocalMux I__5753 (
            .O(N__27474),
            .I(N__27465));
    Span4Mux_v I__5752 (
            .O(N__27471),
            .I(N__27462));
    LocalMux I__5751 (
            .O(N__27468),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__5750 (
            .O(N__27465),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__5749 (
            .O(N__27462),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__5748 (
            .O(N__27455),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__5747 (
            .O(N__27452),
            .I(N__27448));
    InMux I__5746 (
            .O(N__27451),
            .I(N__27444));
    LocalMux I__5745 (
            .O(N__27448),
            .I(N__27441));
    InMux I__5744 (
            .O(N__27447),
            .I(N__27438));
    LocalMux I__5743 (
            .O(N__27444),
            .I(N__27435));
    Span4Mux_v I__5742 (
            .O(N__27441),
            .I(N__27432));
    LocalMux I__5741 (
            .O(N__27438),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    Odrv4 I__5740 (
            .O(N__27435),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    Odrv4 I__5739 (
            .O(N__27432),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__5738 (
            .O(N__27425),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__5737 (
            .O(N__27422),
            .I(N__27418));
    InMux I__5736 (
            .O(N__27421),
            .I(N__27414));
    LocalMux I__5735 (
            .O(N__27418),
            .I(N__27411));
    InMux I__5734 (
            .O(N__27417),
            .I(N__27408));
    LocalMux I__5733 (
            .O(N__27414),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__5732 (
            .O(N__27411),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__5731 (
            .O(N__27408),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__5730 (
            .O(N__27401),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    CascadeMux I__5729 (
            .O(N__27398),
            .I(N__27395));
    InMux I__5728 (
            .O(N__27395),
            .I(N__27391));
    InMux I__5727 (
            .O(N__27394),
            .I(N__27387));
    LocalMux I__5726 (
            .O(N__27391),
            .I(N__27384));
    InMux I__5725 (
            .O(N__27390),
            .I(N__27381));
    LocalMux I__5724 (
            .O(N__27387),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__5723 (
            .O(N__27384),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5722 (
            .O(N__27381),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__5721 (
            .O(N__27374),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__5720 (
            .O(N__27371),
            .I(N__27368));
    LocalMux I__5719 (
            .O(N__27368),
            .I(N__27364));
    InMux I__5718 (
            .O(N__27367),
            .I(N__27361));
    Span4Mux_v I__5717 (
            .O(N__27364),
            .I(N__27357));
    LocalMux I__5716 (
            .O(N__27361),
            .I(N__27354));
    InMux I__5715 (
            .O(N__27360),
            .I(N__27351));
    Span4Mux_h I__5714 (
            .O(N__27357),
            .I(N__27348));
    Span4Mux_h I__5713 (
            .O(N__27354),
            .I(N__27345));
    LocalMux I__5712 (
            .O(N__27351),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__5711 (
            .O(N__27348),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__5710 (
            .O(N__27345),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__5709 (
            .O(N__27338),
            .I(bfn_7_27_0_));
    InMux I__5708 (
            .O(N__27335),
            .I(N__27332));
    LocalMux I__5707 (
            .O(N__27332),
            .I(N__27329));
    Odrv4 I__5706 (
            .O(N__27329),
            .I(scaler_4_data_5));
    CascadeMux I__5705 (
            .O(N__27326),
            .I(N__27323));
    InMux I__5704 (
            .O(N__27323),
            .I(N__27320));
    LocalMux I__5703 (
            .O(N__27320),
            .I(N__27316));
    InMux I__5702 (
            .O(N__27319),
            .I(N__27313));
    Span12Mux_s7_h I__5701 (
            .O(N__27316),
            .I(N__27310));
    LocalMux I__5700 (
            .O(N__27313),
            .I(N__27307));
    Odrv12 I__5699 (
            .O(N__27310),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    Odrv12 I__5698 (
            .O(N__27307),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    CEMux I__5697 (
            .O(N__27302),
            .I(N__27298));
    CEMux I__5696 (
            .O(N__27301),
            .I(N__27295));
    LocalMux I__5695 (
            .O(N__27298),
            .I(N__27290));
    LocalMux I__5694 (
            .O(N__27295),
            .I(N__27287));
    CEMux I__5693 (
            .O(N__27294),
            .I(N__27284));
    CEMux I__5692 (
            .O(N__27293),
            .I(N__27280));
    Span4Mux_v I__5691 (
            .O(N__27290),
            .I(N__27277));
    Span4Mux_v I__5690 (
            .O(N__27287),
            .I(N__27274));
    LocalMux I__5689 (
            .O(N__27284),
            .I(N__27271));
    CEMux I__5688 (
            .O(N__27283),
            .I(N__27268));
    LocalMux I__5687 (
            .O(N__27280),
            .I(N__27264));
    Span4Mux_s2_h I__5686 (
            .O(N__27277),
            .I(N__27261));
    Span4Mux_h I__5685 (
            .O(N__27274),
            .I(N__27256));
    Span4Mux_h I__5684 (
            .O(N__27271),
            .I(N__27256));
    LocalMux I__5683 (
            .O(N__27268),
            .I(N__27253));
    CEMux I__5682 (
            .O(N__27267),
            .I(N__27250));
    Odrv12 I__5681 (
            .O(N__27264),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__5680 (
            .O(N__27261),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__5679 (
            .O(N__27256),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv12 I__5678 (
            .O(N__27253),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    LocalMux I__5677 (
            .O(N__27250),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    CascadeMux I__5676 (
            .O(N__27239),
            .I(N__27236));
    InMux I__5675 (
            .O(N__27236),
            .I(N__27233));
    LocalMux I__5674 (
            .O(N__27233),
            .I(N__27230));
    Span4Mux_h I__5673 (
            .O(N__27230),
            .I(N__27227));
    Odrv4 I__5672 (
            .O(N__27227),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__5671 (
            .O(N__27224),
            .I(N__27221));
    LocalMux I__5670 (
            .O(N__27221),
            .I(N__27218));
    Span4Mux_h I__5669 (
            .O(N__27218),
            .I(N__27215));
    Odrv4 I__5668 (
            .O(N__27215),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__5667 (
            .O(N__27212),
            .I(N__27209));
    LocalMux I__5666 (
            .O(N__27209),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__5665 (
            .O(N__27206),
            .I(N__27203));
    LocalMux I__5664 (
            .O(N__27203),
            .I(N__27200));
    Span4Mux_v I__5663 (
            .O(N__27200),
            .I(N__27197));
    Span4Mux_h I__5662 (
            .O(N__27197),
            .I(N__27194));
    Odrv4 I__5661 (
            .O(N__27194),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__5660 (
            .O(N__27191),
            .I(N__27188));
    LocalMux I__5659 (
            .O(N__27188),
            .I(N__27185));
    Span4Mux_h I__5658 (
            .O(N__27185),
            .I(N__27182));
    Odrv4 I__5657 (
            .O(N__27182),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    CascadeMux I__5656 (
            .O(N__27179),
            .I(N__27176));
    InMux I__5655 (
            .O(N__27176),
            .I(N__27173));
    LocalMux I__5654 (
            .O(N__27173),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__5653 (
            .O(N__27170),
            .I(N__27167));
    LocalMux I__5652 (
            .O(N__27167),
            .I(N__27164));
    Span4Mux_h I__5651 (
            .O(N__27164),
            .I(N__27161));
    Odrv4 I__5650 (
            .O(N__27161),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__5649 (
            .O(N__27158),
            .I(N__27155));
    LocalMux I__5648 (
            .O(N__27155),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    InMux I__5647 (
            .O(N__27152),
            .I(N__27149));
    LocalMux I__5646 (
            .O(N__27149),
            .I(N__27146));
    Span4Mux_h I__5645 (
            .O(N__27146),
            .I(N__27143));
    Odrv4 I__5644 (
            .O(N__27143),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__5643 (
            .O(N__27140),
            .I(N__27137));
    LocalMux I__5642 (
            .O(N__27137),
            .I(N__27134));
    Odrv4 I__5641 (
            .O(N__27134),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    CascadeMux I__5640 (
            .O(N__27131),
            .I(N__27128));
    InMux I__5639 (
            .O(N__27128),
            .I(N__27125));
    LocalMux I__5638 (
            .O(N__27125),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    CascadeMux I__5637 (
            .O(N__27122),
            .I(N__27114));
    InMux I__5636 (
            .O(N__27121),
            .I(N__27098));
    InMux I__5635 (
            .O(N__27120),
            .I(N__27098));
    InMux I__5634 (
            .O(N__27119),
            .I(N__27098));
    InMux I__5633 (
            .O(N__27118),
            .I(N__27093));
    InMux I__5632 (
            .O(N__27117),
            .I(N__27093));
    InMux I__5631 (
            .O(N__27114),
            .I(N__27080));
    InMux I__5630 (
            .O(N__27113),
            .I(N__27080));
    InMux I__5629 (
            .O(N__27112),
            .I(N__27080));
    InMux I__5628 (
            .O(N__27111),
            .I(N__27080));
    InMux I__5627 (
            .O(N__27110),
            .I(N__27080));
    InMux I__5626 (
            .O(N__27109),
            .I(N__27080));
    InMux I__5625 (
            .O(N__27108),
            .I(N__27071));
    InMux I__5624 (
            .O(N__27107),
            .I(N__27071));
    InMux I__5623 (
            .O(N__27106),
            .I(N__27071));
    InMux I__5622 (
            .O(N__27105),
            .I(N__27071));
    LocalMux I__5621 (
            .O(N__27098),
            .I(N__27068));
    LocalMux I__5620 (
            .O(N__27093),
            .I(N__27065));
    LocalMux I__5619 (
            .O(N__27080),
            .I(N__27060));
    LocalMux I__5618 (
            .O(N__27071),
            .I(N__27060));
    Span4Mux_h I__5617 (
            .O(N__27068),
            .I(N__27053));
    Span4Mux_h I__5616 (
            .O(N__27065),
            .I(N__27053));
    Span4Mux_v I__5615 (
            .O(N__27060),
            .I(N__27053));
    Span4Mux_v I__5614 (
            .O(N__27053),
            .I(N__27050));
    Span4Mux_v I__5613 (
            .O(N__27050),
            .I(N__27047));
    Odrv4 I__5612 (
            .O(N__27047),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__5611 (
            .O(N__27044),
            .I(N__27041));
    LocalMux I__5610 (
            .O(N__27041),
            .I(N__27038));
    Span4Mux_v I__5609 (
            .O(N__27038),
            .I(N__27035));
    Span4Mux_h I__5608 (
            .O(N__27035),
            .I(N__27032));
    Span4Mux_v I__5607 (
            .O(N__27032),
            .I(N__27029));
    Odrv4 I__5606 (
            .O(N__27029),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    InMux I__5605 (
            .O(N__27026),
            .I(N__27023));
    LocalMux I__5604 (
            .O(N__27023),
            .I(N__27020));
    Span4Mux_v I__5603 (
            .O(N__27020),
            .I(N__27017));
    Odrv4 I__5602 (
            .O(N__27017),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    CEMux I__5601 (
            .O(N__27014),
            .I(N__27010));
    CEMux I__5600 (
            .O(N__27013),
            .I(N__27007));
    LocalMux I__5599 (
            .O(N__27010),
            .I(N__27004));
    LocalMux I__5598 (
            .O(N__27007),
            .I(N__27001));
    Span4Mux_h I__5597 (
            .O(N__27004),
            .I(N__26998));
    Span4Mux_v I__5596 (
            .O(N__27001),
            .I(N__26994));
    IoSpan4Mux I__5595 (
            .O(N__26998),
            .I(N__26991));
    CEMux I__5594 (
            .O(N__26997),
            .I(N__26988));
    Span4Mux_h I__5593 (
            .O(N__26994),
            .I(N__26983));
    Span4Mux_s2_v I__5592 (
            .O(N__26991),
            .I(N__26983));
    LocalMux I__5591 (
            .O(N__26988),
            .I(N__26980));
    Span4Mux_h I__5590 (
            .O(N__26983),
            .I(N__26975));
    Span4Mux_v I__5589 (
            .O(N__26980),
            .I(N__26975));
    Span4Mux_h I__5588 (
            .O(N__26975),
            .I(N__26972));
    Odrv4 I__5587 (
            .O(N__26972),
            .I(\ppm_encoder_1.N_1014_0 ));
    CascadeMux I__5586 (
            .O(N__26969),
            .I(N__26965));
    InMux I__5585 (
            .O(N__26968),
            .I(N__26962));
    InMux I__5584 (
            .O(N__26965),
            .I(N__26959));
    LocalMux I__5583 (
            .O(N__26962),
            .I(N__26954));
    LocalMux I__5582 (
            .O(N__26959),
            .I(N__26954));
    Span4Mux_v I__5581 (
            .O(N__26954),
            .I(N__26951));
    Span4Mux_h I__5580 (
            .O(N__26951),
            .I(N__26948));
    Odrv4 I__5579 (
            .O(N__26948),
            .I(\ppm_encoder_1.N_1014_i ));
    InMux I__5578 (
            .O(N__26945),
            .I(N__26938));
    InMux I__5577 (
            .O(N__26944),
            .I(N__26938));
    InMux I__5576 (
            .O(N__26943),
            .I(N__26935));
    LocalMux I__5575 (
            .O(N__26938),
            .I(N__26932));
    LocalMux I__5574 (
            .O(N__26935),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__5573 (
            .O(N__26932),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    CascadeMux I__5572 (
            .O(N__26927),
            .I(N__26924));
    InMux I__5571 (
            .O(N__26924),
            .I(N__26918));
    InMux I__5570 (
            .O(N__26923),
            .I(N__26918));
    LocalMux I__5569 (
            .O(N__26918),
            .I(N__26915));
    Odrv4 I__5568 (
            .O(N__26915),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__5567 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__5566 (
            .O(N__26909),
            .I(N__26905));
    InMux I__5565 (
            .O(N__26908),
            .I(N__26902));
    Span4Mux_v I__5564 (
            .O(N__26905),
            .I(N__26899));
    LocalMux I__5563 (
            .O(N__26902),
            .I(N__26896));
    Span4Mux_v I__5562 (
            .O(N__26899),
            .I(N__26893));
    Odrv4 I__5561 (
            .O(N__26896),
            .I(scaler_4_data_11));
    Odrv4 I__5560 (
            .O(N__26893),
            .I(scaler_4_data_11));
    InMux I__5559 (
            .O(N__26888),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__5558 (
            .O(N__26885),
            .I(N__26882));
    InMux I__5557 (
            .O(N__26882),
            .I(N__26876));
    InMux I__5556 (
            .O(N__26881),
            .I(N__26876));
    LocalMux I__5555 (
            .O(N__26876),
            .I(N__26873));
    Odrv12 I__5554 (
            .O(N__26873),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__5553 (
            .O(N__26870),
            .I(N__26866));
    InMux I__5552 (
            .O(N__26869),
            .I(N__26863));
    LocalMux I__5551 (
            .O(N__26866),
            .I(N__26860));
    LocalMux I__5550 (
            .O(N__26863),
            .I(N__26857));
    Span4Mux_v I__5549 (
            .O(N__26860),
            .I(N__26854));
    Span4Mux_h I__5548 (
            .O(N__26857),
            .I(N__26849));
    Span4Mux_v I__5547 (
            .O(N__26854),
            .I(N__26849));
    Odrv4 I__5546 (
            .O(N__26849),
            .I(scaler_4_data_12));
    InMux I__5545 (
            .O(N__26846),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__5544 (
            .O(N__26843),
            .I(N__26840));
    LocalMux I__5543 (
            .O(N__26840),
            .I(N__26836));
    InMux I__5542 (
            .O(N__26839),
            .I(N__26833));
    Odrv4 I__5541 (
            .O(N__26836),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__5540 (
            .O(N__26833),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    CascadeMux I__5539 (
            .O(N__26828),
            .I(N__26825));
    InMux I__5538 (
            .O(N__26825),
            .I(N__26822));
    LocalMux I__5537 (
            .O(N__26822),
            .I(N__26819));
    Odrv4 I__5536 (
            .O(N__26819),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    CascadeMux I__5535 (
            .O(N__26816),
            .I(N__26812));
    InMux I__5534 (
            .O(N__26815),
            .I(N__26809));
    InMux I__5533 (
            .O(N__26812),
            .I(N__26806));
    LocalMux I__5532 (
            .O(N__26809),
            .I(N__26803));
    LocalMux I__5531 (
            .O(N__26806),
            .I(N__26798));
    Span4Mux_v I__5530 (
            .O(N__26803),
            .I(N__26798));
    Span4Mux_v I__5529 (
            .O(N__26798),
            .I(N__26795));
    Odrv4 I__5528 (
            .O(N__26795),
            .I(scaler_4_data_13));
    InMux I__5527 (
            .O(N__26792),
            .I(bfn_7_22_0_));
    InMux I__5526 (
            .O(N__26789),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__5525 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__5524 (
            .O(N__26783),
            .I(N__26780));
    Span4Mux_v I__5523 (
            .O(N__26780),
            .I(N__26777));
    Span4Mux_v I__5522 (
            .O(N__26777),
            .I(N__26774));
    Odrv4 I__5521 (
            .O(N__26774),
            .I(scaler_4_data_14));
    InMux I__5520 (
            .O(N__26771),
            .I(N__26767));
    CascadeMux I__5519 (
            .O(N__26770),
            .I(N__26764));
    LocalMux I__5518 (
            .O(N__26767),
            .I(N__26759));
    InMux I__5517 (
            .O(N__26764),
            .I(N__26754));
    InMux I__5516 (
            .O(N__26763),
            .I(N__26754));
    InMux I__5515 (
            .O(N__26762),
            .I(N__26751));
    Span4Mux_v I__5514 (
            .O(N__26759),
            .I(N__26746));
    LocalMux I__5513 (
            .O(N__26754),
            .I(N__26746));
    LocalMux I__5512 (
            .O(N__26751),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__5511 (
            .O(N__26746),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__5510 (
            .O(N__26741),
            .I(N__26735));
    InMux I__5509 (
            .O(N__26740),
            .I(N__26732));
    InMux I__5508 (
            .O(N__26739),
            .I(N__26729));
    CascadeMux I__5507 (
            .O(N__26738),
            .I(N__26726));
    LocalMux I__5506 (
            .O(N__26735),
            .I(N__26719));
    LocalMux I__5505 (
            .O(N__26732),
            .I(N__26719));
    LocalMux I__5504 (
            .O(N__26729),
            .I(N__26719));
    InMux I__5503 (
            .O(N__26726),
            .I(N__26716));
    Span4Mux_v I__5502 (
            .O(N__26719),
            .I(N__26711));
    LocalMux I__5501 (
            .O(N__26716),
            .I(N__26711));
    Odrv4 I__5500 (
            .O(N__26711),
            .I(frame_decoder_OFF4data_0));
    InMux I__5499 (
            .O(N__26708),
            .I(N__26703));
    InMux I__5498 (
            .O(N__26707),
            .I(N__26700));
    InMux I__5497 (
            .O(N__26706),
            .I(N__26697));
    LocalMux I__5496 (
            .O(N__26703),
            .I(N__26691));
    LocalMux I__5495 (
            .O(N__26700),
            .I(N__26691));
    LocalMux I__5494 (
            .O(N__26697),
            .I(N__26688));
    InMux I__5493 (
            .O(N__26696),
            .I(N__26685));
    Odrv12 I__5492 (
            .O(N__26691),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__5491 (
            .O(N__26688),
            .I(frame_decoder_CH4data_0));
    LocalMux I__5490 (
            .O(N__26685),
            .I(frame_decoder_CH4data_0));
    InMux I__5489 (
            .O(N__26678),
            .I(N__26674));
    InMux I__5488 (
            .O(N__26677),
            .I(N__26671));
    LocalMux I__5487 (
            .O(N__26674),
            .I(N__26666));
    LocalMux I__5486 (
            .O(N__26671),
            .I(N__26666));
    Odrv12 I__5485 (
            .O(N__26666),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    CascadeMux I__5484 (
            .O(N__26663),
            .I(N__26659));
    InMux I__5483 (
            .O(N__26662),
            .I(N__26656));
    InMux I__5482 (
            .O(N__26659),
            .I(N__26653));
    LocalMux I__5481 (
            .O(N__26656),
            .I(scaler_4_data_4));
    LocalMux I__5480 (
            .O(N__26653),
            .I(scaler_4_data_4));
    InMux I__5479 (
            .O(N__26648),
            .I(N__26645));
    LocalMux I__5478 (
            .O(N__26645),
            .I(N__26642));
    Span4Mux_s3_v I__5477 (
            .O(N__26642),
            .I(N__26638));
    InMux I__5476 (
            .O(N__26641),
            .I(N__26635));
    Span4Mux_h I__5475 (
            .O(N__26638),
            .I(N__26632));
    LocalMux I__5474 (
            .O(N__26635),
            .I(N__26629));
    Odrv4 I__5473 (
            .O(N__26632),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv12 I__5472 (
            .O(N__26629),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    InMux I__5471 (
            .O(N__26624),
            .I(N__26621));
    LocalMux I__5470 (
            .O(N__26621),
            .I(\scaler_4.N_905_i_l_ofxZ0 ));
    CascadeMux I__5469 (
            .O(N__26618),
            .I(N__26615));
    InMux I__5468 (
            .O(N__26615),
            .I(N__26612));
    LocalMux I__5467 (
            .O(N__26612),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ));
    InMux I__5466 (
            .O(N__26609),
            .I(N__26605));
    InMux I__5465 (
            .O(N__26608),
            .I(N__26602));
    LocalMux I__5464 (
            .O(N__26605),
            .I(N__26599));
    LocalMux I__5463 (
            .O(N__26602),
            .I(N__26596));
    Span4Mux_v I__5462 (
            .O(N__26599),
            .I(N__26593));
    Span4Mux_v I__5461 (
            .O(N__26596),
            .I(N__26588));
    Span4Mux_v I__5460 (
            .O(N__26593),
            .I(N__26588));
    Odrv4 I__5459 (
            .O(N__26588),
            .I(scaler_4_data_6));
    InMux I__5458 (
            .O(N__26585),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__5457 (
            .O(N__26582),
            .I(N__26579));
    InMux I__5456 (
            .O(N__26579),
            .I(N__26573));
    InMux I__5455 (
            .O(N__26578),
            .I(N__26573));
    LocalMux I__5454 (
            .O(N__26573),
            .I(N__26570));
    Odrv4 I__5453 (
            .O(N__26570),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__5452 (
            .O(N__26567),
            .I(N__26563));
    InMux I__5451 (
            .O(N__26566),
            .I(N__26560));
    LocalMux I__5450 (
            .O(N__26563),
            .I(N__26557));
    LocalMux I__5449 (
            .O(N__26560),
            .I(N__26554));
    Span4Mux_v I__5448 (
            .O(N__26557),
            .I(N__26551));
    Span4Mux_h I__5447 (
            .O(N__26554),
            .I(N__26546));
    Span4Mux_v I__5446 (
            .O(N__26551),
            .I(N__26546));
    Odrv4 I__5445 (
            .O(N__26546),
            .I(scaler_4_data_7));
    InMux I__5444 (
            .O(N__26543),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    CascadeMux I__5443 (
            .O(N__26540),
            .I(N__26537));
    InMux I__5442 (
            .O(N__26537),
            .I(N__26531));
    InMux I__5441 (
            .O(N__26536),
            .I(N__26531));
    LocalMux I__5440 (
            .O(N__26531),
            .I(N__26528));
    Odrv4 I__5439 (
            .O(N__26528),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    CascadeMux I__5438 (
            .O(N__26525),
            .I(N__26521));
    InMux I__5437 (
            .O(N__26524),
            .I(N__26518));
    InMux I__5436 (
            .O(N__26521),
            .I(N__26515));
    LocalMux I__5435 (
            .O(N__26518),
            .I(N__26512));
    LocalMux I__5434 (
            .O(N__26515),
            .I(N__26509));
    Span4Mux_v I__5433 (
            .O(N__26512),
            .I(N__26506));
    Span4Mux_v I__5432 (
            .O(N__26509),
            .I(N__26503));
    Span4Mux_v I__5431 (
            .O(N__26506),
            .I(N__26500));
    Odrv4 I__5430 (
            .O(N__26503),
            .I(scaler_4_data_8));
    Odrv4 I__5429 (
            .O(N__26500),
            .I(scaler_4_data_8));
    InMux I__5428 (
            .O(N__26495),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    CascadeMux I__5427 (
            .O(N__26492),
            .I(N__26489));
    InMux I__5426 (
            .O(N__26489),
            .I(N__26483));
    InMux I__5425 (
            .O(N__26488),
            .I(N__26483));
    LocalMux I__5424 (
            .O(N__26483),
            .I(N__26480));
    Odrv4 I__5423 (
            .O(N__26480),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__5422 (
            .O(N__26477),
            .I(N__26474));
    LocalMux I__5421 (
            .O(N__26474),
            .I(N__26470));
    InMux I__5420 (
            .O(N__26473),
            .I(N__26467));
    Span4Mux_v I__5419 (
            .O(N__26470),
            .I(N__26464));
    LocalMux I__5418 (
            .O(N__26467),
            .I(N__26461));
    Span4Mux_h I__5417 (
            .O(N__26464),
            .I(N__26456));
    Span4Mux_v I__5416 (
            .O(N__26461),
            .I(N__26456));
    Span4Mux_v I__5415 (
            .O(N__26456),
            .I(N__26453));
    Odrv4 I__5414 (
            .O(N__26453),
            .I(scaler_4_data_9));
    InMux I__5413 (
            .O(N__26450),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__5412 (
            .O(N__26447),
            .I(N__26444));
    InMux I__5411 (
            .O(N__26444),
            .I(N__26438));
    InMux I__5410 (
            .O(N__26443),
            .I(N__26438));
    LocalMux I__5409 (
            .O(N__26438),
            .I(N__26435));
    Odrv12 I__5408 (
            .O(N__26435),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__5407 (
            .O(N__26432),
            .I(N__26428));
    InMux I__5406 (
            .O(N__26431),
            .I(N__26425));
    LocalMux I__5405 (
            .O(N__26428),
            .I(N__26422));
    LocalMux I__5404 (
            .O(N__26425),
            .I(N__26417));
    Span4Mux_v I__5403 (
            .O(N__26422),
            .I(N__26417));
    Span4Mux_v I__5402 (
            .O(N__26417),
            .I(N__26414));
    Odrv4 I__5401 (
            .O(N__26414),
            .I(scaler_4_data_10));
    InMux I__5400 (
            .O(N__26411),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    InMux I__5399 (
            .O(N__26408),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__5398 (
            .O(N__26405),
            .I(N__26402));
    LocalMux I__5397 (
            .O(N__26402),
            .I(N__26399));
    Odrv4 I__5396 (
            .O(N__26399),
            .I(frame_decoder_OFF4data_2));
    CascadeMux I__5395 (
            .O(N__26396),
            .I(N__26393));
    InMux I__5394 (
            .O(N__26393),
            .I(N__26390));
    LocalMux I__5393 (
            .O(N__26390),
            .I(frame_decoder_CH4data_2));
    InMux I__5392 (
            .O(N__26387),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__5391 (
            .O(N__26384),
            .I(N__26381));
    LocalMux I__5390 (
            .O(N__26381),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__5389 (
            .O(N__26378),
            .I(N__26375));
    InMux I__5388 (
            .O(N__26375),
            .I(N__26372));
    LocalMux I__5387 (
            .O(N__26372),
            .I(N__26369));
    Odrv12 I__5386 (
            .O(N__26369),
            .I(frame_decoder_OFF4data_3));
    InMux I__5385 (
            .O(N__26366),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__5384 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__5383 (
            .O(N__26360),
            .I(N__26357));
    Odrv12 I__5382 (
            .O(N__26357),
            .I(frame_decoder_OFF4data_4));
    CascadeMux I__5381 (
            .O(N__26354),
            .I(N__26351));
    InMux I__5380 (
            .O(N__26351),
            .I(N__26348));
    LocalMux I__5379 (
            .O(N__26348),
            .I(frame_decoder_CH4data_4));
    InMux I__5378 (
            .O(N__26345),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__5377 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5376 (
            .O(N__26339),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__5375 (
            .O(N__26336),
            .I(N__26333));
    InMux I__5374 (
            .O(N__26333),
            .I(N__26330));
    LocalMux I__5373 (
            .O(N__26330),
            .I(N__26327));
    Odrv12 I__5372 (
            .O(N__26327),
            .I(frame_decoder_OFF4data_5));
    InMux I__5371 (
            .O(N__26324),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__5370 (
            .O(N__26321),
            .I(N__26318));
    LocalMux I__5369 (
            .O(N__26318),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__5368 (
            .O(N__26315),
            .I(N__26312));
    InMux I__5367 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__5366 (
            .O(N__26309),
            .I(N__26306));
    Odrv12 I__5365 (
            .O(N__26306),
            .I(frame_decoder_OFF4data_6));
    InMux I__5364 (
            .O(N__26303),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__5363 (
            .O(N__26300),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__5362 (
            .O(N__26297),
            .I(bfn_7_20_0_));
    InMux I__5361 (
            .O(N__26294),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CEMux I__5360 (
            .O(N__26291),
            .I(N__26288));
    LocalMux I__5359 (
            .O(N__26288),
            .I(N__26285));
    Span4Mux_v I__5358 (
            .O(N__26285),
            .I(N__26282));
    Odrv4 I__5357 (
            .O(N__26282),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__5356 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__5355 (
            .O(N__26276),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__5354 (
            .O(N__26273),
            .I(N__26270));
    InMux I__5353 (
            .O(N__26270),
            .I(N__26267));
    LocalMux I__5352 (
            .O(N__26267),
            .I(N__26264));
    Odrv4 I__5351 (
            .O(N__26264),
            .I(frame_decoder_OFF4data_1));
    InMux I__5350 (
            .O(N__26261),
            .I(N__26256));
    InMux I__5349 (
            .O(N__26260),
            .I(N__26253));
    InMux I__5348 (
            .O(N__26259),
            .I(N__26250));
    LocalMux I__5347 (
            .O(N__26256),
            .I(N__26245));
    LocalMux I__5346 (
            .O(N__26253),
            .I(N__26245));
    LocalMux I__5345 (
            .O(N__26250),
            .I(N__26242));
    Span4Mux_h I__5344 (
            .O(N__26245),
            .I(N__26239));
    Span4Mux_h I__5343 (
            .O(N__26242),
            .I(N__26236));
    Odrv4 I__5342 (
            .O(N__26239),
            .I(uart_drone_data_5));
    Odrv4 I__5341 (
            .O(N__26236),
            .I(uart_drone_data_5));
    InMux I__5340 (
            .O(N__26231),
            .I(N__26226));
    CascadeMux I__5339 (
            .O(N__26230),
            .I(N__26222));
    InMux I__5338 (
            .O(N__26229),
            .I(N__26219));
    LocalMux I__5337 (
            .O(N__26226),
            .I(N__26216));
    InMux I__5336 (
            .O(N__26225),
            .I(N__26213));
    InMux I__5335 (
            .O(N__26222),
            .I(N__26210));
    LocalMux I__5334 (
            .O(N__26219),
            .I(N__26207));
    Span4Mux_h I__5333 (
            .O(N__26216),
            .I(N__26204));
    LocalMux I__5332 (
            .O(N__26213),
            .I(N__26199));
    LocalMux I__5331 (
            .O(N__26210),
            .I(N__26199));
    Span12Mux_s7_h I__5330 (
            .O(N__26207),
            .I(N__26196));
    Span4Mux_v I__5329 (
            .O(N__26204),
            .I(N__26193));
    Span4Mux_h I__5328 (
            .O(N__26199),
            .I(N__26190));
    Odrv12 I__5327 (
            .O(N__26196),
            .I(uart_drone_data_6));
    Odrv4 I__5326 (
            .O(N__26193),
            .I(uart_drone_data_6));
    Odrv4 I__5325 (
            .O(N__26190),
            .I(uart_drone_data_6));
    InMux I__5324 (
            .O(N__26183),
            .I(N__26180));
    LocalMux I__5323 (
            .O(N__26180),
            .I(N__26175));
    InMux I__5322 (
            .O(N__26179),
            .I(N__26172));
    InMux I__5321 (
            .O(N__26178),
            .I(N__26169));
    Span4Mux_h I__5320 (
            .O(N__26175),
            .I(N__26166));
    LocalMux I__5319 (
            .O(N__26172),
            .I(N__26163));
    LocalMux I__5318 (
            .O(N__26169),
            .I(N__26160));
    Span4Mux_v I__5317 (
            .O(N__26166),
            .I(N__26157));
    Span12Mux_s7_h I__5316 (
            .O(N__26163),
            .I(N__26154));
    Span4Mux_h I__5315 (
            .O(N__26160),
            .I(N__26151));
    Odrv4 I__5314 (
            .O(N__26157),
            .I(uart_drone_data_7));
    Odrv12 I__5313 (
            .O(N__26154),
            .I(uart_drone_data_7));
    Odrv4 I__5312 (
            .O(N__26151),
            .I(uart_drone_data_7));
    CascadeMux I__5311 (
            .O(N__26144),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    IoInMux I__5310 (
            .O(N__26141),
            .I(N__26138));
    LocalMux I__5309 (
            .O(N__26138),
            .I(N__26135));
    Span12Mux_s4_v I__5308 (
            .O(N__26135),
            .I(N__26132));
    Span12Mux_v I__5307 (
            .O(N__26132),
            .I(N__26129));
    Odrv12 I__5306 (
            .O(N__26129),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__5305 (
            .O(N__26126),
            .I(N__26122));
    InMux I__5304 (
            .O(N__26125),
            .I(N__26119));
    LocalMux I__5303 (
            .O(N__26122),
            .I(N__26115));
    LocalMux I__5302 (
            .O(N__26119),
            .I(N__26112));
    InMux I__5301 (
            .O(N__26118),
            .I(N__26109));
    Span4Mux_v I__5300 (
            .O(N__26115),
            .I(N__26106));
    Span4Mux_v I__5299 (
            .O(N__26112),
            .I(N__26101));
    LocalMux I__5298 (
            .O(N__26109),
            .I(N__26101));
    Span4Mux_h I__5297 (
            .O(N__26106),
            .I(N__26098));
    Span4Mux_h I__5296 (
            .O(N__26101),
            .I(N__26095));
    Odrv4 I__5295 (
            .O(N__26098),
            .I(uart_drone_data_0));
    Odrv4 I__5294 (
            .O(N__26095),
            .I(uart_drone_data_0));
    InMux I__5293 (
            .O(N__26090),
            .I(N__26086));
    InMux I__5292 (
            .O(N__26089),
            .I(N__26083));
    LocalMux I__5291 (
            .O(N__26086),
            .I(N__26076));
    LocalMux I__5290 (
            .O(N__26083),
            .I(N__26076));
    InMux I__5289 (
            .O(N__26082),
            .I(N__26073));
    InMux I__5288 (
            .O(N__26081),
            .I(N__26070));
    Span4Mux_v I__5287 (
            .O(N__26076),
            .I(N__26067));
    LocalMux I__5286 (
            .O(N__26073),
            .I(N__26062));
    LocalMux I__5285 (
            .O(N__26070),
            .I(N__26062));
    Span4Mux_h I__5284 (
            .O(N__26067),
            .I(N__26059));
    Span4Mux_h I__5283 (
            .O(N__26062),
            .I(N__26056));
    Odrv4 I__5282 (
            .O(N__26059),
            .I(uart_drone_data_1));
    Odrv4 I__5281 (
            .O(N__26056),
            .I(uart_drone_data_1));
    InMux I__5280 (
            .O(N__26051),
            .I(N__26047));
    CascadeMux I__5279 (
            .O(N__26050),
            .I(N__26043));
    LocalMux I__5278 (
            .O(N__26047),
            .I(N__26040));
    InMux I__5277 (
            .O(N__26046),
            .I(N__26037));
    InMux I__5276 (
            .O(N__26043),
            .I(N__26034));
    Span4Mux_h I__5275 (
            .O(N__26040),
            .I(N__26031));
    LocalMux I__5274 (
            .O(N__26037),
            .I(N__26028));
    LocalMux I__5273 (
            .O(N__26034),
            .I(N__26025));
    Span4Mux_v I__5272 (
            .O(N__26031),
            .I(N__26022));
    Span4Mux_h I__5271 (
            .O(N__26028),
            .I(N__26019));
    Span4Mux_h I__5270 (
            .O(N__26025),
            .I(N__26016));
    Odrv4 I__5269 (
            .O(N__26022),
            .I(uart_drone_data_2));
    Odrv4 I__5268 (
            .O(N__26019),
            .I(uart_drone_data_2));
    Odrv4 I__5267 (
            .O(N__26016),
            .I(uart_drone_data_2));
    InMux I__5266 (
            .O(N__26009),
            .I(N__26006));
    LocalMux I__5265 (
            .O(N__26006),
            .I(N__26000));
    InMux I__5264 (
            .O(N__26005),
            .I(N__25997));
    InMux I__5263 (
            .O(N__26004),
            .I(N__25994));
    InMux I__5262 (
            .O(N__26003),
            .I(N__25991));
    Span4Mux_v I__5261 (
            .O(N__26000),
            .I(N__25988));
    LocalMux I__5260 (
            .O(N__25997),
            .I(N__25985));
    LocalMux I__5259 (
            .O(N__25994),
            .I(N__25980));
    LocalMux I__5258 (
            .O(N__25991),
            .I(N__25980));
    Span4Mux_h I__5257 (
            .O(N__25988),
            .I(N__25977));
    Span4Mux_h I__5256 (
            .O(N__25985),
            .I(N__25974));
    Span4Mux_h I__5255 (
            .O(N__25980),
            .I(N__25971));
    Odrv4 I__5254 (
            .O(N__25977),
            .I(uart_drone_data_3));
    Odrv4 I__5253 (
            .O(N__25974),
            .I(uart_drone_data_3));
    Odrv4 I__5252 (
            .O(N__25971),
            .I(uart_drone_data_3));
    InMux I__5251 (
            .O(N__25964),
            .I(N__25959));
    InMux I__5250 (
            .O(N__25963),
            .I(N__25955));
    InMux I__5249 (
            .O(N__25962),
            .I(N__25952));
    LocalMux I__5248 (
            .O(N__25959),
            .I(N__25949));
    InMux I__5247 (
            .O(N__25958),
            .I(N__25946));
    LocalMux I__5246 (
            .O(N__25955),
            .I(N__25943));
    LocalMux I__5245 (
            .O(N__25952),
            .I(N__25940));
    Span4Mux_v I__5244 (
            .O(N__25949),
            .I(N__25937));
    LocalMux I__5243 (
            .O(N__25946),
            .I(N__25934));
    Span4Mux_h I__5242 (
            .O(N__25943),
            .I(N__25931));
    Span4Mux_v I__5241 (
            .O(N__25940),
            .I(N__25928));
    Span4Mux_v I__5240 (
            .O(N__25937),
            .I(N__25923));
    Span4Mux_v I__5239 (
            .O(N__25934),
            .I(N__25923));
    Odrv4 I__5238 (
            .O(N__25931),
            .I(uart_drone_data_4));
    Odrv4 I__5237 (
            .O(N__25928),
            .I(uart_drone_data_4));
    Odrv4 I__5236 (
            .O(N__25923),
            .I(uart_drone_data_4));
    InMux I__5235 (
            .O(N__25916),
            .I(N__25913));
    LocalMux I__5234 (
            .O(N__25913),
            .I(N__25907));
    InMux I__5233 (
            .O(N__25912),
            .I(N__25902));
    InMux I__5232 (
            .O(N__25911),
            .I(N__25902));
    CascadeMux I__5231 (
            .O(N__25910),
            .I(N__25898));
    Span4Mux_v I__5230 (
            .O(N__25907),
            .I(N__25892));
    LocalMux I__5229 (
            .O(N__25902),
            .I(N__25892));
    InMux I__5228 (
            .O(N__25901),
            .I(N__25885));
    InMux I__5227 (
            .O(N__25898),
            .I(N__25885));
    InMux I__5226 (
            .O(N__25897),
            .I(N__25885));
    Span4Mux_v I__5225 (
            .O(N__25892),
            .I(N__25882));
    LocalMux I__5224 (
            .O(N__25885),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__5223 (
            .O(N__25882),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    CEMux I__5222 (
            .O(N__25877),
            .I(N__25874));
    LocalMux I__5221 (
            .O(N__25874),
            .I(N__25871));
    Span4Mux_h I__5220 (
            .O(N__25871),
            .I(N__25868));
    Odrv4 I__5219 (
            .O(N__25868),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    CascadeMux I__5218 (
            .O(N__25865),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ));
    InMux I__5217 (
            .O(N__25862),
            .I(N__25859));
    LocalMux I__5216 (
            .O(N__25859),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_3_2 ));
    CascadeMux I__5215 (
            .O(N__25856),
            .I(N__25853));
    InMux I__5214 (
            .O(N__25853),
            .I(N__25847));
    InMux I__5213 (
            .O(N__25852),
            .I(N__25847));
    LocalMux I__5212 (
            .O(N__25847),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    InMux I__5211 (
            .O(N__25844),
            .I(N__25832));
    InMux I__5210 (
            .O(N__25843),
            .I(N__25832));
    InMux I__5209 (
            .O(N__25842),
            .I(N__25832));
    InMux I__5208 (
            .O(N__25841),
            .I(N__25832));
    LocalMux I__5207 (
            .O(N__25832),
            .I(N__25829));
    Span4Mux_v I__5206 (
            .O(N__25829),
            .I(N__25825));
    InMux I__5205 (
            .O(N__25828),
            .I(N__25822));
    Odrv4 I__5204 (
            .O(N__25825),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    LocalMux I__5203 (
            .O(N__25822),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    CascadeMux I__5202 (
            .O(N__25817),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ));
    InMux I__5201 (
            .O(N__25814),
            .I(N__25810));
    InMux I__5200 (
            .O(N__25813),
            .I(N__25807));
    LocalMux I__5199 (
            .O(N__25810),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    LocalMux I__5198 (
            .O(N__25807),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    InMux I__5197 (
            .O(N__25802),
            .I(N__25799));
    LocalMux I__5196 (
            .O(N__25799),
            .I(N__25796));
    Span4Mux_v I__5195 (
            .O(N__25796),
            .I(N__25793));
    Odrv4 I__5194 (
            .O(N__25793),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    InMux I__5193 (
            .O(N__25790),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__5192 (
            .O(N__25787),
            .I(bfn_5_30_0_));
    CascadeMux I__5191 (
            .O(N__25784),
            .I(N__25781));
    InMux I__5190 (
            .O(N__25781),
            .I(N__25778));
    LocalMux I__5189 (
            .O(N__25778),
            .I(N__25774));
    InMux I__5188 (
            .O(N__25777),
            .I(N__25771));
    Span4Mux_v I__5187 (
            .O(N__25774),
            .I(N__25768));
    LocalMux I__5186 (
            .O(N__25771),
            .I(N__25765));
    Span4Mux_h I__5185 (
            .O(N__25768),
            .I(N__25762));
    Odrv12 I__5184 (
            .O(N__25765),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv4 I__5183 (
            .O(N__25762),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    CEMux I__5182 (
            .O(N__25757),
            .I(N__25751));
    CEMux I__5181 (
            .O(N__25756),
            .I(N__25748));
    CEMux I__5180 (
            .O(N__25755),
            .I(N__25745));
    CEMux I__5179 (
            .O(N__25754),
            .I(N__25742));
    LocalMux I__5178 (
            .O(N__25751),
            .I(N__25739));
    LocalMux I__5177 (
            .O(N__25748),
            .I(N__25736));
    LocalMux I__5176 (
            .O(N__25745),
            .I(N__25733));
    LocalMux I__5175 (
            .O(N__25742),
            .I(N__25730));
    Span4Mux_v I__5174 (
            .O(N__25739),
            .I(N__25725));
    Span4Mux_s3_h I__5173 (
            .O(N__25736),
            .I(N__25725));
    Span4Mux_h I__5172 (
            .O(N__25733),
            .I(N__25722));
    Span4Mux_h I__5171 (
            .O(N__25730),
            .I(N__25719));
    Span4Mux_h I__5170 (
            .O(N__25725),
            .I(N__25716));
    Odrv4 I__5169 (
            .O(N__25722),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__5168 (
            .O(N__25719),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__5167 (
            .O(N__25716),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    CEMux I__5166 (
            .O(N__25709),
            .I(N__25706));
    LocalMux I__5165 (
            .O(N__25706),
            .I(N__25700));
    CEMux I__5164 (
            .O(N__25705),
            .I(N__25697));
    CEMux I__5163 (
            .O(N__25704),
            .I(N__25694));
    CEMux I__5162 (
            .O(N__25703),
            .I(N__25691));
    Span4Mux_h I__5161 (
            .O(N__25700),
            .I(N__25686));
    LocalMux I__5160 (
            .O(N__25697),
            .I(N__25686));
    LocalMux I__5159 (
            .O(N__25694),
            .I(N__25683));
    LocalMux I__5158 (
            .O(N__25691),
            .I(N__25680));
    Span4Mux_v I__5157 (
            .O(N__25686),
            .I(N__25677));
    Span4Mux_h I__5156 (
            .O(N__25683),
            .I(N__25674));
    Span4Mux_h I__5155 (
            .O(N__25680),
            .I(N__25671));
    Span4Mux_h I__5154 (
            .O(N__25677),
            .I(N__25668));
    Span4Mux_h I__5153 (
            .O(N__25674),
            .I(N__25665));
    Span4Mux_v I__5152 (
            .O(N__25671),
            .I(N__25660));
    Span4Mux_h I__5151 (
            .O(N__25668),
            .I(N__25660));
    Odrv4 I__5150 (
            .O(N__25665),
            .I(\dron_frame_decoder_1.N_390_0 ));
    Odrv4 I__5149 (
            .O(N__25660),
            .I(\dron_frame_decoder_1.N_390_0 ));
    CascadeMux I__5148 (
            .O(N__25655),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ));
    CEMux I__5147 (
            .O(N__25652),
            .I(N__25649));
    LocalMux I__5146 (
            .O(N__25649),
            .I(N__25645));
    CEMux I__5145 (
            .O(N__25648),
            .I(N__25642));
    Span4Mux_v I__5144 (
            .O(N__25645),
            .I(N__25637));
    LocalMux I__5143 (
            .O(N__25642),
            .I(N__25637));
    Span4Mux_v I__5142 (
            .O(N__25637),
            .I(N__25633));
    CEMux I__5141 (
            .O(N__25636),
            .I(N__25630));
    Span4Mux_h I__5140 (
            .O(N__25633),
            .I(N__25627));
    LocalMux I__5139 (
            .O(N__25630),
            .I(N__25624));
    Odrv4 I__5138 (
            .O(N__25627),
            .I(\dron_frame_decoder_1.N_382_0 ));
    Odrv12 I__5137 (
            .O(N__25624),
            .I(\dron_frame_decoder_1.N_382_0 ));
    CascadeMux I__5136 (
            .O(N__25619),
            .I(N__25614));
    CascadeMux I__5135 (
            .O(N__25618),
            .I(N__25611));
    InMux I__5134 (
            .O(N__25617),
            .I(N__25604));
    InMux I__5133 (
            .O(N__25614),
            .I(N__25604));
    InMux I__5132 (
            .O(N__25611),
            .I(N__25604));
    LocalMux I__5131 (
            .O(N__25604),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    InMux I__5130 (
            .O(N__25601),
            .I(N__25598));
    LocalMux I__5129 (
            .O(N__25598),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__5128 (
            .O(N__25595),
            .I(N__25592));
    LocalMux I__5127 (
            .O(N__25592),
            .I(N__25589));
    Span4Mux_v I__5126 (
            .O(N__25589),
            .I(N__25586));
    Span4Mux_v I__5125 (
            .O(N__25586),
            .I(N__25583));
    Odrv4 I__5124 (
            .O(N__25583),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__5123 (
            .O(N__25580),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__5122 (
            .O(N__25577),
            .I(N__25574));
    LocalMux I__5121 (
            .O(N__25574),
            .I(N__25571));
    Span4Mux_v I__5120 (
            .O(N__25571),
            .I(N__25568));
    Span4Mux_v I__5119 (
            .O(N__25568),
            .I(N__25565));
    Odrv4 I__5118 (
            .O(N__25565),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__5117 (
            .O(N__25562),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    CascadeMux I__5116 (
            .O(N__25559),
            .I(N__25556));
    InMux I__5115 (
            .O(N__25556),
            .I(N__25553));
    LocalMux I__5114 (
            .O(N__25553),
            .I(N__25550));
    Span4Mux_h I__5113 (
            .O(N__25550),
            .I(N__25547));
    Odrv4 I__5112 (
            .O(N__25547),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__5111 (
            .O(N__25544),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__5110 (
            .O(N__25541),
            .I(N__25538));
    LocalMux I__5109 (
            .O(N__25538),
            .I(N__25535));
    Odrv12 I__5108 (
            .O(N__25535),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__5107 (
            .O(N__25532),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    CascadeMux I__5106 (
            .O(N__25529),
            .I(N__25526));
    InMux I__5105 (
            .O(N__25526),
            .I(N__25523));
    LocalMux I__5104 (
            .O(N__25523),
            .I(N__25520));
    Span4Mux_v I__5103 (
            .O(N__25520),
            .I(N__25517));
    Span4Mux_v I__5102 (
            .O(N__25517),
            .I(N__25514));
    Odrv4 I__5101 (
            .O(N__25514),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__5100 (
            .O(N__25511),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__5099 (
            .O(N__25508),
            .I(N__25505));
    LocalMux I__5098 (
            .O(N__25505),
            .I(N__25502));
    Span12Mux_v I__5097 (
            .O(N__25502),
            .I(N__25499));
    Odrv12 I__5096 (
            .O(N__25499),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__5095 (
            .O(N__25496),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__5094 (
            .O(N__25493),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    CascadeMux I__5093 (
            .O(N__25490),
            .I(N__25486));
    InMux I__5092 (
            .O(N__25489),
            .I(N__25482));
    InMux I__5091 (
            .O(N__25486),
            .I(N__25477));
    InMux I__5090 (
            .O(N__25485),
            .I(N__25477));
    LocalMux I__5089 (
            .O(N__25482),
            .I(N__25474));
    LocalMux I__5088 (
            .O(N__25477),
            .I(N__25471));
    Span4Mux_h I__5087 (
            .O(N__25474),
            .I(N__25468));
    Span4Mux_v I__5086 (
            .O(N__25471),
            .I(N__25465));
    Odrv4 I__5085 (
            .O(N__25468),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__5084 (
            .O(N__25465),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    CascadeMux I__5083 (
            .O(N__25460),
            .I(N__25457));
    InMux I__5082 (
            .O(N__25457),
            .I(N__25452));
    InMux I__5081 (
            .O(N__25456),
            .I(N__25449));
    CascadeMux I__5080 (
            .O(N__25455),
            .I(N__25446));
    LocalMux I__5079 (
            .O(N__25452),
            .I(N__25443));
    LocalMux I__5078 (
            .O(N__25449),
            .I(N__25440));
    InMux I__5077 (
            .O(N__25446),
            .I(N__25437));
    Span4Mux_v I__5076 (
            .O(N__25443),
            .I(N__25434));
    Span4Mux_h I__5075 (
            .O(N__25440),
            .I(N__25431));
    LocalMux I__5074 (
            .O(N__25437),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__5073 (
            .O(N__25434),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__5072 (
            .O(N__25431),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__5071 (
            .O(N__25424),
            .I(N__25421));
    LocalMux I__5070 (
            .O(N__25421),
            .I(N__25418));
    Span4Mux_h I__5069 (
            .O(N__25418),
            .I(N__25415));
    Odrv4 I__5068 (
            .O(N__25415),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__5067 (
            .O(N__25412),
            .I(N__25408));
    InMux I__5066 (
            .O(N__25411),
            .I(N__25405));
    LocalMux I__5065 (
            .O(N__25408),
            .I(N__25402));
    LocalMux I__5064 (
            .O(N__25405),
            .I(\ppm_encoder_1.N_238 ));
    Odrv4 I__5063 (
            .O(N__25402),
            .I(\ppm_encoder_1.N_238 ));
    InMux I__5062 (
            .O(N__25397),
            .I(N__25392));
    InMux I__5061 (
            .O(N__25396),
            .I(N__25389));
    InMux I__5060 (
            .O(N__25395),
            .I(N__25386));
    LocalMux I__5059 (
            .O(N__25392),
            .I(N__25383));
    LocalMux I__5058 (
            .O(N__25389),
            .I(N__25377));
    LocalMux I__5057 (
            .O(N__25386),
            .I(N__25377));
    Span4Mux_s2_v I__5056 (
            .O(N__25383),
            .I(N__25374));
    InMux I__5055 (
            .O(N__25382),
            .I(N__25371));
    Odrv4 I__5054 (
            .O(N__25377),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__5053 (
            .O(N__25374),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__5052 (
            .O(N__25371),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    CascadeMux I__5051 (
            .O(N__25364),
            .I(N__25359));
    CascadeMux I__5050 (
            .O(N__25363),
            .I(N__25354));
    InMux I__5049 (
            .O(N__25362),
            .I(N__25351));
    InMux I__5048 (
            .O(N__25359),
            .I(N__25348));
    InMux I__5047 (
            .O(N__25358),
            .I(N__25341));
    InMux I__5046 (
            .O(N__25357),
            .I(N__25341));
    InMux I__5045 (
            .O(N__25354),
            .I(N__25341));
    LocalMux I__5044 (
            .O(N__25351),
            .I(N__25338));
    LocalMux I__5043 (
            .O(N__25348),
            .I(N__25335));
    LocalMux I__5042 (
            .O(N__25341),
            .I(N__25330));
    Span4Mux_v I__5041 (
            .O(N__25338),
            .I(N__25325));
    Span4Mux_v I__5040 (
            .O(N__25335),
            .I(N__25325));
    InMux I__5039 (
            .O(N__25334),
            .I(N__25320));
    InMux I__5038 (
            .O(N__25333),
            .I(N__25320));
    Odrv4 I__5037 (
            .O(N__25330),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__5036 (
            .O(N__25325),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__5035 (
            .O(N__25320),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    IoInMux I__5034 (
            .O(N__25313),
            .I(N__25310));
    LocalMux I__5033 (
            .O(N__25310),
            .I(N__25307));
    Span4Mux_s2_v I__5032 (
            .O(N__25307),
            .I(N__25304));
    Sp12to4 I__5031 (
            .O(N__25304),
            .I(N__25301));
    Odrv12 I__5030 (
            .O(N__25301),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__5029 (
            .O(N__25298),
            .I(N__25293));
    InMux I__5028 (
            .O(N__25297),
            .I(N__25289));
    InMux I__5027 (
            .O(N__25296),
            .I(N__25286));
    LocalMux I__5026 (
            .O(N__25293),
            .I(N__25283));
    InMux I__5025 (
            .O(N__25292),
            .I(N__25280));
    LocalMux I__5024 (
            .O(N__25289),
            .I(N__25274));
    LocalMux I__5023 (
            .O(N__25286),
            .I(N__25274));
    Span4Mux_s3_v I__5022 (
            .O(N__25283),
            .I(N__25271));
    LocalMux I__5021 (
            .O(N__25280),
            .I(N__25268));
    InMux I__5020 (
            .O(N__25279),
            .I(N__25263));
    Span4Mux_s3_v I__5019 (
            .O(N__25274),
            .I(N__25260));
    Span4Mux_h I__5018 (
            .O(N__25271),
            .I(N__25255));
    Span4Mux_s3_v I__5017 (
            .O(N__25268),
            .I(N__25255));
    InMux I__5016 (
            .O(N__25267),
            .I(N__25252));
    InMux I__5015 (
            .O(N__25266),
            .I(N__25249));
    LocalMux I__5014 (
            .O(N__25263),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__5013 (
            .O(N__25260),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__5012 (
            .O(N__25255),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__5011 (
            .O(N__25252),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__5010 (
            .O(N__25249),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__5009 (
            .O(N__25238),
            .I(N__25233));
    InMux I__5008 (
            .O(N__25237),
            .I(N__25230));
    CascadeMux I__5007 (
            .O(N__25236),
            .I(N__25226));
    LocalMux I__5006 (
            .O(N__25233),
            .I(N__25222));
    LocalMux I__5005 (
            .O(N__25230),
            .I(N__25219));
    InMux I__5004 (
            .O(N__25229),
            .I(N__25216));
    InMux I__5003 (
            .O(N__25226),
            .I(N__25210));
    InMux I__5002 (
            .O(N__25225),
            .I(N__25210));
    Span4Mux_s2_v I__5001 (
            .O(N__25222),
            .I(N__25207));
    Span4Mux_s2_v I__5000 (
            .O(N__25219),
            .I(N__25202));
    LocalMux I__4999 (
            .O(N__25216),
            .I(N__25202));
    InMux I__4998 (
            .O(N__25215),
            .I(N__25199));
    LocalMux I__4997 (
            .O(N__25210),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__4996 (
            .O(N__25207),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__4995 (
            .O(N__25202),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4994 (
            .O(N__25199),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    InMux I__4993 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__4992 (
            .O(N__25187),
            .I(N__25181));
    InMux I__4991 (
            .O(N__25186),
            .I(N__25176));
    InMux I__4990 (
            .O(N__25185),
            .I(N__25176));
    InMux I__4989 (
            .O(N__25184),
            .I(N__25173));
    Span4Mux_h I__4988 (
            .O(N__25181),
            .I(N__25168));
    LocalMux I__4987 (
            .O(N__25176),
            .I(N__25168));
    LocalMux I__4986 (
            .O(N__25173),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__4985 (
            .O(N__25168),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__4984 (
            .O(N__25163),
            .I(N__25160));
    LocalMux I__4983 (
            .O(N__25160),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    InMux I__4982 (
            .O(N__25157),
            .I(N__25154));
    LocalMux I__4981 (
            .O(N__25154),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    CascadeMux I__4980 (
            .O(N__25151),
            .I(N__25148));
    InMux I__4979 (
            .O(N__25148),
            .I(N__25145));
    LocalMux I__4978 (
            .O(N__25145),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__4977 (
            .O(N__25142),
            .I(N__25136));
    InMux I__4976 (
            .O(N__25141),
            .I(N__25136));
    LocalMux I__4975 (
            .O(N__25136),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    InMux I__4974 (
            .O(N__25133),
            .I(N__25130));
    LocalMux I__4973 (
            .O(N__25130),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    CascadeMux I__4972 (
            .O(N__25127),
            .I(N__25124));
    InMux I__4971 (
            .O(N__25124),
            .I(N__25121));
    LocalMux I__4970 (
            .O(N__25121),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__4969 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__4968 (
            .O(N__25115),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__4967 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__4966 (
            .O(N__25109),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__4965 (
            .O(N__25106),
            .I(N__25103));
    LocalMux I__4964 (
            .O(N__25103),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__4963 (
            .O(N__25100),
            .I(N__25097));
    LocalMux I__4962 (
            .O(N__25097),
            .I(N__25094));
    Odrv4 I__4961 (
            .O(N__25094),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    CascadeMux I__4960 (
            .O(N__25091),
            .I(N__25088));
    InMux I__4959 (
            .O(N__25088),
            .I(N__25085));
    LocalMux I__4958 (
            .O(N__25085),
            .I(N__25082));
    Span4Mux_v I__4957 (
            .O(N__25082),
            .I(N__25079));
    Odrv4 I__4956 (
            .O(N__25079),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__4955 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__4954 (
            .O(N__25073),
            .I(N__25070));
    Span4Mux_v I__4953 (
            .O(N__25070),
            .I(N__25066));
    InMux I__4952 (
            .O(N__25069),
            .I(N__25063));
    Odrv4 I__4951 (
            .O(N__25066),
            .I(throttle_command_1));
    LocalMux I__4950 (
            .O(N__25063),
            .I(throttle_command_1));
    InMux I__4949 (
            .O(N__25058),
            .I(N__25055));
    LocalMux I__4948 (
            .O(N__25055),
            .I(N__25050));
    InMux I__4947 (
            .O(N__25054),
            .I(N__25047));
    InMux I__4946 (
            .O(N__25053),
            .I(N__25044));
    Span4Mux_h I__4945 (
            .O(N__25050),
            .I(N__25041));
    LocalMux I__4944 (
            .O(N__25047),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    LocalMux I__4943 (
            .O(N__25044),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__4942 (
            .O(N__25041),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    InMux I__4941 (
            .O(N__25034),
            .I(N__25031));
    LocalMux I__4940 (
            .O(N__25031),
            .I(N__25028));
    Span4Mux_h I__4939 (
            .O(N__25028),
            .I(N__25025));
    Odrv4 I__4938 (
            .O(N__25025),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__4937 (
            .O(N__25022),
            .I(N__25018));
    InMux I__4936 (
            .O(N__25021),
            .I(N__25015));
    LocalMux I__4935 (
            .O(N__25018),
            .I(N__25012));
    LocalMux I__4934 (
            .O(N__25015),
            .I(N__25009));
    Span4Mux_v I__4933 (
            .O(N__25012),
            .I(N__25004));
    Span4Mux_v I__4932 (
            .O(N__25009),
            .I(N__25004));
    Odrv4 I__4931 (
            .O(N__25004),
            .I(throttle_command_3));
    CascadeMux I__4930 (
            .O(N__25001),
            .I(N__24993));
    CascadeMux I__4929 (
            .O(N__25000),
            .I(N__24988));
    CascadeMux I__4928 (
            .O(N__24999),
            .I(N__24977));
    CascadeMux I__4927 (
            .O(N__24998),
            .I(N__24974));
    CascadeMux I__4926 (
            .O(N__24997),
            .I(N__24967));
    InMux I__4925 (
            .O(N__24996),
            .I(N__24964));
    InMux I__4924 (
            .O(N__24993),
            .I(N__24957));
    InMux I__4923 (
            .O(N__24992),
            .I(N__24957));
    InMux I__4922 (
            .O(N__24991),
            .I(N__24957));
    InMux I__4921 (
            .O(N__24988),
            .I(N__24948));
    InMux I__4920 (
            .O(N__24987),
            .I(N__24948));
    InMux I__4919 (
            .O(N__24986),
            .I(N__24948));
    InMux I__4918 (
            .O(N__24985),
            .I(N__24948));
    CascadeMux I__4917 (
            .O(N__24984),
            .I(N__24933));
    CascadeMux I__4916 (
            .O(N__24983),
            .I(N__24930));
    CascadeMux I__4915 (
            .O(N__24982),
            .I(N__24925));
    CascadeMux I__4914 (
            .O(N__24981),
            .I(N__24922));
    InMux I__4913 (
            .O(N__24980),
            .I(N__24914));
    InMux I__4912 (
            .O(N__24977),
            .I(N__24914));
    InMux I__4911 (
            .O(N__24974),
            .I(N__24914));
    InMux I__4910 (
            .O(N__24973),
            .I(N__24909));
    InMux I__4909 (
            .O(N__24972),
            .I(N__24909));
    InMux I__4908 (
            .O(N__24971),
            .I(N__24902));
    InMux I__4907 (
            .O(N__24970),
            .I(N__24902));
    InMux I__4906 (
            .O(N__24967),
            .I(N__24902));
    LocalMux I__4905 (
            .O(N__24964),
            .I(N__24897));
    LocalMux I__4904 (
            .O(N__24957),
            .I(N__24897));
    LocalMux I__4903 (
            .O(N__24948),
            .I(N__24894));
    InMux I__4902 (
            .O(N__24947),
            .I(N__24883));
    InMux I__4901 (
            .O(N__24946),
            .I(N__24883));
    InMux I__4900 (
            .O(N__24945),
            .I(N__24883));
    InMux I__4899 (
            .O(N__24944),
            .I(N__24883));
    InMux I__4898 (
            .O(N__24943),
            .I(N__24883));
    CascadeMux I__4897 (
            .O(N__24942),
            .I(N__24880));
    CascadeMux I__4896 (
            .O(N__24941),
            .I(N__24876));
    CascadeMux I__4895 (
            .O(N__24940),
            .I(N__24873));
    CascadeMux I__4894 (
            .O(N__24939),
            .I(N__24870));
    CascadeMux I__4893 (
            .O(N__24938),
            .I(N__24867));
    CascadeMux I__4892 (
            .O(N__24937),
            .I(N__24864));
    CascadeMux I__4891 (
            .O(N__24936),
            .I(N__24861));
    InMux I__4890 (
            .O(N__24933),
            .I(N__24855));
    InMux I__4889 (
            .O(N__24930),
            .I(N__24850));
    InMux I__4888 (
            .O(N__24929),
            .I(N__24850));
    InMux I__4887 (
            .O(N__24928),
            .I(N__24841));
    InMux I__4886 (
            .O(N__24925),
            .I(N__24841));
    InMux I__4885 (
            .O(N__24922),
            .I(N__24841));
    InMux I__4884 (
            .O(N__24921),
            .I(N__24841));
    LocalMux I__4883 (
            .O(N__24914),
            .I(N__24836));
    LocalMux I__4882 (
            .O(N__24909),
            .I(N__24836));
    LocalMux I__4881 (
            .O(N__24902),
            .I(N__24831));
    Span4Mux_v I__4880 (
            .O(N__24897),
            .I(N__24831));
    Span4Mux_v I__4879 (
            .O(N__24894),
            .I(N__24826));
    LocalMux I__4878 (
            .O(N__24883),
            .I(N__24826));
    InMux I__4877 (
            .O(N__24880),
            .I(N__24823));
    InMux I__4876 (
            .O(N__24879),
            .I(N__24816));
    InMux I__4875 (
            .O(N__24876),
            .I(N__24816));
    InMux I__4874 (
            .O(N__24873),
            .I(N__24816));
    InMux I__4873 (
            .O(N__24870),
            .I(N__24801));
    InMux I__4872 (
            .O(N__24867),
            .I(N__24801));
    InMux I__4871 (
            .O(N__24864),
            .I(N__24801));
    InMux I__4870 (
            .O(N__24861),
            .I(N__24801));
    InMux I__4869 (
            .O(N__24860),
            .I(N__24801));
    InMux I__4868 (
            .O(N__24859),
            .I(N__24801));
    InMux I__4867 (
            .O(N__24858),
            .I(N__24801));
    LocalMux I__4866 (
            .O(N__24855),
            .I(N__24796));
    LocalMux I__4865 (
            .O(N__24850),
            .I(N__24796));
    LocalMux I__4864 (
            .O(N__24841),
            .I(N__24793));
    Span4Mux_v I__4863 (
            .O(N__24836),
            .I(N__24786));
    Span4Mux_v I__4862 (
            .O(N__24831),
            .I(N__24786));
    Span4Mux_v I__4861 (
            .O(N__24826),
            .I(N__24786));
    LocalMux I__4860 (
            .O(N__24823),
            .I(pid_altitude_dv));
    LocalMux I__4859 (
            .O(N__24816),
            .I(pid_altitude_dv));
    LocalMux I__4858 (
            .O(N__24801),
            .I(pid_altitude_dv));
    Odrv4 I__4857 (
            .O(N__24796),
            .I(pid_altitude_dv));
    Odrv12 I__4856 (
            .O(N__24793),
            .I(pid_altitude_dv));
    Odrv4 I__4855 (
            .O(N__24786),
            .I(pid_altitude_dv));
    InMux I__4854 (
            .O(N__24773),
            .I(N__24770));
    LocalMux I__4853 (
            .O(N__24770),
            .I(N__24765));
    InMux I__4852 (
            .O(N__24769),
            .I(N__24762));
    InMux I__4851 (
            .O(N__24768),
            .I(N__24759));
    Span4Mux_s2_v I__4850 (
            .O(N__24765),
            .I(N__24756));
    LocalMux I__4849 (
            .O(N__24762),
            .I(N__24753));
    LocalMux I__4848 (
            .O(N__24759),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv4 I__4847 (
            .O(N__24756),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv12 I__4846 (
            .O(N__24753),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__4845 (
            .O(N__24746),
            .I(N__24743));
    LocalMux I__4844 (
            .O(N__24743),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    InMux I__4843 (
            .O(N__24740),
            .I(N__24734));
    InMux I__4842 (
            .O(N__24739),
            .I(N__24729));
    InMux I__4841 (
            .O(N__24738),
            .I(N__24729));
    InMux I__4840 (
            .O(N__24737),
            .I(N__24726));
    LocalMux I__4839 (
            .O(N__24734),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__4838 (
            .O(N__24729),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__4837 (
            .O(N__24726),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    CascadeMux I__4836 (
            .O(N__24719),
            .I(\ppm_encoder_1.N_140_0_cascade_ ));
    InMux I__4835 (
            .O(N__24716),
            .I(N__24713));
    LocalMux I__4834 (
            .O(N__24713),
            .I(\ppm_encoder_1.N_145 ));
    IoInMux I__4833 (
            .O(N__24710),
            .I(N__24707));
    LocalMux I__4832 (
            .O(N__24707),
            .I(N__24704));
    Span4Mux_s0_v I__4831 (
            .O(N__24704),
            .I(N__24701));
    Sp12to4 I__4830 (
            .O(N__24701),
            .I(N__24698));
    Span12Mux_h I__4829 (
            .O(N__24698),
            .I(N__24695));
    Span12Mux_v I__4828 (
            .O(N__24695),
            .I(N__24692));
    Span12Mux_v I__4827 (
            .O(N__24692),
            .I(N__24688));
    InMux I__4826 (
            .O(N__24691),
            .I(N__24685));
    Odrv12 I__4825 (
            .O(N__24688),
            .I(ppm_output_c));
    LocalMux I__4824 (
            .O(N__24685),
            .I(ppm_output_c));
    InMux I__4823 (
            .O(N__24680),
            .I(N__24677));
    LocalMux I__4822 (
            .O(N__24677),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    InMux I__4821 (
            .O(N__24674),
            .I(N__24671));
    LocalMux I__4820 (
            .O(N__24671),
            .I(N__24668));
    Odrv4 I__4819 (
            .O(N__24668),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__4818 (
            .O(N__24665),
            .I(N__24662));
    LocalMux I__4817 (
            .O(N__24662),
            .I(N__24659));
    Odrv4 I__4816 (
            .O(N__24659),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    InMux I__4815 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__4814 (
            .O(N__24653),
            .I(N__24649));
    InMux I__4813 (
            .O(N__24652),
            .I(N__24646));
    Span4Mux_h I__4812 (
            .O(N__24649),
            .I(N__24643));
    LocalMux I__4811 (
            .O(N__24646),
            .I(N__24640));
    Sp12to4 I__4810 (
            .O(N__24643),
            .I(N__24635));
    Sp12to4 I__4809 (
            .O(N__24640),
            .I(N__24635));
    Odrv12 I__4808 (
            .O(N__24635),
            .I(scaler_2_data_6));
    InMux I__4807 (
            .O(N__24632),
            .I(N__24629));
    LocalMux I__4806 (
            .O(N__24629),
            .I(N__24626));
    Span4Mux_h I__4805 (
            .O(N__24626),
            .I(N__24623));
    Span4Mux_v I__4804 (
            .O(N__24623),
            .I(N__24618));
    InMux I__4803 (
            .O(N__24622),
            .I(N__24613));
    InMux I__4802 (
            .O(N__24621),
            .I(N__24613));
    Odrv4 I__4801 (
            .O(N__24618),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__4800 (
            .O(N__24613),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    CascadeMux I__4799 (
            .O(N__24608),
            .I(N__24603));
    InMux I__4798 (
            .O(N__24607),
            .I(N__24600));
    InMux I__4797 (
            .O(N__24606),
            .I(N__24595));
    InMux I__4796 (
            .O(N__24603),
            .I(N__24595));
    LocalMux I__4795 (
            .O(N__24600),
            .I(N__24592));
    LocalMux I__4794 (
            .O(N__24595),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__4793 (
            .O(N__24592),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__4792 (
            .O(N__24587),
            .I(N__24584));
    LocalMux I__4791 (
            .O(N__24584),
            .I(N__24581));
    Span4Mux_v I__4790 (
            .O(N__24581),
            .I(N__24577));
    InMux I__4789 (
            .O(N__24580),
            .I(N__24574));
    Span4Mux_h I__4788 (
            .O(N__24577),
            .I(N__24568));
    LocalMux I__4787 (
            .O(N__24574),
            .I(N__24568));
    InMux I__4786 (
            .O(N__24573),
            .I(N__24565));
    Odrv4 I__4785 (
            .O(N__24568),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__4784 (
            .O(N__24565),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__4783 (
            .O(N__24560),
            .I(N__24556));
    CascadeMux I__4782 (
            .O(N__24559),
            .I(N__24552));
    LocalMux I__4781 (
            .O(N__24556),
            .I(N__24549));
    InMux I__4780 (
            .O(N__24555),
            .I(N__24544));
    InMux I__4779 (
            .O(N__24552),
            .I(N__24544));
    Span4Mux_v I__4778 (
            .O(N__24549),
            .I(N__24541));
    LocalMux I__4777 (
            .O(N__24544),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__4776 (
            .O(N__24541),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__4775 (
            .O(N__24536),
            .I(N__24533));
    LocalMux I__4774 (
            .O(N__24533),
            .I(N__24530));
    Span4Mux_h I__4773 (
            .O(N__24530),
            .I(N__24527));
    Span4Mux_v I__4772 (
            .O(N__24527),
            .I(N__24523));
    InMux I__4771 (
            .O(N__24526),
            .I(N__24520));
    Odrv4 I__4770 (
            .O(N__24523),
            .I(throttle_command_0));
    LocalMux I__4769 (
            .O(N__24520),
            .I(throttle_command_0));
    InMux I__4768 (
            .O(N__24515),
            .I(N__24509));
    InMux I__4767 (
            .O(N__24514),
            .I(N__24509));
    LocalMux I__4766 (
            .O(N__24509),
            .I(N__24504));
    InMux I__4765 (
            .O(N__24508),
            .I(N__24499));
    InMux I__4764 (
            .O(N__24507),
            .I(N__24499));
    Span4Mux_h I__4763 (
            .O(N__24504),
            .I(N__24496));
    LocalMux I__4762 (
            .O(N__24499),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    Odrv4 I__4761 (
            .O(N__24496),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    InMux I__4760 (
            .O(N__24491),
            .I(N__24488));
    LocalMux I__4759 (
            .O(N__24488),
            .I(N__24485));
    Span4Mux_v I__4758 (
            .O(N__24485),
            .I(N__24482));
    Span4Mux_v I__4757 (
            .O(N__24482),
            .I(N__24479));
    Odrv4 I__4756 (
            .O(N__24479),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    InMux I__4755 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__4754 (
            .O(N__24473),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__4753 (
            .O(N__24470),
            .I(\ppm_encoder_1.un1_elevator_cry_7 ));
    CascadeMux I__4752 (
            .O(N__24467),
            .I(N__24464));
    InMux I__4751 (
            .O(N__24464),
            .I(N__24461));
    LocalMux I__4750 (
            .O(N__24461),
            .I(N__24458));
    Span4Mux_v I__4749 (
            .O(N__24458),
            .I(N__24455));
    Odrv4 I__4748 (
            .O(N__24455),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__4747 (
            .O(N__24452),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__4746 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__4745 (
            .O(N__24446),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__4744 (
            .O(N__24443),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__4743 (
            .O(N__24440),
            .I(N__24437));
    LocalMux I__4742 (
            .O(N__24437),
            .I(N__24434));
    Odrv4 I__4741 (
            .O(N__24434),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__4740 (
            .O(N__24431),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__4739 (
            .O(N__24428),
            .I(N__24425));
    LocalMux I__4738 (
            .O(N__24425),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__4737 (
            .O(N__24422),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__4736 (
            .O(N__24419),
            .I(N__24416));
    LocalMux I__4735 (
            .O(N__24416),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__4734 (
            .O(N__24413),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__4733 (
            .O(N__24410),
            .I(bfn_5_23_0_));
    InMux I__4732 (
            .O(N__24407),
            .I(N__24404));
    LocalMux I__4731 (
            .O(N__24404),
            .I(N__24400));
    InMux I__4730 (
            .O(N__24403),
            .I(N__24397));
    Span4Mux_v I__4729 (
            .O(N__24400),
            .I(N__24392));
    LocalMux I__4728 (
            .O(N__24397),
            .I(N__24392));
    Span4Mux_h I__4727 (
            .O(N__24392),
            .I(N__24389));
    Odrv4 I__4726 (
            .O(N__24389),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    CascadeMux I__4725 (
            .O(N__24386),
            .I(N__24382));
    InMux I__4724 (
            .O(N__24385),
            .I(N__24378));
    InMux I__4723 (
            .O(N__24382),
            .I(N__24375));
    InMux I__4722 (
            .O(N__24381),
            .I(N__24371));
    LocalMux I__4721 (
            .O(N__24378),
            .I(N__24368));
    LocalMux I__4720 (
            .O(N__24375),
            .I(N__24365));
    InMux I__4719 (
            .O(N__24374),
            .I(N__24362));
    LocalMux I__4718 (
            .O(N__24371),
            .I(N__24359));
    Span4Mux_h I__4717 (
            .O(N__24368),
            .I(N__24352));
    Span4Mux_h I__4716 (
            .O(N__24365),
            .I(N__24352));
    LocalMux I__4715 (
            .O(N__24362),
            .I(N__24352));
    Span4Mux_h I__4714 (
            .O(N__24359),
            .I(N__24349));
    Odrv4 I__4713 (
            .O(N__24352),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__4712 (
            .O(N__24349),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__4711 (
            .O(N__24344),
            .I(N__24341));
    LocalMux I__4710 (
            .O(N__24341),
            .I(N__24338));
    Odrv4 I__4709 (
            .O(N__24338),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__4708 (
            .O(N__24335),
            .I(N__24332));
    LocalMux I__4707 (
            .O(N__24332),
            .I(N__24329));
    Span4Mux_v I__4706 (
            .O(N__24329),
            .I(N__24324));
    InMux I__4705 (
            .O(N__24328),
            .I(N__24321));
    InMux I__4704 (
            .O(N__24327),
            .I(N__24318));
    Span4Mux_s2_h I__4703 (
            .O(N__24324),
            .I(N__24315));
    LocalMux I__4702 (
            .O(N__24321),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    LocalMux I__4701 (
            .O(N__24318),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    Odrv4 I__4700 (
            .O(N__24315),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    CascadeMux I__4699 (
            .O(N__24308),
            .I(N__24305));
    InMux I__4698 (
            .O(N__24305),
            .I(N__24302));
    LocalMux I__4697 (
            .O(N__24302),
            .I(N__24297));
    InMux I__4696 (
            .O(N__24301),
            .I(N__24294));
    InMux I__4695 (
            .O(N__24300),
            .I(N__24291));
    Span4Mux_h I__4694 (
            .O(N__24297),
            .I(N__24288));
    LocalMux I__4693 (
            .O(N__24294),
            .I(N__24285));
    LocalMux I__4692 (
            .O(N__24291),
            .I(N__24282));
    Span4Mux_v I__4691 (
            .O(N__24288),
            .I(N__24279));
    Span4Mux_s2_v I__4690 (
            .O(N__24285),
            .I(N__24276));
    Span12Mux_v I__4689 (
            .O(N__24282),
            .I(N__24273));
    Odrv4 I__4688 (
            .O(N__24279),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__4687 (
            .O(N__24276),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv12 I__4686 (
            .O(N__24273),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__4685 (
            .O(N__24266),
            .I(N__24263));
    LocalMux I__4684 (
            .O(N__24263),
            .I(N__24260));
    Span4Mux_v I__4683 (
            .O(N__24260),
            .I(N__24255));
    InMux I__4682 (
            .O(N__24259),
            .I(N__24252));
    InMux I__4681 (
            .O(N__24258),
            .I(N__24249));
    Span4Mux_v I__4680 (
            .O(N__24255),
            .I(N__24244));
    LocalMux I__4679 (
            .O(N__24252),
            .I(N__24244));
    LocalMux I__4678 (
            .O(N__24249),
            .I(N__24241));
    Odrv4 I__4677 (
            .O(N__24244),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    Odrv4 I__4676 (
            .O(N__24241),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    CascadeMux I__4675 (
            .O(N__24236),
            .I(N__24233));
    InMux I__4674 (
            .O(N__24233),
            .I(N__24230));
    LocalMux I__4673 (
            .O(N__24230),
            .I(N__24227));
    Span4Mux_h I__4672 (
            .O(N__24227),
            .I(N__24222));
    InMux I__4671 (
            .O(N__24226),
            .I(N__24217));
    InMux I__4670 (
            .O(N__24225),
            .I(N__24217));
    Odrv4 I__4669 (
            .O(N__24222),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    LocalMux I__4668 (
            .O(N__24217),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    InMux I__4667 (
            .O(N__24212),
            .I(N__24209));
    LocalMux I__4666 (
            .O(N__24209),
            .I(N__24206));
    Sp12to4 I__4665 (
            .O(N__24206),
            .I(N__24203));
    Odrv12 I__4664 (
            .O(N__24203),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__4663 (
            .O(N__24200),
            .I(N__24196));
    InMux I__4662 (
            .O(N__24199),
            .I(N__24193));
    LocalMux I__4661 (
            .O(N__24196),
            .I(N__24190));
    LocalMux I__4660 (
            .O(N__24193),
            .I(N__24187));
    Span4Mux_v I__4659 (
            .O(N__24190),
            .I(N__24184));
    Span12Mux_v I__4658 (
            .O(N__24187),
            .I(N__24181));
    Odrv4 I__4657 (
            .O(N__24184),
            .I(scaler_2_data_10));
    Odrv12 I__4656 (
            .O(N__24181),
            .I(scaler_2_data_10));
    InMux I__4655 (
            .O(N__24176),
            .I(N__24173));
    LocalMux I__4654 (
            .O(N__24173),
            .I(N__24170));
    Span4Mux_h I__4653 (
            .O(N__24170),
            .I(N__24167));
    Odrv4 I__4652 (
            .O(N__24167),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__4651 (
            .O(N__24164),
            .I(N__24161));
    LocalMux I__4650 (
            .O(N__24161),
            .I(N__24157));
    InMux I__4649 (
            .O(N__24160),
            .I(N__24154));
    Span4Mux_h I__4648 (
            .O(N__24157),
            .I(N__24148));
    LocalMux I__4647 (
            .O(N__24154),
            .I(N__24148));
    InMux I__4646 (
            .O(N__24153),
            .I(N__24145));
    Span4Mux_v I__4645 (
            .O(N__24148),
            .I(N__24142));
    LocalMux I__4644 (
            .O(N__24145),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__4643 (
            .O(N__24142),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__4642 (
            .O(N__24137),
            .I(N__24134));
    LocalMux I__4641 (
            .O(N__24134),
            .I(N__24130));
    InMux I__4640 (
            .O(N__24133),
            .I(N__24127));
    Span4Mux_h I__4639 (
            .O(N__24130),
            .I(N__24122));
    LocalMux I__4638 (
            .O(N__24127),
            .I(N__24122));
    Span4Mux_v I__4637 (
            .O(N__24122),
            .I(N__24119));
    Odrv4 I__4636 (
            .O(N__24119),
            .I(scaler_2_data_13));
    InMux I__4635 (
            .O(N__24116),
            .I(N__24113));
    LocalMux I__4634 (
            .O(N__24113),
            .I(N__24110));
    Odrv12 I__4633 (
            .O(N__24110),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__4632 (
            .O(N__24107),
            .I(N__24104));
    LocalMux I__4631 (
            .O(N__24104),
            .I(N__24100));
    InMux I__4630 (
            .O(N__24103),
            .I(N__24097));
    Span4Mux_h I__4629 (
            .O(N__24100),
            .I(N__24091));
    LocalMux I__4628 (
            .O(N__24097),
            .I(N__24091));
    InMux I__4627 (
            .O(N__24096),
            .I(N__24088));
    Span4Mux_v I__4626 (
            .O(N__24091),
            .I(N__24085));
    LocalMux I__4625 (
            .O(N__24088),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__4624 (
            .O(N__24085),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__4623 (
            .O(N__24080),
            .I(N__24077));
    LocalMux I__4622 (
            .O(N__24077),
            .I(N__24074));
    Span4Mux_h I__4621 (
            .O(N__24074),
            .I(N__24071));
    Odrv4 I__4620 (
            .O(N__24071),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__4619 (
            .O(N__24068),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__4618 (
            .O(N__24065),
            .I(N__24059));
    InMux I__4617 (
            .O(N__24064),
            .I(N__24054));
    InMux I__4616 (
            .O(N__24063),
            .I(N__24054));
    InMux I__4615 (
            .O(N__24062),
            .I(N__24051));
    LocalMux I__4614 (
            .O(N__24059),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__4613 (
            .O(N__24054),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__4612 (
            .O(N__24051),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    CascadeMux I__4611 (
            .O(N__24044),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ));
    InMux I__4610 (
            .O(N__24041),
            .I(N__24035));
    InMux I__4609 (
            .O(N__24040),
            .I(N__24035));
    LocalMux I__4608 (
            .O(N__24035),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_1 ));
    CascadeMux I__4607 (
            .O(N__24032),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ));
    CascadeMux I__4606 (
            .O(N__24029),
            .I(N__24025));
    InMux I__4605 (
            .O(N__24028),
            .I(N__24021));
    InMux I__4604 (
            .O(N__24025),
            .I(N__24018));
    InMux I__4603 (
            .O(N__24024),
            .I(N__24015));
    LocalMux I__4602 (
            .O(N__24021),
            .I(N__24012));
    LocalMux I__4601 (
            .O(N__24018),
            .I(N__24009));
    LocalMux I__4600 (
            .O(N__24015),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv4 I__4599 (
            .O(N__24012),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv4 I__4598 (
            .O(N__24009),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__4597 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__4596 (
            .O(N__23999),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3 ));
    InMux I__4595 (
            .O(N__23996),
            .I(N__23992));
    IoInMux I__4594 (
            .O(N__23995),
            .I(N__23989));
    LocalMux I__4593 (
            .O(N__23992),
            .I(N__23986));
    LocalMux I__4592 (
            .O(N__23989),
            .I(N__23982));
    Span4Mux_v I__4591 (
            .O(N__23986),
            .I(N__23978));
    InMux I__4590 (
            .O(N__23985),
            .I(N__23975));
    Span12Mux_s9_v I__4589 (
            .O(N__23982),
            .I(N__23972));
    InMux I__4588 (
            .O(N__23981),
            .I(N__23969));
    Span4Mux_v I__4587 (
            .O(N__23978),
            .I(N__23964));
    LocalMux I__4586 (
            .O(N__23975),
            .I(N__23964));
    Odrv12 I__4585 (
            .O(N__23972),
            .I(debug_CH1_0A_c));
    LocalMux I__4584 (
            .O(N__23969),
            .I(debug_CH1_0A_c));
    Odrv4 I__4583 (
            .O(N__23964),
            .I(debug_CH1_0A_c));
    InMux I__4582 (
            .O(N__23957),
            .I(N__23944));
    InMux I__4581 (
            .O(N__23956),
            .I(N__23941));
    CascadeMux I__4580 (
            .O(N__23955),
            .I(N__23936));
    CascadeMux I__4579 (
            .O(N__23954),
            .I(N__23933));
    InMux I__4578 (
            .O(N__23953),
            .I(N__23917));
    InMux I__4577 (
            .O(N__23952),
            .I(N__23917));
    InMux I__4576 (
            .O(N__23951),
            .I(N__23917));
    InMux I__4575 (
            .O(N__23950),
            .I(N__23917));
    InMux I__4574 (
            .O(N__23949),
            .I(N__23917));
    InMux I__4573 (
            .O(N__23948),
            .I(N__23917));
    InMux I__4572 (
            .O(N__23947),
            .I(N__23917));
    LocalMux I__4571 (
            .O(N__23944),
            .I(N__23914));
    LocalMux I__4570 (
            .O(N__23941),
            .I(N__23909));
    InMux I__4569 (
            .O(N__23940),
            .I(N__23898));
    InMux I__4568 (
            .O(N__23939),
            .I(N__23898));
    InMux I__4567 (
            .O(N__23936),
            .I(N__23898));
    InMux I__4566 (
            .O(N__23933),
            .I(N__23898));
    InMux I__4565 (
            .O(N__23932),
            .I(N__23898));
    LocalMux I__4564 (
            .O(N__23917),
            .I(N__23895));
    Span4Mux_v I__4563 (
            .O(N__23914),
            .I(N__23892));
    InMux I__4562 (
            .O(N__23913),
            .I(N__23887));
    InMux I__4561 (
            .O(N__23912),
            .I(N__23887));
    Span4Mux_v I__4560 (
            .O(N__23909),
            .I(N__23882));
    LocalMux I__4559 (
            .O(N__23898),
            .I(N__23879));
    Span4Mux_v I__4558 (
            .O(N__23895),
            .I(N__23872));
    Span4Mux_v I__4557 (
            .O(N__23892),
            .I(N__23872));
    LocalMux I__4556 (
            .O(N__23887),
            .I(N__23872));
    InMux I__4555 (
            .O(N__23886),
            .I(N__23864));
    InMux I__4554 (
            .O(N__23885),
            .I(N__23861));
    Span4Mux_v I__4553 (
            .O(N__23882),
            .I(N__23858));
    Span4Mux_v I__4552 (
            .O(N__23879),
            .I(N__23853));
    Span4Mux_v I__4551 (
            .O(N__23872),
            .I(N__23853));
    InMux I__4550 (
            .O(N__23871),
            .I(N__23846));
    InMux I__4549 (
            .O(N__23870),
            .I(N__23846));
    InMux I__4548 (
            .O(N__23869),
            .I(N__23846));
    InMux I__4547 (
            .O(N__23868),
            .I(N__23843));
    InMux I__4546 (
            .O(N__23867),
            .I(N__23840));
    LocalMux I__4545 (
            .O(N__23864),
            .I(\pid_alt.N_60_i ));
    LocalMux I__4544 (
            .O(N__23861),
            .I(\pid_alt.N_60_i ));
    Odrv4 I__4543 (
            .O(N__23858),
            .I(\pid_alt.N_60_i ));
    Odrv4 I__4542 (
            .O(N__23853),
            .I(\pid_alt.N_60_i ));
    LocalMux I__4541 (
            .O(N__23846),
            .I(\pid_alt.N_60_i ));
    LocalMux I__4540 (
            .O(N__23843),
            .I(\pid_alt.N_60_i ));
    LocalMux I__4539 (
            .O(N__23840),
            .I(\pid_alt.N_60_i ));
    InMux I__4538 (
            .O(N__23825),
            .I(N__23822));
    LocalMux I__4537 (
            .O(N__23822),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    InMux I__4536 (
            .O(N__23819),
            .I(N__23814));
    InMux I__4535 (
            .O(N__23818),
            .I(N__23811));
    CascadeMux I__4534 (
            .O(N__23817),
            .I(N__23808));
    LocalMux I__4533 (
            .O(N__23814),
            .I(N__23805));
    LocalMux I__4532 (
            .O(N__23811),
            .I(N__23801));
    InMux I__4531 (
            .O(N__23808),
            .I(N__23798));
    Span4Mux_v I__4530 (
            .O(N__23805),
            .I(N__23795));
    InMux I__4529 (
            .O(N__23804),
            .I(N__23792));
    Span12Mux_v I__4528 (
            .O(N__23801),
            .I(N__23787));
    LocalMux I__4527 (
            .O(N__23798),
            .I(N__23787));
    Odrv4 I__4526 (
            .O(N__23795),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__4525 (
            .O(N__23792),
            .I(frame_decoder_OFF2data_0));
    Odrv12 I__4524 (
            .O(N__23787),
            .I(frame_decoder_OFF2data_0));
    InMux I__4523 (
            .O(N__23780),
            .I(N__23776));
    InMux I__4522 (
            .O(N__23779),
            .I(N__23773));
    LocalMux I__4521 (
            .O(N__23776),
            .I(N__23770));
    LocalMux I__4520 (
            .O(N__23773),
            .I(N__23766));
    Span4Mux_v I__4519 (
            .O(N__23770),
            .I(N__23763));
    InMux I__4518 (
            .O(N__23769),
            .I(N__23759));
    Span4Mux_v I__4517 (
            .O(N__23766),
            .I(N__23754));
    Span4Mux_h I__4516 (
            .O(N__23763),
            .I(N__23754));
    InMux I__4515 (
            .O(N__23762),
            .I(N__23751));
    LocalMux I__4514 (
            .O(N__23759),
            .I(N__23748));
    Odrv4 I__4513 (
            .O(N__23754),
            .I(frame_decoder_CH2data_0));
    LocalMux I__4512 (
            .O(N__23751),
            .I(frame_decoder_CH2data_0));
    Odrv4 I__4511 (
            .O(N__23748),
            .I(frame_decoder_CH2data_0));
    InMux I__4510 (
            .O(N__23741),
            .I(N__23738));
    LocalMux I__4509 (
            .O(N__23738),
            .I(N__23734));
    CascadeMux I__4508 (
            .O(N__23737),
            .I(N__23731));
    Span4Mux_v I__4507 (
            .O(N__23734),
            .I(N__23728));
    InMux I__4506 (
            .O(N__23731),
            .I(N__23725));
    Odrv4 I__4505 (
            .O(N__23728),
            .I(scaler_2_data_4));
    LocalMux I__4504 (
            .O(N__23725),
            .I(scaler_2_data_4));
    InMux I__4503 (
            .O(N__23720),
            .I(N__23717));
    LocalMux I__4502 (
            .O(N__23717),
            .I(N__23714));
    Span4Mux_h I__4501 (
            .O(N__23714),
            .I(N__23711));
    Odrv4 I__4500 (
            .O(N__23711),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ));
    InMux I__4499 (
            .O(N__23708),
            .I(N__23705));
    LocalMux I__4498 (
            .O(N__23705),
            .I(N__23701));
    InMux I__4497 (
            .O(N__23704),
            .I(N__23698));
    Odrv4 I__4496 (
            .O(N__23701),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ));
    LocalMux I__4495 (
            .O(N__23698),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ));
    InMux I__4494 (
            .O(N__23693),
            .I(N__23690));
    LocalMux I__4493 (
            .O(N__23690),
            .I(N__23685));
    InMux I__4492 (
            .O(N__23689),
            .I(N__23682));
    InMux I__4491 (
            .O(N__23688),
            .I(N__23679));
    Span4Mux_h I__4490 (
            .O(N__23685),
            .I(N__23676));
    LocalMux I__4489 (
            .O(N__23682),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    LocalMux I__4488 (
            .O(N__23679),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__4487 (
            .O(N__23676),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    InMux I__4486 (
            .O(N__23669),
            .I(N__23666));
    LocalMux I__4485 (
            .O(N__23666),
            .I(N__23663));
    Odrv4 I__4484 (
            .O(N__23663),
            .I(frame_decoder_OFF2data_5));
    InMux I__4483 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__4482 (
            .O(N__23657),
            .I(N__23654));
    Odrv4 I__4481 (
            .O(N__23654),
            .I(frame_decoder_OFF2data_6));
    InMux I__4480 (
            .O(N__23651),
            .I(N__23645));
    InMux I__4479 (
            .O(N__23650),
            .I(N__23645));
    LocalMux I__4478 (
            .O(N__23645),
            .I(frame_decoder_OFF2data_7));
    CEMux I__4477 (
            .O(N__23642),
            .I(N__23639));
    LocalMux I__4476 (
            .O(N__23639),
            .I(N__23636));
    Span4Mux_v I__4475 (
            .O(N__23636),
            .I(N__23633));
    Span4Mux_h I__4474 (
            .O(N__23633),
            .I(N__23630));
    Odrv4 I__4473 (
            .O(N__23630),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    CascadeMux I__4472 (
            .O(N__23627),
            .I(N__23624));
    InMux I__4471 (
            .O(N__23624),
            .I(N__23621));
    LocalMux I__4470 (
            .O(N__23621),
            .I(\dron_frame_decoder_1.state_RNO_1Z0Z_0 ));
    InMux I__4469 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__4468 (
            .O(N__23615),
            .I(N__23612));
    Odrv4 I__4467 (
            .O(N__23612),
            .I(\dron_frame_decoder_1.N_194_4 ));
    CascadeMux I__4466 (
            .O(N__23609),
            .I(N__23606));
    InMux I__4465 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__4464 (
            .O(N__23603),
            .I(N__23600));
    Odrv4 I__4463 (
            .O(N__23600),
            .I(\dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ));
    InMux I__4462 (
            .O(N__23597),
            .I(N__23594));
    LocalMux I__4461 (
            .O(N__23594),
            .I(\dron_frame_decoder_1.state_RNO_0Z0Z_0 ));
    CascadeMux I__4460 (
            .O(N__23591),
            .I(N__23588));
    InMux I__4459 (
            .O(N__23588),
            .I(N__23585));
    LocalMux I__4458 (
            .O(N__23585),
            .I(N__23582));
    Odrv12 I__4457 (
            .O(N__23582),
            .I(alt_command_5));
    CascadeMux I__4456 (
            .O(N__23579),
            .I(N__23576));
    InMux I__4455 (
            .O(N__23576),
            .I(N__23573));
    LocalMux I__4454 (
            .O(N__23573),
            .I(N__23570));
    Odrv4 I__4453 (
            .O(N__23570),
            .I(alt_command_6));
    CascadeMux I__4452 (
            .O(N__23567),
            .I(N__23564));
    InMux I__4451 (
            .O(N__23564),
            .I(N__23561));
    LocalMux I__4450 (
            .O(N__23561),
            .I(N__23558));
    Odrv4 I__4449 (
            .O(N__23558),
            .I(alt_command_7));
    CEMux I__4448 (
            .O(N__23555),
            .I(N__23552));
    LocalMux I__4447 (
            .O(N__23552),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    CascadeMux I__4446 (
            .O(N__23549),
            .I(N__23546));
    InMux I__4445 (
            .O(N__23546),
            .I(N__23543));
    LocalMux I__4444 (
            .O(N__23543),
            .I(N__23540));
    Odrv12 I__4443 (
            .O(N__23540),
            .I(frame_decoder_OFF2data_1));
    CascadeMux I__4442 (
            .O(N__23537),
            .I(N__23534));
    InMux I__4441 (
            .O(N__23534),
            .I(N__23531));
    LocalMux I__4440 (
            .O(N__23531),
            .I(N__23528));
    Odrv4 I__4439 (
            .O(N__23528),
            .I(frame_decoder_OFF2data_2));
    CascadeMux I__4438 (
            .O(N__23525),
            .I(N__23522));
    InMux I__4437 (
            .O(N__23522),
            .I(N__23519));
    LocalMux I__4436 (
            .O(N__23519),
            .I(N__23516));
    Odrv4 I__4435 (
            .O(N__23516),
            .I(frame_decoder_OFF2data_3));
    InMux I__4434 (
            .O(N__23513),
            .I(N__23510));
    LocalMux I__4433 (
            .O(N__23510),
            .I(N__23507));
    Span4Mux_s3_h I__4432 (
            .O(N__23507),
            .I(N__23504));
    Odrv4 I__4431 (
            .O(N__23504),
            .I(frame_decoder_OFF2data_4));
    InMux I__4430 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__4429 (
            .O(N__23498),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    InMux I__4428 (
            .O(N__23495),
            .I(N__23492));
    LocalMux I__4427 (
            .O(N__23492),
            .I(N__23489));
    Odrv4 I__4426 (
            .O(N__23489),
            .I(drone_altitude_i_4));
    InMux I__4425 (
            .O(N__23486),
            .I(N__23483));
    LocalMux I__4424 (
            .O(N__23483),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__4423 (
            .O(N__23480),
            .I(N__23477));
    LocalMux I__4422 (
            .O(N__23477),
            .I(N__23474));
    Odrv4 I__4421 (
            .O(N__23474),
            .I(drone_altitude_i_5));
    InMux I__4420 (
            .O(N__23471),
            .I(N__23468));
    LocalMux I__4419 (
            .O(N__23468),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__4418 (
            .O(N__23465),
            .I(N__23462));
    LocalMux I__4417 (
            .O(N__23462),
            .I(N__23459));
    Odrv4 I__4416 (
            .O(N__23459),
            .I(drone_altitude_i_6));
    CascadeMux I__4415 (
            .O(N__23456),
            .I(N__23453));
    InMux I__4414 (
            .O(N__23453),
            .I(N__23450));
    LocalMux I__4413 (
            .O(N__23450),
            .I(N__23447));
    Span4Mux_s3_h I__4412 (
            .O(N__23447),
            .I(N__23444));
    Odrv4 I__4411 (
            .O(N__23444),
            .I(alt_command_4));
    InMux I__4410 (
            .O(N__23441),
            .I(N__23438));
    LocalMux I__4409 (
            .O(N__23438),
            .I(N__23435));
    Span4Mux_v I__4408 (
            .O(N__23435),
            .I(N__23432));
    Odrv4 I__4407 (
            .O(N__23432),
            .I(\ppm_encoder_1.N_301 ));
    InMux I__4406 (
            .O(N__23429),
            .I(N__23426));
    LocalMux I__4405 (
            .O(N__23426),
            .I(N__23423));
    Span4Mux_h I__4404 (
            .O(N__23423),
            .I(N__23418));
    InMux I__4403 (
            .O(N__23422),
            .I(N__23413));
    InMux I__4402 (
            .O(N__23421),
            .I(N__23413));
    Odrv4 I__4401 (
            .O(N__23418),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__4400 (
            .O(N__23413),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__4399 (
            .O(N__23408),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ));
    InMux I__4398 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__4397 (
            .O(N__23402),
            .I(N__23399));
    Span4Mux_s3_v I__4396 (
            .O(N__23399),
            .I(N__23396));
    Odrv4 I__4395 (
            .O(N__23396),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ));
    CascadeMux I__4394 (
            .O(N__23393),
            .I(N__23390));
    InMux I__4393 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__4392 (
            .O(N__23387),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    CascadeMux I__4391 (
            .O(N__23384),
            .I(N__23381));
    InMux I__4390 (
            .O(N__23381),
            .I(N__23378));
    LocalMux I__4389 (
            .O(N__23378),
            .I(N__23375));
    Span4Mux_v I__4388 (
            .O(N__23375),
            .I(N__23372));
    Odrv4 I__4387 (
            .O(N__23372),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    CascadeMux I__4386 (
            .O(N__23369),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ));
    InMux I__4385 (
            .O(N__23366),
            .I(N__23363));
    LocalMux I__4384 (
            .O(N__23363),
            .I(N__23358));
    InMux I__4383 (
            .O(N__23362),
            .I(N__23353));
    InMux I__4382 (
            .O(N__23361),
            .I(N__23353));
    Odrv4 I__4381 (
            .O(N__23358),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__4380 (
            .O(N__23353),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__4379 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__4378 (
            .O(N__23345),
            .I(N__23342));
    Odrv4 I__4377 (
            .O(N__23342),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    InMux I__4376 (
            .O(N__23339),
            .I(N__23334));
    InMux I__4375 (
            .O(N__23338),
            .I(N__23331));
    InMux I__4374 (
            .O(N__23337),
            .I(N__23328));
    LocalMux I__4373 (
            .O(N__23334),
            .I(N__23325));
    LocalMux I__4372 (
            .O(N__23331),
            .I(N__23322));
    LocalMux I__4371 (
            .O(N__23328),
            .I(N__23319));
    Span4Mux_h I__4370 (
            .O(N__23325),
            .I(N__23316));
    Span4Mux_s1_v I__4369 (
            .O(N__23322),
            .I(N__23309));
    Span4Mux_h I__4368 (
            .O(N__23319),
            .I(N__23309));
    Span4Mux_v I__4367 (
            .O(N__23316),
            .I(N__23309));
    Odrv4 I__4366 (
            .O(N__23309),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__4365 (
            .O(N__23306),
            .I(N__23303));
    LocalMux I__4364 (
            .O(N__23303),
            .I(N__23300));
    Odrv4 I__4363 (
            .O(N__23300),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__4362 (
            .O(N__23297),
            .I(N__23289));
    CascadeMux I__4361 (
            .O(N__23296),
            .I(N__23285));
    InMux I__4360 (
            .O(N__23295),
            .I(N__23277));
    InMux I__4359 (
            .O(N__23294),
            .I(N__23277));
    InMux I__4358 (
            .O(N__23293),
            .I(N__23277));
    InMux I__4357 (
            .O(N__23292),
            .I(N__23274));
    LocalMux I__4356 (
            .O(N__23289),
            .I(N__23271));
    InMux I__4355 (
            .O(N__23288),
            .I(N__23264));
    InMux I__4354 (
            .O(N__23285),
            .I(N__23264));
    InMux I__4353 (
            .O(N__23284),
            .I(N__23264));
    LocalMux I__4352 (
            .O(N__23277),
            .I(N__23261));
    LocalMux I__4351 (
            .O(N__23274),
            .I(N__23254));
    Span4Mux_h I__4350 (
            .O(N__23271),
            .I(N__23254));
    LocalMux I__4349 (
            .O(N__23264),
            .I(N__23254));
    Span4Mux_s3_v I__4348 (
            .O(N__23261),
            .I(N__23250));
    Span4Mux_v I__4347 (
            .O(N__23254),
            .I(N__23247));
    InMux I__4346 (
            .O(N__23253),
            .I(N__23244));
    Odrv4 I__4345 (
            .O(N__23250),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    Odrv4 I__4344 (
            .O(N__23247),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__4343 (
            .O(N__23244),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    InMux I__4342 (
            .O(N__23237),
            .I(N__23224));
    InMux I__4341 (
            .O(N__23236),
            .I(N__23219));
    InMux I__4340 (
            .O(N__23235),
            .I(N__23219));
    CascadeMux I__4339 (
            .O(N__23234),
            .I(N__23216));
    CascadeMux I__4338 (
            .O(N__23233),
            .I(N__23213));
    CascadeMux I__4337 (
            .O(N__23232),
            .I(N__23208));
    CascadeMux I__4336 (
            .O(N__23231),
            .I(N__23205));
    InMux I__4335 (
            .O(N__23230),
            .I(N__23202));
    CascadeMux I__4334 (
            .O(N__23229),
            .I(N__23198));
    CascadeMux I__4333 (
            .O(N__23228),
            .I(N__23195));
    InMux I__4332 (
            .O(N__23227),
            .I(N__23188));
    LocalMux I__4331 (
            .O(N__23224),
            .I(N__23183));
    LocalMux I__4330 (
            .O(N__23219),
            .I(N__23183));
    InMux I__4329 (
            .O(N__23216),
            .I(N__23178));
    InMux I__4328 (
            .O(N__23213),
            .I(N__23178));
    InMux I__4327 (
            .O(N__23212),
            .I(N__23173));
    InMux I__4326 (
            .O(N__23211),
            .I(N__23173));
    InMux I__4325 (
            .O(N__23208),
            .I(N__23168));
    InMux I__4324 (
            .O(N__23205),
            .I(N__23168));
    LocalMux I__4323 (
            .O(N__23202),
            .I(N__23164));
    InMux I__4322 (
            .O(N__23201),
            .I(N__23161));
    InMux I__4321 (
            .O(N__23198),
            .I(N__23156));
    InMux I__4320 (
            .O(N__23195),
            .I(N__23156));
    InMux I__4319 (
            .O(N__23194),
            .I(N__23151));
    InMux I__4318 (
            .O(N__23193),
            .I(N__23151));
    CascadeMux I__4317 (
            .O(N__23192),
            .I(N__23148));
    CascadeMux I__4316 (
            .O(N__23191),
            .I(N__23145));
    LocalMux I__4315 (
            .O(N__23188),
            .I(N__23142));
    Span4Mux_v I__4314 (
            .O(N__23183),
            .I(N__23137));
    LocalMux I__4313 (
            .O(N__23178),
            .I(N__23137));
    LocalMux I__4312 (
            .O(N__23173),
            .I(N__23132));
    LocalMux I__4311 (
            .O(N__23168),
            .I(N__23132));
    InMux I__4310 (
            .O(N__23167),
            .I(N__23129));
    Span4Mux_h I__4309 (
            .O(N__23164),
            .I(N__23122));
    LocalMux I__4308 (
            .O(N__23161),
            .I(N__23122));
    LocalMux I__4307 (
            .O(N__23156),
            .I(N__23122));
    LocalMux I__4306 (
            .O(N__23151),
            .I(N__23119));
    InMux I__4305 (
            .O(N__23148),
            .I(N__23114));
    InMux I__4304 (
            .O(N__23145),
            .I(N__23114));
    Span4Mux_s1_v I__4303 (
            .O(N__23142),
            .I(N__23105));
    Span4Mux_s1_v I__4302 (
            .O(N__23137),
            .I(N__23105));
    Span4Mux_s2_h I__4301 (
            .O(N__23132),
            .I(N__23105));
    LocalMux I__4300 (
            .O(N__23129),
            .I(N__23105));
    Odrv4 I__4299 (
            .O(N__23122),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__4298 (
            .O(N__23119),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__4297 (
            .O(N__23114),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__4296 (
            .O(N__23105),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__4295 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__4294 (
            .O(N__23093),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    CascadeMux I__4293 (
            .O(N__23090),
            .I(N__23077));
    InMux I__4292 (
            .O(N__23089),
            .I(N__23072));
    InMux I__4291 (
            .O(N__23088),
            .I(N__23069));
    InMux I__4290 (
            .O(N__23087),
            .I(N__23064));
    InMux I__4289 (
            .O(N__23086),
            .I(N__23064));
    CascadeMux I__4288 (
            .O(N__23085),
            .I(N__23056));
    CascadeMux I__4287 (
            .O(N__23084),
            .I(N__23052));
    CascadeMux I__4286 (
            .O(N__23083),
            .I(N__23048));
    InMux I__4285 (
            .O(N__23082),
            .I(N__23041));
    InMux I__4284 (
            .O(N__23081),
            .I(N__23036));
    InMux I__4283 (
            .O(N__23080),
            .I(N__23036));
    InMux I__4282 (
            .O(N__23077),
            .I(N__23031));
    InMux I__4281 (
            .O(N__23076),
            .I(N__23031));
    InMux I__4280 (
            .O(N__23075),
            .I(N__23026));
    LocalMux I__4279 (
            .O(N__23072),
            .I(N__23023));
    LocalMux I__4278 (
            .O(N__23069),
            .I(N__23018));
    LocalMux I__4277 (
            .O(N__23064),
            .I(N__23018));
    InMux I__4276 (
            .O(N__23063),
            .I(N__23011));
    InMux I__4275 (
            .O(N__23062),
            .I(N__23011));
    InMux I__4274 (
            .O(N__23061),
            .I(N__23011));
    InMux I__4273 (
            .O(N__23060),
            .I(N__23002));
    InMux I__4272 (
            .O(N__23059),
            .I(N__23002));
    InMux I__4271 (
            .O(N__23056),
            .I(N__23002));
    InMux I__4270 (
            .O(N__23055),
            .I(N__23002));
    InMux I__4269 (
            .O(N__23052),
            .I(N__22997));
    InMux I__4268 (
            .O(N__23051),
            .I(N__22997));
    InMux I__4267 (
            .O(N__23048),
            .I(N__22994));
    InMux I__4266 (
            .O(N__23047),
            .I(N__22989));
    InMux I__4265 (
            .O(N__23046),
            .I(N__22989));
    CascadeMux I__4264 (
            .O(N__23045),
            .I(N__22986));
    CascadeMux I__4263 (
            .O(N__23044),
            .I(N__22979));
    LocalMux I__4262 (
            .O(N__23041),
            .I(N__22971));
    LocalMux I__4261 (
            .O(N__23036),
            .I(N__22971));
    LocalMux I__4260 (
            .O(N__23031),
            .I(N__22971));
    InMux I__4259 (
            .O(N__23030),
            .I(N__22966));
    InMux I__4258 (
            .O(N__23029),
            .I(N__22966));
    LocalMux I__4257 (
            .O(N__23026),
            .I(N__22963));
    Span4Mux_v I__4256 (
            .O(N__23023),
            .I(N__22960));
    Span4Mux_h I__4255 (
            .O(N__23018),
            .I(N__22951));
    LocalMux I__4254 (
            .O(N__23011),
            .I(N__22951));
    LocalMux I__4253 (
            .O(N__23002),
            .I(N__22951));
    LocalMux I__4252 (
            .O(N__22997),
            .I(N__22951));
    LocalMux I__4251 (
            .O(N__22994),
            .I(N__22937));
    LocalMux I__4250 (
            .O(N__22989),
            .I(N__22937));
    InMux I__4249 (
            .O(N__22986),
            .I(N__22928));
    InMux I__4248 (
            .O(N__22985),
            .I(N__22928));
    InMux I__4247 (
            .O(N__22984),
            .I(N__22928));
    InMux I__4246 (
            .O(N__22983),
            .I(N__22928));
    InMux I__4245 (
            .O(N__22982),
            .I(N__22921));
    InMux I__4244 (
            .O(N__22979),
            .I(N__22921));
    InMux I__4243 (
            .O(N__22978),
            .I(N__22921));
    Span4Mux_s2_v I__4242 (
            .O(N__22971),
            .I(N__22916));
    LocalMux I__4241 (
            .O(N__22966),
            .I(N__22916));
    Span4Mux_v I__4240 (
            .O(N__22963),
            .I(N__22909));
    Span4Mux_v I__4239 (
            .O(N__22960),
            .I(N__22909));
    Span4Mux_v I__4238 (
            .O(N__22951),
            .I(N__22909));
    InMux I__4237 (
            .O(N__22950),
            .I(N__22902));
    InMux I__4236 (
            .O(N__22949),
            .I(N__22902));
    InMux I__4235 (
            .O(N__22948),
            .I(N__22902));
    InMux I__4234 (
            .O(N__22947),
            .I(N__22893));
    InMux I__4233 (
            .O(N__22946),
            .I(N__22893));
    InMux I__4232 (
            .O(N__22945),
            .I(N__22893));
    InMux I__4231 (
            .O(N__22944),
            .I(N__22893));
    InMux I__4230 (
            .O(N__22943),
            .I(N__22888));
    InMux I__4229 (
            .O(N__22942),
            .I(N__22888));
    Odrv4 I__4228 (
            .O(N__22937),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4227 (
            .O(N__22928),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4226 (
            .O(N__22921),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__4225 (
            .O(N__22916),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__4224 (
            .O(N__22909),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4223 (
            .O(N__22902),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4222 (
            .O(N__22893),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__4221 (
            .O(N__22888),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    InMux I__4220 (
            .O(N__22871),
            .I(N__22868));
    LocalMux I__4219 (
            .O(N__22868),
            .I(N__22865));
    Odrv4 I__4218 (
            .O(N__22865),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__4217 (
            .O(N__22862),
            .I(N__22859));
    LocalMux I__4216 (
            .O(N__22859),
            .I(N__22856));
    Odrv12 I__4215 (
            .O(N__22856),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__4214 (
            .O(N__22853),
            .I(N__22850));
    LocalMux I__4213 (
            .O(N__22850),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__4212 (
            .O(N__22847),
            .I(N__22844));
    LocalMux I__4211 (
            .O(N__22844),
            .I(N__22841));
    Span4Mux_v I__4210 (
            .O(N__22841),
            .I(N__22838));
    Span4Mux_h I__4209 (
            .O(N__22838),
            .I(N__22835));
    Span4Mux_v I__4208 (
            .O(N__22835),
            .I(N__22832));
    Odrv4 I__4207 (
            .O(N__22832),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__4206 (
            .O(N__22829),
            .I(N__22826));
    LocalMux I__4205 (
            .O(N__22826),
            .I(N__22823));
    Span4Mux_v I__4204 (
            .O(N__22823),
            .I(N__22820));
    Odrv4 I__4203 (
            .O(N__22820),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    CascadeMux I__4202 (
            .O(N__22817),
            .I(N__22814));
    InMux I__4201 (
            .O(N__22814),
            .I(N__22811));
    LocalMux I__4200 (
            .O(N__22811),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__4199 (
            .O(N__22808),
            .I(N__22805));
    LocalMux I__4198 (
            .O(N__22805),
            .I(N__22802));
    Span4Mux_v I__4197 (
            .O(N__22802),
            .I(N__22799));
    Odrv4 I__4196 (
            .O(N__22799),
            .I(\ppm_encoder_1.N_300 ));
    InMux I__4195 (
            .O(N__22796),
            .I(N__22793));
    LocalMux I__4194 (
            .O(N__22793),
            .I(N__22788));
    InMux I__4193 (
            .O(N__22792),
            .I(N__22783));
    InMux I__4192 (
            .O(N__22791),
            .I(N__22783));
    Odrv12 I__4191 (
            .O(N__22788),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__4190 (
            .O(N__22783),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__4189 (
            .O(N__22778),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__4188 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__4187 (
            .O(N__22772),
            .I(N__22768));
    InMux I__4186 (
            .O(N__22771),
            .I(N__22765));
    Span4Mux_v I__4185 (
            .O(N__22768),
            .I(N__22759));
    LocalMux I__4184 (
            .O(N__22765),
            .I(N__22759));
    InMux I__4183 (
            .O(N__22764),
            .I(N__22756));
    Span4Mux_v I__4182 (
            .O(N__22759),
            .I(N__22753));
    LocalMux I__4181 (
            .O(N__22756),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__4180 (
            .O(N__22753),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    CascadeMux I__4179 (
            .O(N__22748),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__4178 (
            .O(N__22745),
            .I(N__22742));
    LocalMux I__4177 (
            .O(N__22742),
            .I(N__22739));
    Span4Mux_h I__4176 (
            .O(N__22739),
            .I(N__22736));
    Odrv4 I__4175 (
            .O(N__22736),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    InMux I__4174 (
            .O(N__22733),
            .I(N__22730));
    LocalMux I__4173 (
            .O(N__22730),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__4172 (
            .O(N__22727),
            .I(\ppm_encoder_1.N_145_17_cascade_ ));
    CascadeMux I__4171 (
            .O(N__22724),
            .I(N__22721));
    InMux I__4170 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__4169 (
            .O(N__22718),
            .I(\ppm_encoder_1.N_145_17 ));
    CascadeMux I__4168 (
            .O(N__22715),
            .I(\ppm_encoder_1.N_238_cascade_ ));
    InMux I__4167 (
            .O(N__22712),
            .I(N__22709));
    LocalMux I__4166 (
            .O(N__22709),
            .I(N__22706));
    Span4Mux_h I__4165 (
            .O(N__22706),
            .I(N__22703));
    Odrv4 I__4164 (
            .O(N__22703),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__4163 (
            .O(N__22700),
            .I(N__22697));
    LocalMux I__4162 (
            .O(N__22697),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__4161 (
            .O(N__22694),
            .I(N__22691));
    LocalMux I__4160 (
            .O(N__22691),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__4159 (
            .O(N__22688),
            .I(N__22685));
    LocalMux I__4158 (
            .O(N__22685),
            .I(N__22682));
    Odrv12 I__4157 (
            .O(N__22682),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__4156 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__4155 (
            .O(N__22676),
            .I(N__22673));
    Span4Mux_h I__4154 (
            .O(N__22673),
            .I(N__22670));
    Odrv4 I__4153 (
            .O(N__22670),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    CascadeMux I__4152 (
            .O(N__22667),
            .I(N__22664));
    InMux I__4151 (
            .O(N__22664),
            .I(N__22661));
    LocalMux I__4150 (
            .O(N__22661),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    CascadeMux I__4149 (
            .O(N__22658),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ));
    CascadeMux I__4148 (
            .O(N__22655),
            .I(N__22652));
    InMux I__4147 (
            .O(N__22652),
            .I(N__22649));
    LocalMux I__4146 (
            .O(N__22649),
            .I(N__22646));
    Span4Mux_h I__4145 (
            .O(N__22646),
            .I(N__22643));
    Odrv4 I__4144 (
            .O(N__22643),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ));
    InMux I__4143 (
            .O(N__22640),
            .I(N__22636));
    InMux I__4142 (
            .O(N__22639),
            .I(N__22633));
    LocalMux I__4141 (
            .O(N__22636),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    LocalMux I__4140 (
            .O(N__22633),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    InMux I__4139 (
            .O(N__22628),
            .I(N__22624));
    InMux I__4138 (
            .O(N__22627),
            .I(N__22621));
    LocalMux I__4137 (
            .O(N__22624),
            .I(N__22618));
    LocalMux I__4136 (
            .O(N__22621),
            .I(N__22615));
    Span4Mux_v I__4135 (
            .O(N__22618),
            .I(N__22610));
    Span4Mux_v I__4134 (
            .O(N__22615),
            .I(N__22610));
    Odrv4 I__4133 (
            .O(N__22610),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    InMux I__4132 (
            .O(N__22607),
            .I(N__22603));
    InMux I__4131 (
            .O(N__22606),
            .I(N__22600));
    LocalMux I__4130 (
            .O(N__22603),
            .I(N__22596));
    LocalMux I__4129 (
            .O(N__22600),
            .I(N__22593));
    InMux I__4128 (
            .O(N__22599),
            .I(N__22590));
    Span4Mux_v I__4127 (
            .O(N__22596),
            .I(N__22585));
    Span4Mux_v I__4126 (
            .O(N__22593),
            .I(N__22585));
    LocalMux I__4125 (
            .O(N__22590),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__4124 (
            .O(N__22585),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    CascadeMux I__4123 (
            .O(N__22580),
            .I(\ppm_encoder_1.N_302_cascade_ ));
    InMux I__4122 (
            .O(N__22577),
            .I(N__22571));
    InMux I__4121 (
            .O(N__22576),
            .I(N__22568));
    InMux I__4120 (
            .O(N__22575),
            .I(N__22565));
    InMux I__4119 (
            .O(N__22574),
            .I(N__22562));
    LocalMux I__4118 (
            .O(N__22571),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4117 (
            .O(N__22568),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4116 (
            .O(N__22565),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4115 (
            .O(N__22562),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__4114 (
            .O(N__22553),
            .I(N__22550));
    LocalMux I__4113 (
            .O(N__22550),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ));
    CascadeMux I__4112 (
            .O(N__22547),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ));
    InMux I__4111 (
            .O(N__22544),
            .I(N__22539));
    InMux I__4110 (
            .O(N__22543),
            .I(N__22534));
    InMux I__4109 (
            .O(N__22542),
            .I(N__22534));
    LocalMux I__4108 (
            .O(N__22539),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__4107 (
            .O(N__22534),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__4106 (
            .O(N__22529),
            .I(N__22524));
    CascadeMux I__4105 (
            .O(N__22528),
            .I(N__22521));
    InMux I__4104 (
            .O(N__22527),
            .I(N__22516));
    InMux I__4103 (
            .O(N__22524),
            .I(N__22516));
    InMux I__4102 (
            .O(N__22521),
            .I(N__22513));
    LocalMux I__4101 (
            .O(N__22516),
            .I(N__22510));
    LocalMux I__4100 (
            .O(N__22513),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    Odrv4 I__4099 (
            .O(N__22510),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__4098 (
            .O(N__22505),
            .I(N__22501));
    InMux I__4097 (
            .O(N__22504),
            .I(N__22497));
    InMux I__4096 (
            .O(N__22501),
            .I(N__22494));
    InMux I__4095 (
            .O(N__22500),
            .I(N__22491));
    LocalMux I__4094 (
            .O(N__22497),
            .I(N__22488));
    LocalMux I__4093 (
            .O(N__22494),
            .I(N__22485));
    LocalMux I__4092 (
            .O(N__22491),
            .I(N__22478));
    Sp12to4 I__4091 (
            .O(N__22488),
            .I(N__22473));
    Span12Mux_s4_h I__4090 (
            .O(N__22485),
            .I(N__22473));
    InMux I__4089 (
            .O(N__22484),
            .I(N__22468));
    InMux I__4088 (
            .O(N__22483),
            .I(N__22468));
    InMux I__4087 (
            .O(N__22482),
            .I(N__22465));
    InMux I__4086 (
            .O(N__22481),
            .I(N__22462));
    Odrv4 I__4085 (
            .O(N__22478),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv12 I__4084 (
            .O(N__22473),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__4083 (
            .O(N__22468),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__4082 (
            .O(N__22465),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__4081 (
            .O(N__22462),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__4080 (
            .O(N__22451),
            .I(N__22447));
    InMux I__4079 (
            .O(N__22450),
            .I(N__22443));
    InMux I__4078 (
            .O(N__22447),
            .I(N__22438));
    InMux I__4077 (
            .O(N__22446),
            .I(N__22438));
    LocalMux I__4076 (
            .O(N__22443),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__4075 (
            .O(N__22438),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__4074 (
            .O(N__22433),
            .I(N__22429));
    InMux I__4073 (
            .O(N__22432),
            .I(N__22426));
    LocalMux I__4072 (
            .O(N__22429),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    LocalMux I__4071 (
            .O(N__22426),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    InMux I__4070 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__4069 (
            .O(N__22418),
            .I(N__22414));
    InMux I__4068 (
            .O(N__22417),
            .I(N__22411));
    Span4Mux_h I__4067 (
            .O(N__22414),
            .I(N__22408));
    LocalMux I__4066 (
            .O(N__22411),
            .I(N__22402));
    Span4Mux_v I__4065 (
            .O(N__22408),
            .I(N__22398));
    InMux I__4064 (
            .O(N__22407),
            .I(N__22395));
    CascadeMux I__4063 (
            .O(N__22406),
            .I(N__22392));
    CascadeMux I__4062 (
            .O(N__22405),
            .I(N__22389));
    Span12Mux_s6_v I__4061 (
            .O(N__22402),
            .I(N__22386));
    InMux I__4060 (
            .O(N__22401),
            .I(N__22383));
    Span4Mux_v I__4059 (
            .O(N__22398),
            .I(N__22378));
    LocalMux I__4058 (
            .O(N__22395),
            .I(N__22378));
    InMux I__4057 (
            .O(N__22392),
            .I(N__22375));
    InMux I__4056 (
            .O(N__22389),
            .I(N__22372));
    Odrv12 I__4055 (
            .O(N__22386),
            .I(\ppm_encoder_1.N_227 ));
    LocalMux I__4054 (
            .O(N__22383),
            .I(\ppm_encoder_1.N_227 ));
    Odrv4 I__4053 (
            .O(N__22378),
            .I(\ppm_encoder_1.N_227 ));
    LocalMux I__4052 (
            .O(N__22375),
            .I(\ppm_encoder_1.N_227 ));
    LocalMux I__4051 (
            .O(N__22372),
            .I(\ppm_encoder_1.N_227 ));
    CascadeMux I__4050 (
            .O(N__22361),
            .I(N__22355));
    CascadeMux I__4049 (
            .O(N__22360),
            .I(N__22350));
    CascadeMux I__4048 (
            .O(N__22359),
            .I(N__22347));
    CascadeMux I__4047 (
            .O(N__22358),
            .I(N__22344));
    InMux I__4046 (
            .O(N__22355),
            .I(N__22338));
    InMux I__4045 (
            .O(N__22354),
            .I(N__22333));
    InMux I__4044 (
            .O(N__22353),
            .I(N__22333));
    InMux I__4043 (
            .O(N__22350),
            .I(N__22330));
    InMux I__4042 (
            .O(N__22347),
            .I(N__22327));
    InMux I__4041 (
            .O(N__22344),
            .I(N__22324));
    CascadeMux I__4040 (
            .O(N__22343),
            .I(N__22321));
    CascadeMux I__4039 (
            .O(N__22342),
            .I(N__22318));
    CascadeMux I__4038 (
            .O(N__22341),
            .I(N__22315));
    LocalMux I__4037 (
            .O(N__22338),
            .I(N__22311));
    LocalMux I__4036 (
            .O(N__22333),
            .I(N__22308));
    LocalMux I__4035 (
            .O(N__22330),
            .I(N__22305));
    LocalMux I__4034 (
            .O(N__22327),
            .I(N__22302));
    LocalMux I__4033 (
            .O(N__22324),
            .I(N__22299));
    InMux I__4032 (
            .O(N__22321),
            .I(N__22296));
    InMux I__4031 (
            .O(N__22318),
            .I(N__22291));
    InMux I__4030 (
            .O(N__22315),
            .I(N__22291));
    InMux I__4029 (
            .O(N__22314),
            .I(N__22288));
    Span4Mux_s2_h I__4028 (
            .O(N__22311),
            .I(N__22283));
    Span4Mux_v I__4027 (
            .O(N__22308),
            .I(N__22283));
    Span4Mux_s3_h I__4026 (
            .O(N__22305),
            .I(N__22280));
    Odrv4 I__4025 (
            .O(N__22302),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__4024 (
            .O(N__22299),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__4023 (
            .O(N__22296),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__4022 (
            .O(N__22291),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__4021 (
            .O(N__22288),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__4020 (
            .O(N__22283),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__4019 (
            .O(N__22280),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    CascadeMux I__4018 (
            .O(N__22265),
            .I(N__22257));
    CascadeMux I__4017 (
            .O(N__22264),
            .I(N__22253));
    InMux I__4016 (
            .O(N__22263),
            .I(N__22246));
    InMux I__4015 (
            .O(N__22262),
            .I(N__22243));
    InMux I__4014 (
            .O(N__22261),
            .I(N__22240));
    InMux I__4013 (
            .O(N__22260),
            .I(N__22237));
    InMux I__4012 (
            .O(N__22257),
            .I(N__22228));
    InMux I__4011 (
            .O(N__22256),
            .I(N__22228));
    InMux I__4010 (
            .O(N__22253),
            .I(N__22228));
    InMux I__4009 (
            .O(N__22252),
            .I(N__22228));
    InMux I__4008 (
            .O(N__22251),
            .I(N__22225));
    InMux I__4007 (
            .O(N__22250),
            .I(N__22219));
    InMux I__4006 (
            .O(N__22249),
            .I(N__22216));
    LocalMux I__4005 (
            .O(N__22246),
            .I(N__22209));
    LocalMux I__4004 (
            .O(N__22243),
            .I(N__22209));
    LocalMux I__4003 (
            .O(N__22240),
            .I(N__22209));
    LocalMux I__4002 (
            .O(N__22237),
            .I(N__22206));
    LocalMux I__4001 (
            .O(N__22228),
            .I(N__22203));
    LocalMux I__4000 (
            .O(N__22225),
            .I(N__22199));
    InMux I__3999 (
            .O(N__22224),
            .I(N__22194));
    InMux I__3998 (
            .O(N__22223),
            .I(N__22194));
    InMux I__3997 (
            .O(N__22222),
            .I(N__22191));
    LocalMux I__3996 (
            .O(N__22219),
            .I(N__22188));
    LocalMux I__3995 (
            .O(N__22216),
            .I(N__22179));
    Span4Mux_v I__3994 (
            .O(N__22209),
            .I(N__22179));
    Span4Mux_v I__3993 (
            .O(N__22206),
            .I(N__22179));
    Span4Mux_s2_h I__3992 (
            .O(N__22203),
            .I(N__22179));
    InMux I__3991 (
            .O(N__22202),
            .I(N__22176));
    Odrv4 I__3990 (
            .O(N__22199),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3989 (
            .O(N__22194),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3988 (
            .O(N__22191),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3987 (
            .O(N__22188),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3986 (
            .O(N__22179),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3985 (
            .O(N__22176),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    InMux I__3984 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__3983 (
            .O(N__22160),
            .I(N__22156));
    InMux I__3982 (
            .O(N__22159),
            .I(N__22153));
    Odrv4 I__3981 (
            .O(N__22156),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    LocalMux I__3980 (
            .O(N__22153),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    CascadeMux I__3979 (
            .O(N__22148),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ));
    CascadeMux I__3978 (
            .O(N__22145),
            .I(N__22142));
    InMux I__3977 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__3976 (
            .O(N__22139),
            .I(N__22136));
    Span4Mux_v I__3975 (
            .O(N__22136),
            .I(N__22133));
    Odrv4 I__3974 (
            .O(N__22133),
            .I(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ));
    CascadeMux I__3973 (
            .O(N__22130),
            .I(N__22126));
    InMux I__3972 (
            .O(N__22129),
            .I(N__22120));
    InMux I__3971 (
            .O(N__22126),
            .I(N__22117));
    CascadeMux I__3970 (
            .O(N__22125),
            .I(N__22114));
    CascadeMux I__3969 (
            .O(N__22124),
            .I(N__22111));
    CascadeMux I__3968 (
            .O(N__22123),
            .I(N__22107));
    LocalMux I__3967 (
            .O(N__22120),
            .I(N__22102));
    LocalMux I__3966 (
            .O(N__22117),
            .I(N__22099));
    InMux I__3965 (
            .O(N__22114),
            .I(N__22096));
    InMux I__3964 (
            .O(N__22111),
            .I(N__22092));
    CascadeMux I__3963 (
            .O(N__22110),
            .I(N__22089));
    InMux I__3962 (
            .O(N__22107),
            .I(N__22086));
    CascadeMux I__3961 (
            .O(N__22106),
            .I(N__22083));
    CascadeMux I__3960 (
            .O(N__22105),
            .I(N__22079));
    Span4Mux_s3_h I__3959 (
            .O(N__22102),
            .I(N__22075));
    Span4Mux_v I__3958 (
            .O(N__22099),
            .I(N__22070));
    LocalMux I__3957 (
            .O(N__22096),
            .I(N__22070));
    InMux I__3956 (
            .O(N__22095),
            .I(N__22067));
    LocalMux I__3955 (
            .O(N__22092),
            .I(N__22064));
    InMux I__3954 (
            .O(N__22089),
            .I(N__22061));
    LocalMux I__3953 (
            .O(N__22086),
            .I(N__22058));
    InMux I__3952 (
            .O(N__22083),
            .I(N__22055));
    InMux I__3951 (
            .O(N__22082),
            .I(N__22048));
    InMux I__3950 (
            .O(N__22079),
            .I(N__22048));
    InMux I__3949 (
            .O(N__22078),
            .I(N__22048));
    Odrv4 I__3948 (
            .O(N__22075),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__3947 (
            .O(N__22070),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3946 (
            .O(N__22067),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__3945 (
            .O(N__22064),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3944 (
            .O(N__22061),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__3943 (
            .O(N__22058),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3942 (
            .O(N__22055),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3941 (
            .O(N__22048),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    CascadeMux I__3940 (
            .O(N__22031),
            .I(N__22027));
    InMux I__3939 (
            .O(N__22030),
            .I(N__22023));
    InMux I__3938 (
            .O(N__22027),
            .I(N__22020));
    InMux I__3937 (
            .O(N__22026),
            .I(N__22017));
    LocalMux I__3936 (
            .O(N__22023),
            .I(N__22013));
    LocalMux I__3935 (
            .O(N__22020),
            .I(N__22010));
    LocalMux I__3934 (
            .O(N__22017),
            .I(N__22007));
    CascadeMux I__3933 (
            .O(N__22016),
            .I(N__22003));
    Span4Mux_s3_h I__3932 (
            .O(N__22013),
            .I(N__21993));
    Span4Mux_s3_h I__3931 (
            .O(N__22010),
            .I(N__21990));
    Span4Mux_s3_h I__3930 (
            .O(N__22007),
            .I(N__21987));
    InMux I__3929 (
            .O(N__22006),
            .I(N__21984));
    InMux I__3928 (
            .O(N__22003),
            .I(N__21979));
    InMux I__3927 (
            .O(N__22002),
            .I(N__21979));
    InMux I__3926 (
            .O(N__22001),
            .I(N__21976));
    InMux I__3925 (
            .O(N__22000),
            .I(N__21973));
    InMux I__3924 (
            .O(N__21999),
            .I(N__21970));
    InMux I__3923 (
            .O(N__21998),
            .I(N__21963));
    InMux I__3922 (
            .O(N__21997),
            .I(N__21963));
    InMux I__3921 (
            .O(N__21996),
            .I(N__21963));
    Odrv4 I__3920 (
            .O(N__21993),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__3919 (
            .O(N__21990),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__3918 (
            .O(N__21987),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3917 (
            .O(N__21984),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3916 (
            .O(N__21979),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3915 (
            .O(N__21976),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3914 (
            .O(N__21973),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3913 (
            .O(N__21970),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3912 (
            .O(N__21963),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__3911 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__3910 (
            .O(N__21941),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8 ));
    InMux I__3909 (
            .O(N__21938),
            .I(N__21929));
    InMux I__3908 (
            .O(N__21937),
            .I(N__21929));
    InMux I__3907 (
            .O(N__21936),
            .I(N__21929));
    LocalMux I__3906 (
            .O(N__21929),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    CascadeMux I__3905 (
            .O(N__21926),
            .I(N__21923));
    InMux I__3904 (
            .O(N__21923),
            .I(N__21919));
    InMux I__3903 (
            .O(N__21922),
            .I(N__21916));
    LocalMux I__3902 (
            .O(N__21919),
            .I(N__21913));
    LocalMux I__3901 (
            .O(N__21916),
            .I(N__21910));
    Span4Mux_h I__3900 (
            .O(N__21913),
            .I(N__21904));
    Span4Mux_s3_h I__3899 (
            .O(N__21910),
            .I(N__21904));
    InMux I__3898 (
            .O(N__21909),
            .I(N__21901));
    Span4Mux_v I__3897 (
            .O(N__21904),
            .I(N__21898));
    LocalMux I__3896 (
            .O(N__21901),
            .I(throttle_command_8));
    Odrv4 I__3895 (
            .O(N__21898),
            .I(throttle_command_8));
    InMux I__3894 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__3893 (
            .O(N__21890),
            .I(N__21887));
    Odrv4 I__3892 (
            .O(N__21887),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__3891 (
            .O(N__21884),
            .I(N__21875));
    InMux I__3890 (
            .O(N__21883),
            .I(N__21875));
    InMux I__3889 (
            .O(N__21882),
            .I(N__21875));
    LocalMux I__3888 (
            .O(N__21875),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__3887 (
            .O(N__21872),
            .I(N__21868));
    InMux I__3886 (
            .O(N__21871),
            .I(N__21865));
    LocalMux I__3885 (
            .O(N__21868),
            .I(N__21860));
    LocalMux I__3884 (
            .O(N__21865),
            .I(N__21860));
    Span4Mux_v I__3883 (
            .O(N__21860),
            .I(N__21857));
    Odrv4 I__3882 (
            .O(N__21857),
            .I(scaler_2_data_8));
    InMux I__3881 (
            .O(N__21854),
            .I(N__21851));
    LocalMux I__3880 (
            .O(N__21851),
            .I(N__21848));
    Odrv4 I__3879 (
            .O(N__21848),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__3878 (
            .O(N__21845),
            .I(N__21840));
    InMux I__3877 (
            .O(N__21844),
            .I(N__21837));
    InMux I__3876 (
            .O(N__21843),
            .I(N__21834));
    LocalMux I__3875 (
            .O(N__21840),
            .I(N__21829));
    LocalMux I__3874 (
            .O(N__21837),
            .I(N__21829));
    LocalMux I__3873 (
            .O(N__21834),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__3872 (
            .O(N__21829),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__3871 (
            .O(N__21824),
            .I(N__21821));
    LocalMux I__3870 (
            .O(N__21821),
            .I(N__21818));
    Odrv4 I__3869 (
            .O(N__21818),
            .I(\ppm_encoder_1.N_296 ));
    InMux I__3868 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__3867 (
            .O(N__21812),
            .I(N__21808));
    InMux I__3866 (
            .O(N__21811),
            .I(N__21805));
    Odrv12 I__3865 (
            .O(N__21808),
            .I(throttle_command_4));
    LocalMux I__3864 (
            .O(N__21805),
            .I(throttle_command_4));
    InMux I__3863 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__3862 (
            .O(N__21797),
            .I(N__21794));
    Span4Mux_h I__3861 (
            .O(N__21794),
            .I(N__21791));
    Odrv4 I__3860 (
            .O(N__21791),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__3859 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__3858 (
            .O(N__21785),
            .I(N__21782));
    Span4Mux_h I__3857 (
            .O(N__21782),
            .I(N__21778));
    InMux I__3856 (
            .O(N__21781),
            .I(N__21775));
    Odrv4 I__3855 (
            .O(N__21778),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    LocalMux I__3854 (
            .O(N__21775),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    CascadeMux I__3853 (
            .O(N__21770),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    CascadeMux I__3852 (
            .O(N__21767),
            .I(N__21764));
    InMux I__3851 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__3850 (
            .O(N__21761),
            .I(N__21758));
    Span4Mux_v I__3849 (
            .O(N__21758),
            .I(N__21755));
    Odrv4 I__3848 (
            .O(N__21755),
            .I(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ));
    InMux I__3847 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__3846 (
            .O(N__21749),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    CascadeMux I__3845 (
            .O(N__21746),
            .I(\ppm_encoder_1.N_304_cascade_ ));
    CascadeMux I__3844 (
            .O(N__21743),
            .I(N__21739));
    InMux I__3843 (
            .O(N__21742),
            .I(N__21736));
    InMux I__3842 (
            .O(N__21739),
            .I(N__21733));
    LocalMux I__3841 (
            .O(N__21736),
            .I(N__21730));
    LocalMux I__3840 (
            .O(N__21733),
            .I(N__21727));
    Span4Mux_v I__3839 (
            .O(N__21730),
            .I(N__21724));
    Odrv12 I__3838 (
            .O(N__21727),
            .I(scaler_2_data_12));
    Odrv4 I__3837 (
            .O(N__21724),
            .I(scaler_2_data_12));
    InMux I__3836 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__3835 (
            .O(N__21716),
            .I(N__21713));
    Odrv4 I__3834 (
            .O(N__21713),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__3833 (
            .O(N__21710),
            .I(N__21701));
    InMux I__3832 (
            .O(N__21709),
            .I(N__21701));
    InMux I__3831 (
            .O(N__21708),
            .I(N__21701));
    LocalMux I__3830 (
            .O(N__21701),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__3829 (
            .O(N__21698),
            .I(N__21689));
    InMux I__3828 (
            .O(N__21697),
            .I(N__21689));
    InMux I__3827 (
            .O(N__21696),
            .I(N__21689));
    LocalMux I__3826 (
            .O(N__21689),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__3825 (
            .O(N__21686),
            .I(N__21682));
    InMux I__3824 (
            .O(N__21685),
            .I(N__21679));
    LocalMux I__3823 (
            .O(N__21682),
            .I(N__21676));
    LocalMux I__3822 (
            .O(N__21679),
            .I(N__21673));
    Span4Mux_h I__3821 (
            .O(N__21676),
            .I(N__21670));
    Span4Mux_s2_h I__3820 (
            .O(N__21673),
            .I(N__21667));
    Odrv4 I__3819 (
            .O(N__21670),
            .I(throttle_command_12));
    Odrv4 I__3818 (
            .O(N__21667),
            .I(throttle_command_12));
    InMux I__3817 (
            .O(N__21662),
            .I(N__21659));
    LocalMux I__3816 (
            .O(N__21659),
            .I(N__21656));
    Span4Mux_h I__3815 (
            .O(N__21656),
            .I(N__21653));
    Odrv4 I__3814 (
            .O(N__21653),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__3813 (
            .O(N__21650),
            .I(N__21641));
    InMux I__3812 (
            .O(N__21649),
            .I(N__21641));
    InMux I__3811 (
            .O(N__21648),
            .I(N__21641));
    LocalMux I__3810 (
            .O(N__21641),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    InMux I__3809 (
            .O(N__21638),
            .I(N__21614));
    InMux I__3808 (
            .O(N__21637),
            .I(N__21614));
    InMux I__3807 (
            .O(N__21636),
            .I(N__21614));
    InMux I__3806 (
            .O(N__21635),
            .I(N__21614));
    InMux I__3805 (
            .O(N__21634),
            .I(N__21611));
    InMux I__3804 (
            .O(N__21633),
            .I(N__21608));
    InMux I__3803 (
            .O(N__21632),
            .I(N__21605));
    InMux I__3802 (
            .O(N__21631),
            .I(N__21592));
    InMux I__3801 (
            .O(N__21630),
            .I(N__21592));
    InMux I__3800 (
            .O(N__21629),
            .I(N__21592));
    InMux I__3799 (
            .O(N__21628),
            .I(N__21592));
    InMux I__3798 (
            .O(N__21627),
            .I(N__21592));
    InMux I__3797 (
            .O(N__21626),
            .I(N__21592));
    InMux I__3796 (
            .O(N__21625),
            .I(N__21589));
    InMux I__3795 (
            .O(N__21624),
            .I(N__21586));
    InMux I__3794 (
            .O(N__21623),
            .I(N__21583));
    LocalMux I__3793 (
            .O(N__21614),
            .I(N__21566));
    LocalMux I__3792 (
            .O(N__21611),
            .I(N__21563));
    LocalMux I__3791 (
            .O(N__21608),
            .I(N__21560));
    LocalMux I__3790 (
            .O(N__21605),
            .I(N__21557));
    LocalMux I__3789 (
            .O(N__21592),
            .I(N__21554));
    LocalMux I__3788 (
            .O(N__21589),
            .I(N__21551));
    LocalMux I__3787 (
            .O(N__21586),
            .I(N__21548));
    LocalMux I__3786 (
            .O(N__21583),
            .I(N__21545));
    SRMux I__3785 (
            .O(N__21582),
            .I(N__21500));
    SRMux I__3784 (
            .O(N__21581),
            .I(N__21500));
    SRMux I__3783 (
            .O(N__21580),
            .I(N__21500));
    SRMux I__3782 (
            .O(N__21579),
            .I(N__21500));
    SRMux I__3781 (
            .O(N__21578),
            .I(N__21500));
    SRMux I__3780 (
            .O(N__21577),
            .I(N__21500));
    SRMux I__3779 (
            .O(N__21576),
            .I(N__21500));
    SRMux I__3778 (
            .O(N__21575),
            .I(N__21500));
    SRMux I__3777 (
            .O(N__21574),
            .I(N__21500));
    SRMux I__3776 (
            .O(N__21573),
            .I(N__21500));
    SRMux I__3775 (
            .O(N__21572),
            .I(N__21500));
    SRMux I__3774 (
            .O(N__21571),
            .I(N__21500));
    SRMux I__3773 (
            .O(N__21570),
            .I(N__21500));
    SRMux I__3772 (
            .O(N__21569),
            .I(N__21500));
    Glb2LocalMux I__3771 (
            .O(N__21566),
            .I(N__21500));
    Glb2LocalMux I__3770 (
            .O(N__21563),
            .I(N__21500));
    Glb2LocalMux I__3769 (
            .O(N__21560),
            .I(N__21500));
    Glb2LocalMux I__3768 (
            .O(N__21557),
            .I(N__21500));
    Glb2LocalMux I__3767 (
            .O(N__21554),
            .I(N__21500));
    Glb2LocalMux I__3766 (
            .O(N__21551),
            .I(N__21500));
    Glb2LocalMux I__3765 (
            .O(N__21548),
            .I(N__21500));
    Glb2LocalMux I__3764 (
            .O(N__21545),
            .I(N__21500));
    GlobalMux I__3763 (
            .O(N__21500),
            .I(N__21497));
    gio2CtrlBuf I__3762 (
            .O(N__21497),
            .I(N_423_g));
    IoInMux I__3761 (
            .O(N__21494),
            .I(N__21491));
    LocalMux I__3760 (
            .O(N__21491),
            .I(N__21488));
    Span12Mux_s11_v I__3759 (
            .O(N__21488),
            .I(N__21485));
    Odrv12 I__3758 (
            .O(N__21485),
            .I(\pid_alt.N_422_0 ));
    CEMux I__3757 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__3756 (
            .O(N__21479),
            .I(\pid_alt.state_1_0_0 ));
    InMux I__3755 (
            .O(N__21476),
            .I(N__21472));
    InMux I__3754 (
            .O(N__21475),
            .I(N__21469));
    LocalMux I__3753 (
            .O(N__21472),
            .I(N__21465));
    LocalMux I__3752 (
            .O(N__21469),
            .I(N__21462));
    InMux I__3751 (
            .O(N__21468),
            .I(N__21459));
    Span12Mux_s4_h I__3750 (
            .O(N__21465),
            .I(N__21456));
    Span4Mux_h I__3749 (
            .O(N__21462),
            .I(N__21453));
    LocalMux I__3748 (
            .O(N__21459),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv12 I__3747 (
            .O(N__21456),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__3746 (
            .O(N__21453),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__3745 (
            .O(N__21446),
            .I(N__21442));
    CascadeMux I__3744 (
            .O(N__21445),
            .I(N__21439));
    LocalMux I__3743 (
            .O(N__21442),
            .I(N__21436));
    InMux I__3742 (
            .O(N__21439),
            .I(N__21433));
    Span4Mux_v I__3741 (
            .O(N__21436),
            .I(N__21427));
    LocalMux I__3740 (
            .O(N__21433),
            .I(N__21427));
    InMux I__3739 (
            .O(N__21432),
            .I(N__21424));
    Span4Mux_v I__3738 (
            .O(N__21427),
            .I(N__21421));
    LocalMux I__3737 (
            .O(N__21424),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__3736 (
            .O(N__21421),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    InMux I__3735 (
            .O(N__21416),
            .I(N__21412));
    CascadeMux I__3734 (
            .O(N__21415),
            .I(N__21408));
    LocalMux I__3733 (
            .O(N__21412),
            .I(N__21405));
    InMux I__3732 (
            .O(N__21411),
            .I(N__21402));
    InMux I__3731 (
            .O(N__21408),
            .I(N__21399));
    Span4Mux_v I__3730 (
            .O(N__21405),
            .I(N__21396));
    LocalMux I__3729 (
            .O(N__21402),
            .I(N__21393));
    LocalMux I__3728 (
            .O(N__21399),
            .I(throttle_command_10));
    Odrv4 I__3727 (
            .O(N__21396),
            .I(throttle_command_10));
    Odrv12 I__3726 (
            .O(N__21393),
            .I(throttle_command_10));
    CascadeMux I__3725 (
            .O(N__21386),
            .I(N__21383));
    InMux I__3724 (
            .O(N__21383),
            .I(N__21380));
    LocalMux I__3723 (
            .O(N__21380),
            .I(N__21377));
    Span4Mux_v I__3722 (
            .O(N__21377),
            .I(N__21374));
    Odrv4 I__3721 (
            .O(N__21374),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__3720 (
            .O(N__21371),
            .I(N__21367));
    InMux I__3719 (
            .O(N__21370),
            .I(N__21364));
    LocalMux I__3718 (
            .O(N__21367),
            .I(N__21361));
    LocalMux I__3717 (
            .O(N__21364),
            .I(N__21358));
    Span4Mux_v I__3716 (
            .O(N__21361),
            .I(N__21353));
    Span4Mux_v I__3715 (
            .O(N__21358),
            .I(N__21353));
    Odrv4 I__3714 (
            .O(N__21353),
            .I(throttle_command_13));
    InMux I__3713 (
            .O(N__21350),
            .I(N__21347));
    LocalMux I__3712 (
            .O(N__21347),
            .I(N__21344));
    Span4Mux_h I__3711 (
            .O(N__21344),
            .I(N__21341));
    Odrv4 I__3710 (
            .O(N__21341),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__3709 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__3708 (
            .O(N__21335),
            .I(N__21332));
    Span4Mux_h I__3707 (
            .O(N__21332),
            .I(N__21329));
    Odrv4 I__3706 (
            .O(N__21329),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    CascadeMux I__3705 (
            .O(N__21326),
            .I(N__21323));
    InMux I__3704 (
            .O(N__21323),
            .I(N__21319));
    InMux I__3703 (
            .O(N__21322),
            .I(N__21316));
    LocalMux I__3702 (
            .O(N__21319),
            .I(N__21313));
    LocalMux I__3701 (
            .O(N__21316),
            .I(N__21310));
    Span4Mux_v I__3700 (
            .O(N__21313),
            .I(N__21307));
    Span4Mux_s3_h I__3699 (
            .O(N__21310),
            .I(N__21304));
    Odrv4 I__3698 (
            .O(N__21307),
            .I(throttle_command_2));
    Odrv4 I__3697 (
            .O(N__21304),
            .I(throttle_command_2));
    CascadeMux I__3696 (
            .O(N__21299),
            .I(N__21296));
    InMux I__3695 (
            .O(N__21296),
            .I(N__21290));
    InMux I__3694 (
            .O(N__21295),
            .I(N__21290));
    LocalMux I__3693 (
            .O(N__21290),
            .I(N__21287));
    Span4Mux_h I__3692 (
            .O(N__21287),
            .I(N__21284));
    Odrv4 I__3691 (
            .O(N__21284),
            .I(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ));
    InMux I__3690 (
            .O(N__21281),
            .I(\scaler_2.un2_source_data_0_cry_5 ));
    CascadeMux I__3689 (
            .O(N__21278),
            .I(N__21275));
    InMux I__3688 (
            .O(N__21275),
            .I(N__21269));
    InMux I__3687 (
            .O(N__21274),
            .I(N__21269));
    LocalMux I__3686 (
            .O(N__21269),
            .I(N__21266));
    Span4Mux_h I__3685 (
            .O(N__21266),
            .I(N__21263));
    Odrv4 I__3684 (
            .O(N__21263),
            .I(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ));
    CascadeMux I__3683 (
            .O(N__21260),
            .I(N__21257));
    InMux I__3682 (
            .O(N__21257),
            .I(N__21253));
    InMux I__3681 (
            .O(N__21256),
            .I(N__21250));
    LocalMux I__3680 (
            .O(N__21253),
            .I(N__21247));
    LocalMux I__3679 (
            .O(N__21250),
            .I(N__21244));
    Span12Mux_s4_h I__3678 (
            .O(N__21247),
            .I(N__21241));
    Span4Mux_v I__3677 (
            .O(N__21244),
            .I(N__21238));
    Odrv12 I__3676 (
            .O(N__21241),
            .I(scaler_2_data_11));
    Odrv4 I__3675 (
            .O(N__21238),
            .I(scaler_2_data_11));
    InMux I__3674 (
            .O(N__21233),
            .I(\scaler_2.un2_source_data_0_cry_6 ));
    CascadeMux I__3673 (
            .O(N__21230),
            .I(N__21227));
    InMux I__3672 (
            .O(N__21227),
            .I(N__21221));
    InMux I__3671 (
            .O(N__21226),
            .I(N__21221));
    LocalMux I__3670 (
            .O(N__21221),
            .I(N__21218));
    Span4Mux_h I__3669 (
            .O(N__21218),
            .I(N__21215));
    Odrv4 I__3668 (
            .O(N__21215),
            .I(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ));
    InMux I__3667 (
            .O(N__21212),
            .I(\scaler_2.un2_source_data_0_cry_7 ));
    InMux I__3666 (
            .O(N__21209),
            .I(N__21205));
    InMux I__3665 (
            .O(N__21208),
            .I(N__21202));
    LocalMux I__3664 (
            .O(N__21205),
            .I(N__21199));
    LocalMux I__3663 (
            .O(N__21202),
            .I(N__21196));
    Span4Mux_h I__3662 (
            .O(N__21199),
            .I(N__21193));
    Span4Mux_h I__3661 (
            .O(N__21196),
            .I(N__21190));
    Odrv4 I__3660 (
            .O(N__21193),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    Odrv4 I__3659 (
            .O(N__21190),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    CascadeMux I__3658 (
            .O(N__21185),
            .I(N__21182));
    InMux I__3657 (
            .O(N__21182),
            .I(N__21179));
    LocalMux I__3656 (
            .O(N__21179),
            .I(N__21176));
    Span4Mux_h I__3655 (
            .O(N__21176),
            .I(N__21173));
    Odrv4 I__3654 (
            .O(N__21173),
            .I(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ));
    InMux I__3653 (
            .O(N__21170),
            .I(bfn_4_17_0_));
    InMux I__3652 (
            .O(N__21167),
            .I(\scaler_2.un2_source_data_0_cry_9 ));
    InMux I__3651 (
            .O(N__21164),
            .I(N__21161));
    LocalMux I__3650 (
            .O(N__21161),
            .I(N__21158));
    Span4Mux_h I__3649 (
            .O(N__21158),
            .I(N__21155));
    Span4Mux_v I__3648 (
            .O(N__21155),
            .I(N__21152));
    Odrv4 I__3647 (
            .O(N__21152),
            .I(scaler_2_data_14));
    InMux I__3646 (
            .O(N__21149),
            .I(N__21146));
    LocalMux I__3645 (
            .O(N__21146),
            .I(N__21143));
    Span12Mux_v I__3644 (
            .O(N__21143),
            .I(N__21140));
    Odrv12 I__3643 (
            .O(N__21140),
            .I(alt_ki_7));
    InMux I__3642 (
            .O(N__21137),
            .I(N__21134));
    LocalMux I__3641 (
            .O(N__21134),
            .I(N__21131));
    Span4Mux_h I__3640 (
            .O(N__21131),
            .I(N__21127));
    InMux I__3639 (
            .O(N__21130),
            .I(N__21124));
    Odrv4 I__3638 (
            .O(N__21127),
            .I(\pid_alt.un1_pid_prereg_0_axb_1 ));
    LocalMux I__3637 (
            .O(N__21124),
            .I(\pid_alt.un1_pid_prereg_0_axb_1 ));
    CascadeMux I__3636 (
            .O(N__21119),
            .I(N__21116));
    InMux I__3635 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__3634 (
            .O(N__21113),
            .I(N__21110));
    Span4Mux_v I__3633 (
            .O(N__21110),
            .I(N__21107));
    Odrv4 I__3632 (
            .O(N__21107),
            .I(\pid_alt.un1_pid_prereg_0_cry_0_THRU_CO ));
    InMux I__3631 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__3630 (
            .O(N__21101),
            .I(N__21098));
    Span4Mux_h I__3629 (
            .O(N__21098),
            .I(N__21093));
    InMux I__3628 (
            .O(N__21097),
            .I(N__21090));
    InMux I__3627 (
            .O(N__21096),
            .I(N__21087));
    Odrv4 I__3626 (
            .O(N__21093),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    LocalMux I__3625 (
            .O(N__21090),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    LocalMux I__3624 (
            .O(N__21087),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__3623 (
            .O(N__21080),
            .I(N__21077));
    LocalMux I__3622 (
            .O(N__21077),
            .I(N__21074));
    Odrv4 I__3621 (
            .O(N__21074),
            .I(\scaler_2.N_881_i_l_ofxZ0 ));
    InMux I__3620 (
            .O(N__21071),
            .I(N__21065));
    InMux I__3619 (
            .O(N__21070),
            .I(N__21065));
    LocalMux I__3618 (
            .O(N__21065),
            .I(frame_decoder_CH2data_7));
    InMux I__3617 (
            .O(N__21062),
            .I(N__21059));
    LocalMux I__3616 (
            .O(N__21059),
            .I(N__21056));
    Span4Mux_h I__3615 (
            .O(N__21056),
            .I(N__21053));
    Odrv4 I__3614 (
            .O(N__21053),
            .I(\scaler_2.un3_source_data_0_axb_7 ));
    InMux I__3613 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__3612 (
            .O(N__21047),
            .I(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ));
    CascadeMux I__3611 (
            .O(N__21044),
            .I(N__21038));
    CascadeMux I__3610 (
            .O(N__21043),
            .I(N__21035));
    InMux I__3609 (
            .O(N__21042),
            .I(N__21032));
    InMux I__3608 (
            .O(N__21041),
            .I(N__21029));
    InMux I__3607 (
            .O(N__21038),
            .I(N__21026));
    InMux I__3606 (
            .O(N__21035),
            .I(N__21023));
    LocalMux I__3605 (
            .O(N__21032),
            .I(N__21020));
    LocalMux I__3604 (
            .O(N__21029),
            .I(N__21017));
    LocalMux I__3603 (
            .O(N__21026),
            .I(N__21012));
    LocalMux I__3602 (
            .O(N__21023),
            .I(N__21012));
    Span4Mux_v I__3601 (
            .O(N__21020),
            .I(N__21009));
    Span4Mux_v I__3600 (
            .O(N__21017),
            .I(N__21004));
    Span4Mux_h I__3599 (
            .O(N__21012),
            .I(N__21004));
    Odrv4 I__3598 (
            .O(N__21009),
            .I(\scaler_2.un2_source_data_0 ));
    Odrv4 I__3597 (
            .O(N__21004),
            .I(\scaler_2.un2_source_data_0 ));
    InMux I__3596 (
            .O(N__20999),
            .I(\scaler_2.un2_source_data_0_cry_1 ));
    CascadeMux I__3595 (
            .O(N__20996),
            .I(N__20993));
    InMux I__3594 (
            .O(N__20993),
            .I(N__20987));
    InMux I__3593 (
            .O(N__20992),
            .I(N__20987));
    LocalMux I__3592 (
            .O(N__20987),
            .I(N__20984));
    Span4Mux_v I__3591 (
            .O(N__20984),
            .I(N__20981));
    Odrv4 I__3590 (
            .O(N__20981),
            .I(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ));
    InMux I__3589 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__3588 (
            .O(N__20975),
            .I(N__20971));
    InMux I__3587 (
            .O(N__20974),
            .I(N__20968));
    Span4Mux_h I__3586 (
            .O(N__20971),
            .I(N__20963));
    LocalMux I__3585 (
            .O(N__20968),
            .I(N__20963));
    Span4Mux_v I__3584 (
            .O(N__20963),
            .I(N__20960));
    Odrv4 I__3583 (
            .O(N__20960),
            .I(scaler_2_data_7));
    InMux I__3582 (
            .O(N__20957),
            .I(\scaler_2.un2_source_data_0_cry_2 ));
    CascadeMux I__3581 (
            .O(N__20954),
            .I(N__20951));
    InMux I__3580 (
            .O(N__20951),
            .I(N__20945));
    InMux I__3579 (
            .O(N__20950),
            .I(N__20945));
    LocalMux I__3578 (
            .O(N__20945),
            .I(N__20942));
    Span4Mux_v I__3577 (
            .O(N__20942),
            .I(N__20939));
    Odrv4 I__3576 (
            .O(N__20939),
            .I(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ));
    InMux I__3575 (
            .O(N__20936),
            .I(\scaler_2.un2_source_data_0_cry_3 ));
    CascadeMux I__3574 (
            .O(N__20933),
            .I(N__20930));
    InMux I__3573 (
            .O(N__20930),
            .I(N__20924));
    InMux I__3572 (
            .O(N__20929),
            .I(N__20924));
    LocalMux I__3571 (
            .O(N__20924),
            .I(N__20921));
    Span4Mux_v I__3570 (
            .O(N__20921),
            .I(N__20918));
    Odrv4 I__3569 (
            .O(N__20918),
            .I(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ));
    InMux I__3568 (
            .O(N__20915),
            .I(N__20912));
    LocalMux I__3567 (
            .O(N__20912),
            .I(N__20909));
    Span4Mux_v I__3566 (
            .O(N__20909),
            .I(N__20905));
    InMux I__3565 (
            .O(N__20908),
            .I(N__20902));
    Span4Mux_h I__3564 (
            .O(N__20905),
            .I(N__20899));
    LocalMux I__3563 (
            .O(N__20902),
            .I(N__20896));
    Span4Mux_v I__3562 (
            .O(N__20899),
            .I(N__20893));
    Span4Mux_v I__3561 (
            .O(N__20896),
            .I(N__20890));
    Odrv4 I__3560 (
            .O(N__20893),
            .I(scaler_2_data_9));
    Odrv4 I__3559 (
            .O(N__20890),
            .I(scaler_2_data_9));
    InMux I__3558 (
            .O(N__20885),
            .I(\scaler_2.un2_source_data_0_cry_4 ));
    InMux I__3557 (
            .O(N__20882),
            .I(N__20878));
    CascadeMux I__3556 (
            .O(N__20881),
            .I(N__20875));
    LocalMux I__3555 (
            .O(N__20878),
            .I(N__20870));
    InMux I__3554 (
            .O(N__20875),
            .I(N__20867));
    InMux I__3553 (
            .O(N__20874),
            .I(N__20862));
    InMux I__3552 (
            .O(N__20873),
            .I(N__20862));
    Span4Mux_v I__3551 (
            .O(N__20870),
            .I(N__20856));
    LocalMux I__3550 (
            .O(N__20867),
            .I(N__20856));
    LocalMux I__3549 (
            .O(N__20862),
            .I(N__20853));
    InMux I__3548 (
            .O(N__20861),
            .I(N__20850));
    Span4Mux_v I__3547 (
            .O(N__20856),
            .I(N__20847));
    Span4Mux_h I__3546 (
            .O(N__20853),
            .I(N__20841));
    LocalMux I__3545 (
            .O(N__20850),
            .I(N__20838));
    Sp12to4 I__3544 (
            .O(N__20847),
            .I(N__20835));
    InMux I__3543 (
            .O(N__20846),
            .I(N__20828));
    InMux I__3542 (
            .O(N__20845),
            .I(N__20828));
    InMux I__3541 (
            .O(N__20844),
            .I(N__20828));
    Span4Mux_v I__3540 (
            .O(N__20841),
            .I(N__20825));
    Span4Mux_h I__3539 (
            .O(N__20838),
            .I(N__20822));
    Span12Mux_s1_h I__3538 (
            .O(N__20835),
            .I(N__20817));
    LocalMux I__3537 (
            .O(N__20828),
            .I(N__20817));
    Odrv4 I__3536 (
            .O(N__20825),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    Odrv4 I__3535 (
            .O(N__20822),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    Odrv12 I__3534 (
            .O(N__20817),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__3533 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__3532 (
            .O(N__20807),
            .I(N__20804));
    Span4Mux_v I__3531 (
            .O(N__20804),
            .I(N__20800));
    InMux I__3530 (
            .O(N__20803),
            .I(N__20796));
    Span4Mux_h I__3529 (
            .O(N__20800),
            .I(N__20793));
    CascadeMux I__3528 (
            .O(N__20799),
            .I(N__20790));
    LocalMux I__3527 (
            .O(N__20796),
            .I(N__20785));
    Sp12to4 I__3526 (
            .O(N__20793),
            .I(N__20782));
    InMux I__3525 (
            .O(N__20790),
            .I(N__20775));
    InMux I__3524 (
            .O(N__20789),
            .I(N__20775));
    InMux I__3523 (
            .O(N__20788),
            .I(N__20775));
    Span4Mux_v I__3522 (
            .O(N__20785),
            .I(N__20772));
    Span12Mux_h I__3521 (
            .O(N__20782),
            .I(N__20767));
    LocalMux I__3520 (
            .O(N__20775),
            .I(N__20767));
    Span4Mux_h I__3519 (
            .O(N__20772),
            .I(N__20764));
    Span12Mux_v I__3518 (
            .O(N__20767),
            .I(N__20761));
    Odrv4 I__3517 (
            .O(N__20764),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    Odrv12 I__3516 (
            .O(N__20761),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    CascadeMux I__3515 (
            .O(N__20756),
            .I(N__20753));
    InMux I__3514 (
            .O(N__20753),
            .I(N__20750));
    LocalMux I__3513 (
            .O(N__20750),
            .I(N__20747));
    Span4Mux_h I__3512 (
            .O(N__20747),
            .I(N__20744));
    Sp12to4 I__3511 (
            .O(N__20744),
            .I(N__20741));
    Odrv12 I__3510 (
            .O(N__20741),
            .I(\pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20 ));
    InMux I__3509 (
            .O(N__20738),
            .I(N__20735));
    LocalMux I__3508 (
            .O(N__20735),
            .I(N__20732));
    Odrv4 I__3507 (
            .O(N__20732),
            .I(frame_decoder_CH2data_1));
    InMux I__3506 (
            .O(N__20729),
            .I(N__20726));
    LocalMux I__3505 (
            .O(N__20726),
            .I(N__20723));
    Odrv4 I__3504 (
            .O(N__20723),
            .I(frame_decoder_CH2data_2));
    InMux I__3503 (
            .O(N__20720),
            .I(N__20717));
    LocalMux I__3502 (
            .O(N__20717),
            .I(N__20714));
    Odrv4 I__3501 (
            .O(N__20714),
            .I(frame_decoder_CH2data_3));
    CascadeMux I__3500 (
            .O(N__20711),
            .I(N__20708));
    InMux I__3499 (
            .O(N__20708),
            .I(N__20705));
    LocalMux I__3498 (
            .O(N__20705),
            .I(N__20702));
    Odrv4 I__3497 (
            .O(N__20702),
            .I(frame_decoder_CH2data_4));
    CascadeMux I__3496 (
            .O(N__20699),
            .I(N__20696));
    InMux I__3495 (
            .O(N__20696),
            .I(N__20693));
    LocalMux I__3494 (
            .O(N__20693),
            .I(N__20690));
    Odrv4 I__3493 (
            .O(N__20690),
            .I(frame_decoder_CH2data_5));
    CascadeMux I__3492 (
            .O(N__20687),
            .I(N__20684));
    InMux I__3491 (
            .O(N__20684),
            .I(N__20681));
    LocalMux I__3490 (
            .O(N__20681),
            .I(N__20678));
    Odrv4 I__3489 (
            .O(N__20678),
            .I(frame_decoder_CH2data_6));
    InMux I__3488 (
            .O(N__20675),
            .I(N__20672));
    LocalMux I__3487 (
            .O(N__20672),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    InMux I__3486 (
            .O(N__20669),
            .I(N__20666));
    LocalMux I__3485 (
            .O(N__20666),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    InMux I__3484 (
            .O(N__20663),
            .I(N__20660));
    LocalMux I__3483 (
            .O(N__20660),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__3482 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__3481 (
            .O(N__20654),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__3480 (
            .O(N__20651),
            .I(N__20648));
    LocalMux I__3479 (
            .O(N__20648),
            .I(drone_altitude_14));
    InMux I__3478 (
            .O(N__20645),
            .I(N__20642));
    LocalMux I__3477 (
            .O(N__20642),
            .I(drone_altitude_2));
    InMux I__3476 (
            .O(N__20639),
            .I(N__20636));
    LocalMux I__3475 (
            .O(N__20636),
            .I(drone_altitude_3));
    CascadeMux I__3474 (
            .O(N__20633),
            .I(N__20630));
    InMux I__3473 (
            .O(N__20630),
            .I(N__20626));
    InMux I__3472 (
            .O(N__20629),
            .I(N__20623));
    LocalMux I__3471 (
            .O(N__20626),
            .I(N__20615));
    LocalMux I__3470 (
            .O(N__20623),
            .I(N__20615));
    InMux I__3469 (
            .O(N__20622),
            .I(N__20612));
    InMux I__3468 (
            .O(N__20621),
            .I(N__20607));
    InMux I__3467 (
            .O(N__20620),
            .I(N__20607));
    Span4Mux_v I__3466 (
            .O(N__20615),
            .I(N__20604));
    LocalMux I__3465 (
            .O(N__20612),
            .I(N__20601));
    LocalMux I__3464 (
            .O(N__20607),
            .I(N__20598));
    Span4Mux_v I__3463 (
            .O(N__20604),
            .I(N__20595));
    Span4Mux_h I__3462 (
            .O(N__20601),
            .I(N__20590));
    Span4Mux_v I__3461 (
            .O(N__20598),
            .I(N__20590));
    Odrv4 I__3460 (
            .O(N__20595),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    Odrv4 I__3459 (
            .O(N__20590),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    CascadeMux I__3458 (
            .O(N__20585),
            .I(N__20582));
    InMux I__3457 (
            .O(N__20582),
            .I(N__20576));
    InMux I__3456 (
            .O(N__20581),
            .I(N__20576));
    LocalMux I__3455 (
            .O(N__20576),
            .I(N__20573));
    Span4Mux_h I__3454 (
            .O(N__20573),
            .I(N__20569));
    InMux I__3453 (
            .O(N__20572),
            .I(N__20566));
    Span4Mux_v I__3452 (
            .O(N__20569),
            .I(N__20561));
    LocalMux I__3451 (
            .O(N__20566),
            .I(N__20561));
    Span4Mux_v I__3450 (
            .O(N__20561),
            .I(N__20558));
    Span4Mux_v I__3449 (
            .O(N__20558),
            .I(N__20555));
    Odrv4 I__3448 (
            .O(N__20555),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__3447 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__3446 (
            .O(N__20549),
            .I(N__20546));
    Span4Mux_h I__3445 (
            .O(N__20546),
            .I(N__20543));
    Span4Mux_v I__3444 (
            .O(N__20543),
            .I(N__20540));
    Odrv4 I__3443 (
            .O(N__20540),
            .I(\pid_alt.error_p_reg_esr_RNIF43KZ0Z_18 ));
    CascadeMux I__3442 (
            .O(N__20537),
            .I(N__20534));
    InMux I__3441 (
            .O(N__20534),
            .I(N__20530));
    InMux I__3440 (
            .O(N__20533),
            .I(N__20525));
    LocalMux I__3439 (
            .O(N__20530),
            .I(N__20522));
    InMux I__3438 (
            .O(N__20529),
            .I(N__20519));
    InMux I__3437 (
            .O(N__20528),
            .I(N__20516));
    LocalMux I__3436 (
            .O(N__20525),
            .I(N__20513));
    Span4Mux_s1_v I__3435 (
            .O(N__20522),
            .I(N__20508));
    LocalMux I__3434 (
            .O(N__20519),
            .I(N__20508));
    LocalMux I__3433 (
            .O(N__20516),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__3432 (
            .O(N__20513),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__3431 (
            .O(N__20508),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    InMux I__3430 (
            .O(N__20501),
            .I(N__20498));
    LocalMux I__3429 (
            .O(N__20498),
            .I(N__20495));
    Span4Mux_h I__3428 (
            .O(N__20495),
            .I(N__20492));
    Odrv4 I__3427 (
            .O(N__20492),
            .I(alt_kp_7));
    InMux I__3426 (
            .O(N__20489),
            .I(N__20486));
    LocalMux I__3425 (
            .O(N__20486),
            .I(N__20482));
    InMux I__3424 (
            .O(N__20485),
            .I(N__20479));
    Span4Mux_h I__3423 (
            .O(N__20482),
            .I(N__20476));
    LocalMux I__3422 (
            .O(N__20479),
            .I(alt_kp_4));
    Odrv4 I__3421 (
            .O(N__20476),
            .I(alt_kp_4));
    InMux I__3420 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__3419 (
            .O(N__20468),
            .I(N__20465));
    Span4Mux_h I__3418 (
            .O(N__20465),
            .I(N__20462));
    Odrv4 I__3417 (
            .O(N__20462),
            .I(\pid_alt.O_10 ));
    InMux I__3416 (
            .O(N__20459),
            .I(N__20455));
    InMux I__3415 (
            .O(N__20458),
            .I(N__20452));
    LocalMux I__3414 (
            .O(N__20455),
            .I(N__20449));
    LocalMux I__3413 (
            .O(N__20452),
            .I(N__20446));
    Span4Mux_v I__3412 (
            .O(N__20449),
            .I(N__20443));
    Span12Mux_v I__3411 (
            .O(N__20446),
            .I(N__20440));
    Odrv4 I__3410 (
            .O(N__20443),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    Odrv12 I__3409 (
            .O(N__20440),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    CascadeMux I__3408 (
            .O(N__20435),
            .I(N__20431));
    InMux I__3407 (
            .O(N__20434),
            .I(N__20428));
    InMux I__3406 (
            .O(N__20431),
            .I(N__20425));
    LocalMux I__3405 (
            .O(N__20428),
            .I(N__20422));
    LocalMux I__3404 (
            .O(N__20425),
            .I(N__20418));
    Span4Mux_v I__3403 (
            .O(N__20422),
            .I(N__20415));
    InMux I__3402 (
            .O(N__20421),
            .I(N__20412));
    Span4Mux_v I__3401 (
            .O(N__20418),
            .I(N__20409));
    Span4Mux_v I__3400 (
            .O(N__20415),
            .I(N__20406));
    LocalMux I__3399 (
            .O(N__20412),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    Odrv4 I__3398 (
            .O(N__20409),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    Odrv4 I__3397 (
            .O(N__20406),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__3396 (
            .O(N__20399),
            .I(N__20394));
    InMux I__3395 (
            .O(N__20398),
            .I(N__20391));
    CascadeMux I__3394 (
            .O(N__20397),
            .I(N__20387));
    LocalMux I__3393 (
            .O(N__20394),
            .I(N__20384));
    LocalMux I__3392 (
            .O(N__20391),
            .I(N__20381));
    InMux I__3391 (
            .O(N__20390),
            .I(N__20378));
    InMux I__3390 (
            .O(N__20387),
            .I(N__20375));
    Span4Mux_h I__3389 (
            .O(N__20384),
            .I(N__20372));
    Span4Mux_h I__3388 (
            .O(N__20381),
            .I(N__20367));
    LocalMux I__3387 (
            .O(N__20378),
            .I(N__20367));
    LocalMux I__3386 (
            .O(N__20375),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__3385 (
            .O(N__20372),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__3384 (
            .O(N__20367),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    CascadeMux I__3383 (
            .O(N__20360),
            .I(N__20357));
    InMux I__3382 (
            .O(N__20357),
            .I(N__20354));
    LocalMux I__3381 (
            .O(N__20354),
            .I(N__20351));
    Span4Mux_h I__3380 (
            .O(N__20351),
            .I(N__20348));
    Sp12to4 I__3379 (
            .O(N__20348),
            .I(N__20345));
    Odrv12 I__3378 (
            .O(N__20345),
            .I(\pid_alt.error_p_reg_esr_RNI69J71Z0Z_6 ));
    CascadeMux I__3377 (
            .O(N__20342),
            .I(\pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_ ));
    InMux I__3376 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__3375 (
            .O(N__20336),
            .I(N__20333));
    Span4Mux_v I__3374 (
            .O(N__20333),
            .I(N__20330));
    Span4Mux_v I__3373 (
            .O(N__20330),
            .I(N__20327));
    Odrv4 I__3372 (
            .O(N__20327),
            .I(\pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7 ));
    InMux I__3371 (
            .O(N__20324),
            .I(N__20321));
    LocalMux I__3370 (
            .O(N__20321),
            .I(N__20318));
    Span4Mux_h I__3369 (
            .O(N__20318),
            .I(N__20315));
    Odrv4 I__3368 (
            .O(N__20315),
            .I(\pid_alt.O_11 ));
    CEMux I__3367 (
            .O(N__20312),
            .I(N__20270));
    CEMux I__3366 (
            .O(N__20311),
            .I(N__20270));
    CEMux I__3365 (
            .O(N__20310),
            .I(N__20270));
    CEMux I__3364 (
            .O(N__20309),
            .I(N__20270));
    CEMux I__3363 (
            .O(N__20308),
            .I(N__20270));
    CEMux I__3362 (
            .O(N__20307),
            .I(N__20270));
    CEMux I__3361 (
            .O(N__20306),
            .I(N__20270));
    CEMux I__3360 (
            .O(N__20305),
            .I(N__20270));
    CEMux I__3359 (
            .O(N__20304),
            .I(N__20270));
    CEMux I__3358 (
            .O(N__20303),
            .I(N__20270));
    CEMux I__3357 (
            .O(N__20302),
            .I(N__20270));
    CEMux I__3356 (
            .O(N__20301),
            .I(N__20270));
    CEMux I__3355 (
            .O(N__20300),
            .I(N__20270));
    CEMux I__3354 (
            .O(N__20299),
            .I(N__20270));
    GlobalMux I__3353 (
            .O(N__20270),
            .I(N__20267));
    gio2CtrlBuf I__3352 (
            .O(N__20267),
            .I(\pid_alt.N_422_0_g ));
    InMux I__3351 (
            .O(N__20264),
            .I(N__20258));
    InMux I__3350 (
            .O(N__20263),
            .I(N__20258));
    LocalMux I__3349 (
            .O(N__20258),
            .I(N__20255));
    Span4Mux_v I__3348 (
            .O(N__20255),
            .I(N__20252));
    Odrv4 I__3347 (
            .O(N__20252),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    CascadeMux I__3346 (
            .O(N__20249),
            .I(N__20246));
    InMux I__3345 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__3344 (
            .O(N__20243),
            .I(N__20240));
    Span4Mux_h I__3343 (
            .O(N__20240),
            .I(N__20235));
    InMux I__3342 (
            .O(N__20239),
            .I(N__20230));
    InMux I__3341 (
            .O(N__20238),
            .I(N__20230));
    Odrv4 I__3340 (
            .O(N__20235),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    LocalMux I__3339 (
            .O(N__20230),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__3338 (
            .O(N__20225),
            .I(N__20217));
    InMux I__3337 (
            .O(N__20224),
            .I(N__20217));
    InMux I__3336 (
            .O(N__20223),
            .I(N__20214));
    CascadeMux I__3335 (
            .O(N__20222),
            .I(N__20211));
    LocalMux I__3334 (
            .O(N__20217),
            .I(N__20208));
    LocalMux I__3333 (
            .O(N__20214),
            .I(N__20205));
    InMux I__3332 (
            .O(N__20211),
            .I(N__20202));
    Span4Mux_h I__3331 (
            .O(N__20208),
            .I(N__20197));
    Span4Mux_v I__3330 (
            .O(N__20205),
            .I(N__20197));
    LocalMux I__3329 (
            .O(N__20202),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv4 I__3328 (
            .O(N__20197),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    CascadeMux I__3327 (
            .O(N__20192),
            .I(N__20188));
    CascadeMux I__3326 (
            .O(N__20191),
            .I(N__20185));
    InMux I__3325 (
            .O(N__20188),
            .I(N__20182));
    InMux I__3324 (
            .O(N__20185),
            .I(N__20179));
    LocalMux I__3323 (
            .O(N__20182),
            .I(N__20176));
    LocalMux I__3322 (
            .O(N__20179),
            .I(N__20171));
    Span12Mux_v I__3321 (
            .O(N__20176),
            .I(N__20171));
    Odrv12 I__3320 (
            .O(N__20171),
            .I(\pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7 ));
    CascadeMux I__3319 (
            .O(N__20168),
            .I(N__20165));
    InMux I__3318 (
            .O(N__20165),
            .I(N__20161));
    InMux I__3317 (
            .O(N__20164),
            .I(N__20158));
    LocalMux I__3316 (
            .O(N__20161),
            .I(N__20155));
    LocalMux I__3315 (
            .O(N__20158),
            .I(N__20152));
    Span4Mux_s3_h I__3314 (
            .O(N__20155),
            .I(N__20149));
    Odrv12 I__3313 (
            .O(N__20152),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    Odrv4 I__3312 (
            .O(N__20149),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    InMux I__3311 (
            .O(N__20144),
            .I(N__20141));
    LocalMux I__3310 (
            .O(N__20141),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__3309 (
            .O(N__20138),
            .I(N__20129));
    InMux I__3308 (
            .O(N__20137),
            .I(N__20129));
    InMux I__3307 (
            .O(N__20136),
            .I(N__20129));
    LocalMux I__3306 (
            .O(N__20129),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__3305 (
            .O(N__20126),
            .I(N__20114));
    InMux I__3304 (
            .O(N__20125),
            .I(N__20114));
    InMux I__3303 (
            .O(N__20124),
            .I(N__20114));
    InMux I__3302 (
            .O(N__20123),
            .I(N__20109));
    InMux I__3301 (
            .O(N__20122),
            .I(N__20109));
    InMux I__3300 (
            .O(N__20121),
            .I(N__20102));
    LocalMux I__3299 (
            .O(N__20114),
            .I(N__20095));
    LocalMux I__3298 (
            .O(N__20109),
            .I(N__20095));
    InMux I__3297 (
            .O(N__20108),
            .I(N__20092));
    InMux I__3296 (
            .O(N__20107),
            .I(N__20085));
    InMux I__3295 (
            .O(N__20106),
            .I(N__20085));
    InMux I__3294 (
            .O(N__20105),
            .I(N__20085));
    LocalMux I__3293 (
            .O(N__20102),
            .I(N__20079));
    InMux I__3292 (
            .O(N__20101),
            .I(N__20074));
    InMux I__3291 (
            .O(N__20100),
            .I(N__20074));
    Span4Mux_v I__3290 (
            .O(N__20095),
            .I(N__20068));
    LocalMux I__3289 (
            .O(N__20092),
            .I(N__20065));
    LocalMux I__3288 (
            .O(N__20085),
            .I(N__20062));
    InMux I__3287 (
            .O(N__20084),
            .I(N__20059));
    InMux I__3286 (
            .O(N__20083),
            .I(N__20054));
    InMux I__3285 (
            .O(N__20082),
            .I(N__20054));
    Span4Mux_v I__3284 (
            .O(N__20079),
            .I(N__20049));
    LocalMux I__3283 (
            .O(N__20074),
            .I(N__20049));
    InMux I__3282 (
            .O(N__20073),
            .I(N__20042));
    InMux I__3281 (
            .O(N__20072),
            .I(N__20042));
    InMux I__3280 (
            .O(N__20071),
            .I(N__20042));
    Odrv4 I__3279 (
            .O(N__20068),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__3278 (
            .O(N__20065),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv12 I__3277 (
            .O(N__20062),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3276 (
            .O(N__20059),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3275 (
            .O(N__20054),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__3274 (
            .O(N__20049),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__3273 (
            .O(N__20042),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__3272 (
            .O(N__20027),
            .I(N__20024));
    LocalMux I__3271 (
            .O(N__20024),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__3270 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__3269 (
            .O(N__20018),
            .I(N__20015));
    Span4Mux_s2_v I__3268 (
            .O(N__20015),
            .I(N__20012));
    Odrv4 I__3267 (
            .O(N__20012),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__3266 (
            .O(N__20009),
            .I(N__20000));
    InMux I__3265 (
            .O(N__20008),
            .I(N__20000));
    InMux I__3264 (
            .O(N__20007),
            .I(N__20000));
    LocalMux I__3263 (
            .O(N__20000),
            .I(N__19997));
    Span4Mux_h I__3262 (
            .O(N__19997),
            .I(N__19994));
    Odrv4 I__3261 (
            .O(N__19994),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    CascadeMux I__3260 (
            .O(N__19991),
            .I(N__19988));
    InMux I__3259 (
            .O(N__19988),
            .I(N__19985));
    LocalMux I__3258 (
            .O(N__19985),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    CascadeMux I__3257 (
            .O(N__19982),
            .I(\ppm_encoder_1.N_319_cascade_ ));
    InMux I__3256 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__3255 (
            .O(N__19976),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    CascadeMux I__3254 (
            .O(N__19973),
            .I(N__19970));
    InMux I__3253 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__3252 (
            .O(N__19967),
            .I(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ));
    CascadeMux I__3251 (
            .O(N__19964),
            .I(N__19961));
    InMux I__3250 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__3249 (
            .O(N__19958),
            .I(N__19955));
    Odrv4 I__3248 (
            .O(N__19955),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__3247 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__3246 (
            .O(N__19949),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__3245 (
            .O(N__19946),
            .I(N__19942));
    InMux I__3244 (
            .O(N__19945),
            .I(N__19939));
    LocalMux I__3243 (
            .O(N__19942),
            .I(N__19930));
    LocalMux I__3242 (
            .O(N__19939),
            .I(N__19930));
    InMux I__3241 (
            .O(N__19938),
            .I(N__19923));
    InMux I__3240 (
            .O(N__19937),
            .I(N__19923));
    InMux I__3239 (
            .O(N__19936),
            .I(N__19923));
    CascadeMux I__3238 (
            .O(N__19935),
            .I(N__19918));
    Span4Mux_v I__3237 (
            .O(N__19930),
            .I(N__19914));
    LocalMux I__3236 (
            .O(N__19923),
            .I(N__19911));
    InMux I__3235 (
            .O(N__19922),
            .I(N__19906));
    InMux I__3234 (
            .O(N__19921),
            .I(N__19906));
    InMux I__3233 (
            .O(N__19918),
            .I(N__19901));
    InMux I__3232 (
            .O(N__19917),
            .I(N__19901));
    Odrv4 I__3231 (
            .O(N__19914),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    Odrv4 I__3230 (
            .O(N__19911),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__3229 (
            .O(N__19906),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__3228 (
            .O(N__19901),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    CascadeMux I__3227 (
            .O(N__19892),
            .I(N__19889));
    InMux I__3226 (
            .O(N__19889),
            .I(N__19886));
    LocalMux I__3225 (
            .O(N__19886),
            .I(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ));
    CascadeMux I__3224 (
            .O(N__19883),
            .I(N__19880));
    InMux I__3223 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__3222 (
            .O(N__19877),
            .I(N__19874));
    Span4Mux_h I__3221 (
            .O(N__19874),
            .I(N__19871));
    Odrv4 I__3220 (
            .O(N__19871),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__3219 (
            .O(N__19868),
            .I(N__19865));
    LocalMux I__3218 (
            .O(N__19865),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__3217 (
            .O(N__19862),
            .I(N__19858));
    InMux I__3216 (
            .O(N__19861),
            .I(N__19855));
    LocalMux I__3215 (
            .O(N__19858),
            .I(N__19852));
    LocalMux I__3214 (
            .O(N__19855),
            .I(N__19849));
    Span4Mux_v I__3213 (
            .O(N__19852),
            .I(N__19846));
    Span4Mux_h I__3212 (
            .O(N__19849),
            .I(N__19843));
    Odrv4 I__3211 (
            .O(N__19846),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    Odrv4 I__3210 (
            .O(N__19843),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    CascadeMux I__3209 (
            .O(N__19838),
            .I(N__19834));
    CascadeMux I__3208 (
            .O(N__19837),
            .I(N__19830));
    InMux I__3207 (
            .O(N__19834),
            .I(N__19825));
    InMux I__3206 (
            .O(N__19833),
            .I(N__19825));
    InMux I__3205 (
            .O(N__19830),
            .I(N__19822));
    LocalMux I__3204 (
            .O(N__19825),
            .I(N__19817));
    LocalMux I__3203 (
            .O(N__19822),
            .I(N__19817));
    Span4Mux_s3_h I__3202 (
            .O(N__19817),
            .I(N__19814));
    Odrv4 I__3201 (
            .O(N__19814),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    CascadeMux I__3200 (
            .O(N__19811),
            .I(N__19808));
    InMux I__3199 (
            .O(N__19808),
            .I(N__19805));
    LocalMux I__3198 (
            .O(N__19805),
            .I(N__19802));
    Odrv4 I__3197 (
            .O(N__19802),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__3196 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__3195 (
            .O(N__19796),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__3194 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__3193 (
            .O(N__19790),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__3192 (
            .O(N__19787),
            .I(N__19784));
    LocalMux I__3191 (
            .O(N__19784),
            .I(N__19781));
    Span4Mux_s2_v I__3190 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__3189 (
            .O(N__19778),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__3188 (
            .O(N__19775),
            .I(N__19771));
    InMux I__3187 (
            .O(N__19774),
            .I(N__19768));
    LocalMux I__3186 (
            .O(N__19771),
            .I(N__19765));
    LocalMux I__3185 (
            .O(N__19768),
            .I(N__19762));
    Odrv12 I__3184 (
            .O(N__19765),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    Odrv4 I__3183 (
            .O(N__19762),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__3182 (
            .O(N__19757),
            .I(N__19754));
    LocalMux I__3181 (
            .O(N__19754),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__3180 (
            .O(N__19751),
            .I(N__19748));
    LocalMux I__3179 (
            .O(N__19748),
            .I(N__19745));
    Odrv4 I__3178 (
            .O(N__19745),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__3177 (
            .O(N__19742),
            .I(N__19739));
    LocalMux I__3176 (
            .O(N__19739),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__3175 (
            .O(N__19736),
            .I(N__19733));
    LocalMux I__3174 (
            .O(N__19733),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__3173 (
            .O(N__19730),
            .I(N__19727));
    LocalMux I__3172 (
            .O(N__19727),
            .I(N__19724));
    Span4Mux_h I__3171 (
            .O(N__19724),
            .I(N__19721));
    Odrv4 I__3170 (
            .O(N__19721),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__3169 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__3168 (
            .O(N__19715),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__3167 (
            .O(N__19712),
            .I(N__19709));
    LocalMux I__3166 (
            .O(N__19709),
            .I(N__19705));
    InMux I__3165 (
            .O(N__19708),
            .I(N__19702));
    Span4Mux_s3_h I__3164 (
            .O(N__19705),
            .I(N__19697));
    LocalMux I__3163 (
            .O(N__19702),
            .I(N__19697));
    Odrv4 I__3162 (
            .O(N__19697),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    InMux I__3161 (
            .O(N__19694),
            .I(N__19685));
    InMux I__3160 (
            .O(N__19693),
            .I(N__19685));
    InMux I__3159 (
            .O(N__19692),
            .I(N__19685));
    LocalMux I__3158 (
            .O(N__19685),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__3157 (
            .O(N__19682),
            .I(N__19679));
    LocalMux I__3156 (
            .O(N__19679),
            .I(N__19676));
    Odrv4 I__3155 (
            .O(N__19676),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    CascadeMux I__3154 (
            .O(N__19673),
            .I(N__19670));
    InMux I__3153 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__3152 (
            .O(N__19667),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__3151 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__3150 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_s3_h I__3149 (
            .O(N__19658),
            .I(N__19655));
    Odrv4 I__3148 (
            .O(N__19655),
            .I(\ppm_encoder_1.un1_init_pulses_11_0 ));
    InMux I__3147 (
            .O(N__19652),
            .I(N__19648));
    InMux I__3146 (
            .O(N__19651),
            .I(N__19645));
    LocalMux I__3145 (
            .O(N__19648),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    LocalMux I__3144 (
            .O(N__19645),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    CascadeMux I__3143 (
            .O(N__19640),
            .I(N__19637));
    InMux I__3142 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__3141 (
            .O(N__19634),
            .I(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ));
    InMux I__3140 (
            .O(N__19631),
            .I(N__19628));
    LocalMux I__3139 (
            .O(N__19628),
            .I(N__19625));
    Span4Mux_h I__3138 (
            .O(N__19625),
            .I(N__19622));
    Odrv4 I__3137 (
            .O(N__19622),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ));
    CascadeMux I__3136 (
            .O(N__19619),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ));
    InMux I__3135 (
            .O(N__19616),
            .I(N__19613));
    LocalMux I__3134 (
            .O(N__19613),
            .I(N__19610));
    Span4Mux_v I__3133 (
            .O(N__19610),
            .I(N__19606));
    InMux I__3132 (
            .O(N__19609),
            .I(N__19603));
    Odrv4 I__3131 (
            .O(N__19606),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    LocalMux I__3130 (
            .O(N__19603),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    InMux I__3129 (
            .O(N__19598),
            .I(N__19593));
    InMux I__3128 (
            .O(N__19597),
            .I(N__19588));
    InMux I__3127 (
            .O(N__19596),
            .I(N__19588));
    LocalMux I__3126 (
            .O(N__19593),
            .I(N__19585));
    LocalMux I__3125 (
            .O(N__19588),
            .I(N__19580));
    Span4Mux_v I__3124 (
            .O(N__19585),
            .I(N__19580));
    Odrv4 I__3123 (
            .O(N__19580),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__3122 (
            .O(N__19577),
            .I(N__19573));
    InMux I__3121 (
            .O(N__19576),
            .I(N__19570));
    LocalMux I__3120 (
            .O(N__19573),
            .I(N__19565));
    LocalMux I__3119 (
            .O(N__19570),
            .I(N__19565));
    Odrv4 I__3118 (
            .O(N__19565),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    InMux I__3117 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__3116 (
            .O(N__19559),
            .I(N__19556));
    Span4Mux_v I__3115 (
            .O(N__19556),
            .I(N__19553));
    Span4Mux_s3_h I__3114 (
            .O(N__19553),
            .I(N__19549));
    InMux I__3113 (
            .O(N__19552),
            .I(N__19546));
    Odrv4 I__3112 (
            .O(N__19549),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    LocalMux I__3111 (
            .O(N__19546),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    InMux I__3110 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__3109 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_h I__3108 (
            .O(N__19535),
            .I(N__19532));
    Odrv4 I__3107 (
            .O(N__19532),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    CascadeMux I__3106 (
            .O(N__19529),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ));
    InMux I__3105 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__3104 (
            .O(N__19523),
            .I(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ));
    CascadeMux I__3103 (
            .O(N__19520),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ));
    CascadeMux I__3102 (
            .O(N__19517),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    InMux I__3101 (
            .O(N__19514),
            .I(N__19511));
    LocalMux I__3100 (
            .O(N__19511),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4 ));
    CascadeMux I__3099 (
            .O(N__19508),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ));
    CascadeMux I__3098 (
            .O(N__19505),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    CascadeMux I__3097 (
            .O(N__19502),
            .I(N__19499));
    InMux I__3096 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__3095 (
            .O(N__19496),
            .I(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ));
    CascadeMux I__3094 (
            .O(N__19493),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    InMux I__3093 (
            .O(N__19490),
            .I(N__19485));
    InMux I__3092 (
            .O(N__19489),
            .I(N__19482));
    InMux I__3091 (
            .O(N__19488),
            .I(N__19477));
    LocalMux I__3090 (
            .O(N__19485),
            .I(N__19472));
    LocalMux I__3089 (
            .O(N__19482),
            .I(N__19472));
    InMux I__3088 (
            .O(N__19481),
            .I(N__19469));
    InMux I__3087 (
            .O(N__19480),
            .I(N__19466));
    LocalMux I__3086 (
            .O(N__19477),
            .I(N__19463));
    Span4Mux_v I__3085 (
            .O(N__19472),
            .I(N__19456));
    LocalMux I__3084 (
            .O(N__19469),
            .I(N__19456));
    LocalMux I__3083 (
            .O(N__19466),
            .I(N__19456));
    Odrv4 I__3082 (
            .O(N__19463),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    Odrv4 I__3081 (
            .O(N__19456),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    CascadeMux I__3080 (
            .O(N__19451),
            .I(\pid_alt.N_88_cascade_ ));
    InMux I__3079 (
            .O(N__19448),
            .I(N__19442));
    InMux I__3078 (
            .O(N__19447),
            .I(N__19442));
    LocalMux I__3077 (
            .O(N__19442),
            .I(N__19438));
    InMux I__3076 (
            .O(N__19441),
            .I(N__19435));
    Odrv4 I__3075 (
            .O(N__19438),
            .I(\pid_alt.N_90 ));
    LocalMux I__3074 (
            .O(N__19435),
            .I(\pid_alt.N_90 ));
    CascadeMux I__3073 (
            .O(N__19430),
            .I(N__19427));
    InMux I__3072 (
            .O(N__19427),
            .I(N__19420));
    InMux I__3071 (
            .O(N__19426),
            .I(N__19420));
    CascadeMux I__3070 (
            .O(N__19425),
            .I(N__19416));
    LocalMux I__3069 (
            .O(N__19420),
            .I(N__19410));
    InMux I__3068 (
            .O(N__19419),
            .I(N__19403));
    InMux I__3067 (
            .O(N__19416),
            .I(N__19403));
    InMux I__3066 (
            .O(N__19415),
            .I(N__19403));
    CascadeMux I__3065 (
            .O(N__19414),
            .I(N__19399));
    CascadeMux I__3064 (
            .O(N__19413),
            .I(N__19395));
    Span4Mux_v I__3063 (
            .O(N__19410),
            .I(N__19391));
    LocalMux I__3062 (
            .O(N__19403),
            .I(N__19388));
    InMux I__3061 (
            .O(N__19402),
            .I(N__19381));
    InMux I__3060 (
            .O(N__19399),
            .I(N__19381));
    InMux I__3059 (
            .O(N__19398),
            .I(N__19381));
    InMux I__3058 (
            .O(N__19395),
            .I(N__19378));
    InMux I__3057 (
            .O(N__19394),
            .I(N__19375));
    Odrv4 I__3056 (
            .O(N__19391),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    Odrv4 I__3055 (
            .O(N__19388),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    LocalMux I__3054 (
            .O(N__19381),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    LocalMux I__3053 (
            .O(N__19378),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    LocalMux I__3052 (
            .O(N__19375),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__3051 (
            .O(N__19364),
            .I(N__19361));
    LocalMux I__3050 (
            .O(N__19361),
            .I(N__19357));
    InMux I__3049 (
            .O(N__19360),
            .I(N__19354));
    Span4Mux_v I__3048 (
            .O(N__19357),
            .I(N__19349));
    LocalMux I__3047 (
            .O(N__19354),
            .I(N__19349));
    Odrv4 I__3046 (
            .O(N__19349),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    CascadeMux I__3045 (
            .O(N__19346),
            .I(\pid_alt.N_90_cascade_ ));
    InMux I__3044 (
            .O(N__19343),
            .I(N__19337));
    InMux I__3043 (
            .O(N__19342),
            .I(N__19337));
    LocalMux I__3042 (
            .O(N__19337),
            .I(N__19327));
    InMux I__3041 (
            .O(N__19336),
            .I(N__19324));
    InMux I__3040 (
            .O(N__19335),
            .I(N__19319));
    InMux I__3039 (
            .O(N__19334),
            .I(N__19310));
    InMux I__3038 (
            .O(N__19333),
            .I(N__19310));
    InMux I__3037 (
            .O(N__19332),
            .I(N__19310));
    InMux I__3036 (
            .O(N__19331),
            .I(N__19310));
    InMux I__3035 (
            .O(N__19330),
            .I(N__19307));
    Span4Mux_v I__3034 (
            .O(N__19327),
            .I(N__19302));
    LocalMux I__3033 (
            .O(N__19324),
            .I(N__19302));
    InMux I__3032 (
            .O(N__19323),
            .I(N__19297));
    InMux I__3031 (
            .O(N__19322),
            .I(N__19297));
    LocalMux I__3030 (
            .O(N__19319),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ));
    LocalMux I__3029 (
            .O(N__19310),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ));
    LocalMux I__3028 (
            .O(N__19307),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ));
    Odrv4 I__3027 (
            .O(N__19302),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ));
    LocalMux I__3026 (
            .O(N__19297),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ));
    CEMux I__3025 (
            .O(N__19286),
            .I(N__19281));
    CEMux I__3024 (
            .O(N__19285),
            .I(N__19278));
    CEMux I__3023 (
            .O(N__19284),
            .I(N__19275));
    LocalMux I__3022 (
            .O(N__19281),
            .I(N__19270));
    LocalMux I__3021 (
            .O(N__19278),
            .I(N__19270));
    LocalMux I__3020 (
            .O(N__19275),
            .I(N__19265));
    Span4Mux_v I__3019 (
            .O(N__19270),
            .I(N__19265));
    Odrv4 I__3018 (
            .O(N__19265),
            .I(\pid_alt.N_60_i_1 ));
    SRMux I__3017 (
            .O(N__19262),
            .I(N__19257));
    SRMux I__3016 (
            .O(N__19261),
            .I(N__19253));
    SRMux I__3015 (
            .O(N__19260),
            .I(N__19250));
    LocalMux I__3014 (
            .O(N__19257),
            .I(N__19246));
    SRMux I__3013 (
            .O(N__19256),
            .I(N__19243));
    LocalMux I__3012 (
            .O(N__19253),
            .I(N__19240));
    LocalMux I__3011 (
            .O(N__19250),
            .I(N__19237));
    SRMux I__3010 (
            .O(N__19249),
            .I(N__19234));
    Odrv4 I__3009 (
            .O(N__19246),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__3008 (
            .O(N__19243),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv12 I__3007 (
            .O(N__19240),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv12 I__3006 (
            .O(N__19237),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__3005 (
            .O(N__19234),
            .I(\pid_alt.un1_reset_0_i ));
    CascadeMux I__3004 (
            .O(N__19223),
            .I(N__19219));
    InMux I__3003 (
            .O(N__19222),
            .I(N__19216));
    InMux I__3002 (
            .O(N__19219),
            .I(N__19213));
    LocalMux I__3001 (
            .O(N__19216),
            .I(N__19210));
    LocalMux I__3000 (
            .O(N__19213),
            .I(N__19207));
    Span4Mux_v I__2999 (
            .O(N__19210),
            .I(N__19204));
    Odrv12 I__2998 (
            .O(N__19207),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    Odrv4 I__2997 (
            .O(N__19204),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__2996 (
            .O(N__19199),
            .I(N__19192));
    InMux I__2995 (
            .O(N__19198),
            .I(N__19192));
    InMux I__2994 (
            .O(N__19197),
            .I(N__19189));
    LocalMux I__2993 (
            .O(N__19192),
            .I(N__19185));
    LocalMux I__2992 (
            .O(N__19189),
            .I(N__19182));
    InMux I__2991 (
            .O(N__19188),
            .I(N__19179));
    Span4Mux_v I__2990 (
            .O(N__19185),
            .I(N__19176));
    Odrv4 I__2989 (
            .O(N__19182),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    LocalMux I__2988 (
            .O(N__19179),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__2987 (
            .O(N__19176),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    CascadeMux I__2986 (
            .O(N__19169),
            .I(N__19166));
    InMux I__2985 (
            .O(N__19166),
            .I(N__19161));
    InMux I__2984 (
            .O(N__19165),
            .I(N__19158));
    InMux I__2983 (
            .O(N__19164),
            .I(N__19155));
    LocalMux I__2982 (
            .O(N__19161),
            .I(N__19151));
    LocalMux I__2981 (
            .O(N__19158),
            .I(N__19146));
    LocalMux I__2980 (
            .O(N__19155),
            .I(N__19146));
    InMux I__2979 (
            .O(N__19154),
            .I(N__19143));
    Span4Mux_v I__2978 (
            .O(N__19151),
            .I(N__19138));
    Span4Mux_v I__2977 (
            .O(N__19146),
            .I(N__19138));
    LocalMux I__2976 (
            .O(N__19143),
            .I(\pid_alt.N_130 ));
    Odrv4 I__2975 (
            .O(N__19138),
            .I(\pid_alt.N_130 ));
    CascadeMux I__2974 (
            .O(N__19133),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ));
    InMux I__2973 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__2972 (
            .O(N__19127),
            .I(N__19123));
    InMux I__2971 (
            .O(N__19126),
            .I(N__19120));
    Span4Mux_v I__2970 (
            .O(N__19123),
            .I(N__19117));
    LocalMux I__2969 (
            .O(N__19120),
            .I(N__19114));
    Span4Mux_v I__2968 (
            .O(N__19117),
            .I(N__19111));
    Span4Mux_h I__2967 (
            .O(N__19114),
            .I(N__19108));
    Odrv4 I__2966 (
            .O(N__19111),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    Odrv4 I__2965 (
            .O(N__19108),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    CascadeMux I__2964 (
            .O(N__19103),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    CascadeMux I__2963 (
            .O(N__19100),
            .I(N__19097));
    InMux I__2962 (
            .O(N__19097),
            .I(N__19094));
    LocalMux I__2961 (
            .O(N__19094),
            .I(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ));
    InMux I__2960 (
            .O(N__19091),
            .I(N__19088));
    LocalMux I__2959 (
            .O(N__19088),
            .I(N__19085));
    Span4Mux_s3_h I__2958 (
            .O(N__19085),
            .I(N__19082));
    Span4Mux_v I__2957 (
            .O(N__19082),
            .I(N__19079));
    Odrv4 I__2956 (
            .O(N__19079),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__2955 (
            .O(N__19076),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__2954 (
            .O(N__19073),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__2953 (
            .O(N__19070),
            .I(N__19067));
    LocalMux I__2952 (
            .O(N__19067),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__2951 (
            .O(N__19064),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__2950 (
            .O(N__19061),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__2949 (
            .O(N__19058),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__2948 (
            .O(N__19055),
            .I(bfn_3_22_0_));
    InMux I__2947 (
            .O(N__19052),
            .I(N__19048));
    InMux I__2946 (
            .O(N__19051),
            .I(N__19045));
    LocalMux I__2945 (
            .O(N__19048),
            .I(N__19042));
    LocalMux I__2944 (
            .O(N__19045),
            .I(N__19039));
    Span4Mux_v I__2943 (
            .O(N__19042),
            .I(N__19036));
    Odrv12 I__2942 (
            .O(N__19039),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    Odrv4 I__2941 (
            .O(N__19036),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    InMux I__2940 (
            .O(N__19031),
            .I(N__19027));
    CascadeMux I__2939 (
            .O(N__19030),
            .I(N__19024));
    LocalMux I__2938 (
            .O(N__19027),
            .I(N__19021));
    InMux I__2937 (
            .O(N__19024),
            .I(N__19018));
    Span4Mux_v I__2936 (
            .O(N__19021),
            .I(N__19013));
    LocalMux I__2935 (
            .O(N__19018),
            .I(N__19013));
    Odrv4 I__2934 (
            .O(N__19013),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    CascadeMux I__2933 (
            .O(N__19010),
            .I(N__19006));
    InMux I__2932 (
            .O(N__19009),
            .I(N__19002));
    InMux I__2931 (
            .O(N__19006),
            .I(N__18995));
    InMux I__2930 (
            .O(N__19005),
            .I(N__18995));
    LocalMux I__2929 (
            .O(N__19002),
            .I(N__18991));
    InMux I__2928 (
            .O(N__19001),
            .I(N__18986));
    InMux I__2927 (
            .O(N__19000),
            .I(N__18986));
    LocalMux I__2926 (
            .O(N__18995),
            .I(N__18983));
    InMux I__2925 (
            .O(N__18994),
            .I(N__18980));
    Span4Mux_v I__2924 (
            .O(N__18991),
            .I(N__18975));
    LocalMux I__2923 (
            .O(N__18986),
            .I(N__18975));
    Odrv12 I__2922 (
            .O(N__18983),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    LocalMux I__2921 (
            .O(N__18980),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__2920 (
            .O(N__18975),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    InMux I__2919 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__2918 (
            .O(N__18965),
            .I(N__18961));
    InMux I__2917 (
            .O(N__18964),
            .I(N__18958));
    Odrv12 I__2916 (
            .O(N__18961),
            .I(\pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6 ));
    LocalMux I__2915 (
            .O(N__18958),
            .I(\pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6 ));
    InMux I__2914 (
            .O(N__18953),
            .I(N__18947));
    InMux I__2913 (
            .O(N__18952),
            .I(N__18947));
    LocalMux I__2912 (
            .O(N__18947),
            .I(N__18944));
    Odrv4 I__2911 (
            .O(N__18944),
            .I(\pid_alt.N_88 ));
    CascadeMux I__2910 (
            .O(N__18941),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ));
    InMux I__2909 (
            .O(N__18938),
            .I(N__18934));
    InMux I__2908 (
            .O(N__18937),
            .I(N__18931));
    LocalMux I__2907 (
            .O(N__18934),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    LocalMux I__2906 (
            .O(N__18931),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    CascadeMux I__2905 (
            .O(N__18926),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ));
    CascadeMux I__2904 (
            .O(N__18923),
            .I(\pid_alt.N_92_cascade_ ));
    CascadeMux I__2903 (
            .O(N__18920),
            .I(\pid_alt.un1_reset_1_cascade_ ));
    InMux I__2902 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__2901 (
            .O(N__18914),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ));
    CascadeMux I__2900 (
            .O(N__18911),
            .I(\pid_alt.un1_reset_0_i_cascade_ ));
    InMux I__2899 (
            .O(N__18908),
            .I(N__18905));
    LocalMux I__2898 (
            .O(N__18905),
            .I(N__18902));
    Sp12to4 I__2897 (
            .O(N__18902),
            .I(N__18899));
    Odrv12 I__2896 (
            .O(N__18899),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__2895 (
            .O(N__18896),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__2894 (
            .O(N__18893),
            .I(\ppm_encoder_1.un1_aileron_cry_7 ));
    InMux I__2893 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__2892 (
            .O(N__18887),
            .I(N__18884));
    Odrv4 I__2891 (
            .O(N__18884),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO ));
    CascadeMux I__2890 (
            .O(N__18881),
            .I(N__18878));
    InMux I__2889 (
            .O(N__18878),
            .I(N__18874));
    InMux I__2888 (
            .O(N__18877),
            .I(N__18871));
    LocalMux I__2887 (
            .O(N__18874),
            .I(N__18865));
    LocalMux I__2886 (
            .O(N__18871),
            .I(N__18865));
    InMux I__2885 (
            .O(N__18870),
            .I(N__18862));
    Span4Mux_v I__2884 (
            .O(N__18865),
            .I(N__18857));
    LocalMux I__2883 (
            .O(N__18862),
            .I(N__18854));
    InMux I__2882 (
            .O(N__18861),
            .I(N__18849));
    InMux I__2881 (
            .O(N__18860),
            .I(N__18849));
    Span4Mux_v I__2880 (
            .O(N__18857),
            .I(N__18846));
    Span4Mux_v I__2879 (
            .O(N__18854),
            .I(N__18841));
    LocalMux I__2878 (
            .O(N__18849),
            .I(N__18841));
    Odrv4 I__2877 (
            .O(N__18846),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    Odrv4 I__2876 (
            .O(N__18841),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__2875 (
            .O(N__18836),
            .I(N__18830));
    InMux I__2874 (
            .O(N__18835),
            .I(N__18830));
    LocalMux I__2873 (
            .O(N__18830),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    InMux I__2872 (
            .O(N__18827),
            .I(N__18824));
    LocalMux I__2871 (
            .O(N__18824),
            .I(N__18821));
    Odrv12 I__2870 (
            .O(N__18821),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO ));
    InMux I__2869 (
            .O(N__18818),
            .I(N__18812));
    InMux I__2868 (
            .O(N__18817),
            .I(N__18812));
    LocalMux I__2867 (
            .O(N__18812),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    CascadeMux I__2866 (
            .O(N__18809),
            .I(N__18806));
    InMux I__2865 (
            .O(N__18806),
            .I(N__18791));
    InMux I__2864 (
            .O(N__18805),
            .I(N__18791));
    InMux I__2863 (
            .O(N__18804),
            .I(N__18791));
    InMux I__2862 (
            .O(N__18803),
            .I(N__18791));
    InMux I__2861 (
            .O(N__18802),
            .I(N__18791));
    LocalMux I__2860 (
            .O(N__18791),
            .I(N__18788));
    Span4Mux_h I__2859 (
            .O(N__18788),
            .I(N__18785));
    Odrv4 I__2858 (
            .O(N__18785),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    CascadeMux I__2857 (
            .O(N__18782),
            .I(\pid_alt.source_pid_9_0_tz_6_cascade_ ));
    InMux I__2856 (
            .O(N__18779),
            .I(N__18776));
    LocalMux I__2855 (
            .O(N__18776),
            .I(N__18771));
    InMux I__2854 (
            .O(N__18775),
            .I(N__18766));
    InMux I__2853 (
            .O(N__18774),
            .I(N__18766));
    Odrv4 I__2852 (
            .O(N__18771),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    LocalMux I__2851 (
            .O(N__18766),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    InMux I__2850 (
            .O(N__18761),
            .I(N__18758));
    LocalMux I__2849 (
            .O(N__18758),
            .I(N__18755));
    Span4Mux_s2_h I__2848 (
            .O(N__18755),
            .I(N__18750));
    InMux I__2847 (
            .O(N__18754),
            .I(N__18747));
    InMux I__2846 (
            .O(N__18753),
            .I(N__18744));
    Odrv4 I__2845 (
            .O(N__18750),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    LocalMux I__2844 (
            .O(N__18747),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    LocalMux I__2843 (
            .O(N__18744),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    InMux I__2842 (
            .O(N__18737),
            .I(N__18733));
    CascadeMux I__2841 (
            .O(N__18736),
            .I(N__18730));
    LocalMux I__2840 (
            .O(N__18733),
            .I(N__18726));
    InMux I__2839 (
            .O(N__18730),
            .I(N__18723));
    InMux I__2838 (
            .O(N__18729),
            .I(N__18720));
    Odrv4 I__2837 (
            .O(N__18726),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    LocalMux I__2836 (
            .O(N__18723),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    LocalMux I__2835 (
            .O(N__18720),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    CascadeMux I__2834 (
            .O(N__18713),
            .I(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ));
    InMux I__2833 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__2832 (
            .O(N__18707),
            .I(N__18702));
    InMux I__2831 (
            .O(N__18706),
            .I(N__18699));
    CascadeMux I__2830 (
            .O(N__18705),
            .I(N__18696));
    Span4Mux_v I__2829 (
            .O(N__18702),
            .I(N__18693));
    LocalMux I__2828 (
            .O(N__18699),
            .I(N__18690));
    InMux I__2827 (
            .O(N__18696),
            .I(N__18687));
    Odrv4 I__2826 (
            .O(N__18693),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    Odrv4 I__2825 (
            .O(N__18690),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    LocalMux I__2824 (
            .O(N__18687),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    CascadeMux I__2823 (
            .O(N__18680),
            .I(N__18677));
    InMux I__2822 (
            .O(N__18677),
            .I(N__18673));
    InMux I__2821 (
            .O(N__18676),
            .I(N__18670));
    LocalMux I__2820 (
            .O(N__18673),
            .I(N__18667));
    LocalMux I__2819 (
            .O(N__18670),
            .I(N__18664));
    Odrv12 I__2818 (
            .O(N__18667),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    Odrv4 I__2817 (
            .O(N__18664),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    InMux I__2816 (
            .O(N__18659),
            .I(N__18656));
    LocalMux I__2815 (
            .O(N__18656),
            .I(N__18651));
    InMux I__2814 (
            .O(N__18655),
            .I(N__18646));
    InMux I__2813 (
            .O(N__18654),
            .I(N__18646));
    Odrv4 I__2812 (
            .O(N__18651),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    LocalMux I__2811 (
            .O(N__18646),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    InMux I__2810 (
            .O(N__18641),
            .I(N__18638));
    LocalMux I__2809 (
            .O(N__18638),
            .I(N__18633));
    InMux I__2808 (
            .O(N__18637),
            .I(N__18628));
    InMux I__2807 (
            .O(N__18636),
            .I(N__18628));
    Odrv4 I__2806 (
            .O(N__18633),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    LocalMux I__2805 (
            .O(N__18628),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    CascadeMux I__2804 (
            .O(N__18623),
            .I(N__18620));
    InMux I__2803 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__2802 (
            .O(N__18617),
            .I(N__18614));
    Odrv4 I__2801 (
            .O(N__18614),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ));
    InMux I__2800 (
            .O(N__18611),
            .I(N__18608));
    LocalMux I__2799 (
            .O(N__18608),
            .I(N__18605));
    Span4Mux_v I__2798 (
            .O(N__18605),
            .I(N__18601));
    InMux I__2797 (
            .O(N__18604),
            .I(N__18598));
    Span4Mux_v I__2796 (
            .O(N__18601),
            .I(N__18591));
    LocalMux I__2795 (
            .O(N__18598),
            .I(N__18591));
    InMux I__2794 (
            .O(N__18597),
            .I(N__18586));
    InMux I__2793 (
            .O(N__18596),
            .I(N__18586));
    Span4Mux_v I__2792 (
            .O(N__18591),
            .I(N__18582));
    LocalMux I__2791 (
            .O(N__18586),
            .I(N__18579));
    InMux I__2790 (
            .O(N__18585),
            .I(N__18576));
    Span4Mux_v I__2789 (
            .O(N__18582),
            .I(N__18573));
    Odrv12 I__2788 (
            .O(N__18579),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    LocalMux I__2787 (
            .O(N__18576),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    Odrv4 I__2786 (
            .O(N__18573),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__2785 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__2784 (
            .O(N__18563),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO ));
    CascadeMux I__2783 (
            .O(N__18560),
            .I(N__18556));
    CascadeMux I__2782 (
            .O(N__18559),
            .I(N__18553));
    InMux I__2781 (
            .O(N__18556),
            .I(N__18549));
    InMux I__2780 (
            .O(N__18553),
            .I(N__18544));
    InMux I__2779 (
            .O(N__18552),
            .I(N__18544));
    LocalMux I__2778 (
            .O(N__18549),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__2777 (
            .O(N__18544),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__2776 (
            .O(N__18539),
            .I(N__18535));
    InMux I__2775 (
            .O(N__18538),
            .I(N__18532));
    LocalMux I__2774 (
            .O(N__18535),
            .I(N__18529));
    LocalMux I__2773 (
            .O(N__18532),
            .I(N__18526));
    Span4Mux_v I__2772 (
            .O(N__18529),
            .I(N__18522));
    Span12Mux_v I__2771 (
            .O(N__18526),
            .I(N__18519));
    InMux I__2770 (
            .O(N__18525),
            .I(N__18516));
    Odrv4 I__2769 (
            .O(N__18522),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    Odrv12 I__2768 (
            .O(N__18519),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    LocalMux I__2767 (
            .O(N__18516),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    InMux I__2766 (
            .O(N__18509),
            .I(N__18504));
    InMux I__2765 (
            .O(N__18508),
            .I(N__18499));
    InMux I__2764 (
            .O(N__18507),
            .I(N__18499));
    LocalMux I__2763 (
            .O(N__18504),
            .I(N__18493));
    LocalMux I__2762 (
            .O(N__18499),
            .I(N__18493));
    CascadeMux I__2761 (
            .O(N__18498),
            .I(N__18490));
    Span4Mux_v I__2760 (
            .O(N__18493),
            .I(N__18486));
    InMux I__2759 (
            .O(N__18490),
            .I(N__18483));
    InMux I__2758 (
            .O(N__18489),
            .I(N__18480));
    Span4Mux_h I__2757 (
            .O(N__18486),
            .I(N__18477));
    LocalMux I__2756 (
            .O(N__18483),
            .I(N__18474));
    LocalMux I__2755 (
            .O(N__18480),
            .I(N__18471));
    Span4Mux_v I__2754 (
            .O(N__18477),
            .I(N__18468));
    Odrv4 I__2753 (
            .O(N__18474),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    Odrv4 I__2752 (
            .O(N__18471),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    Odrv4 I__2751 (
            .O(N__18468),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    CascadeMux I__2750 (
            .O(N__18461),
            .I(N__18458));
    InMux I__2749 (
            .O(N__18458),
            .I(N__18455));
    LocalMux I__2748 (
            .O(N__18455),
            .I(N__18452));
    Span4Mux_h I__2747 (
            .O(N__18452),
            .I(N__18449));
    Odrv4 I__2746 (
            .O(N__18449),
            .I(\pid_alt.error_p_reg_esr_RNIB03KZ0Z_16 ));
    InMux I__2745 (
            .O(N__18446),
            .I(N__18443));
    LocalMux I__2744 (
            .O(N__18443),
            .I(N__18440));
    Span4Mux_v I__2743 (
            .O(N__18440),
            .I(N__18437));
    Span4Mux_v I__2742 (
            .O(N__18437),
            .I(N__18434));
    Odrv4 I__2741 (
            .O(N__18434),
            .I(\ppm_encoder_1.N_306 ));
    CascadeMux I__2740 (
            .O(N__18431),
            .I(\dron_frame_decoder_1.N_194_4_cascade_ ));
    CascadeMux I__2739 (
            .O(N__18428),
            .I(N__18424));
    InMux I__2738 (
            .O(N__18427),
            .I(N__18421));
    InMux I__2737 (
            .O(N__18424),
            .I(N__18418));
    LocalMux I__2736 (
            .O(N__18421),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__2735 (
            .O(N__18418),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__2734 (
            .O(N__18413),
            .I(N__18407));
    InMux I__2733 (
            .O(N__18412),
            .I(N__18407));
    LocalMux I__2732 (
            .O(N__18407),
            .I(\pid_alt.m7_e_4 ));
    InMux I__2731 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__2730 (
            .O(N__18401),
            .I(N__18398));
    Odrv4 I__2729 (
            .O(N__18398),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO ));
    CascadeMux I__2728 (
            .O(N__18395),
            .I(N__18392));
    InMux I__2727 (
            .O(N__18392),
            .I(N__18389));
    LocalMux I__2726 (
            .O(N__18389),
            .I(N__18385));
    CascadeMux I__2725 (
            .O(N__18388),
            .I(N__18382));
    Span4Mux_v I__2724 (
            .O(N__18385),
            .I(N__18378));
    InMux I__2723 (
            .O(N__18382),
            .I(N__18375));
    CascadeMux I__2722 (
            .O(N__18381),
            .I(N__18372));
    Span4Mux_v I__2721 (
            .O(N__18378),
            .I(N__18367));
    LocalMux I__2720 (
            .O(N__18375),
            .I(N__18364));
    InMux I__2719 (
            .O(N__18372),
            .I(N__18357));
    InMux I__2718 (
            .O(N__18371),
            .I(N__18357));
    InMux I__2717 (
            .O(N__18370),
            .I(N__18357));
    Span4Mux_h I__2716 (
            .O(N__18367),
            .I(N__18352));
    Span4Mux_v I__2715 (
            .O(N__18364),
            .I(N__18352));
    LocalMux I__2714 (
            .O(N__18357),
            .I(N__18349));
    Odrv4 I__2713 (
            .O(N__18352),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    Odrv4 I__2712 (
            .O(N__18349),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__2711 (
            .O(N__18344),
            .I(N__18338));
    InMux I__2710 (
            .O(N__18343),
            .I(N__18338));
    LocalMux I__2709 (
            .O(N__18338),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    InMux I__2708 (
            .O(N__18335),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__2707 (
            .O(N__18332),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__2706 (
            .O(N__18329),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__2705 (
            .O(N__18326),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__2704 (
            .O(N__18323),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__2703 (
            .O(N__18320),
            .I(N__18312));
    InMux I__2702 (
            .O(N__18319),
            .I(N__18312));
    InMux I__2701 (
            .O(N__18318),
            .I(N__18307));
    InMux I__2700 (
            .O(N__18317),
            .I(N__18307));
    LocalMux I__2699 (
            .O(N__18312),
            .I(N__18304));
    LocalMux I__2698 (
            .O(N__18307),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__2697 (
            .O(N__18304),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    CEMux I__2696 (
            .O(N__18299),
            .I(N__18281));
    CEMux I__2695 (
            .O(N__18298),
            .I(N__18281));
    CEMux I__2694 (
            .O(N__18297),
            .I(N__18281));
    CEMux I__2693 (
            .O(N__18296),
            .I(N__18281));
    CEMux I__2692 (
            .O(N__18295),
            .I(N__18281));
    CEMux I__2691 (
            .O(N__18294),
            .I(N__18281));
    GlobalMux I__2690 (
            .O(N__18281),
            .I(N__18278));
    gio2CtrlBuf I__2689 (
            .O(N__18278),
            .I(\pid_alt.state_0_g_0 ));
    InMux I__2688 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__2687 (
            .O(N__18272),
            .I(N__18268));
    InMux I__2686 (
            .O(N__18271),
            .I(N__18265));
    Span4Mux_h I__2685 (
            .O(N__18268),
            .I(N__18259));
    LocalMux I__2684 (
            .O(N__18265),
            .I(N__18259));
    InMux I__2683 (
            .O(N__18264),
            .I(N__18256));
    Span4Mux_v I__2682 (
            .O(N__18259),
            .I(N__18253));
    LocalMux I__2681 (
            .O(N__18256),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    Odrv4 I__2680 (
            .O(N__18253),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    CascadeMux I__2679 (
            .O(N__18248),
            .I(N__18244));
    CascadeMux I__2678 (
            .O(N__18247),
            .I(N__18241));
    InMux I__2677 (
            .O(N__18244),
            .I(N__18237));
    InMux I__2676 (
            .O(N__18241),
            .I(N__18234));
    CascadeMux I__2675 (
            .O(N__18240),
            .I(N__18231));
    LocalMux I__2674 (
            .O(N__18237),
            .I(N__18228));
    LocalMux I__2673 (
            .O(N__18234),
            .I(N__18225));
    InMux I__2672 (
            .O(N__18231),
            .I(N__18222));
    Span4Mux_v I__2671 (
            .O(N__18228),
            .I(N__18219));
    Span4Mux_v I__2670 (
            .O(N__18225),
            .I(N__18214));
    LocalMux I__2669 (
            .O(N__18222),
            .I(N__18214));
    Span4Mux_v I__2668 (
            .O(N__18219),
            .I(N__18211));
    Span4Mux_v I__2667 (
            .O(N__18214),
            .I(N__18208));
    Odrv4 I__2666 (
            .O(N__18211),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    Odrv4 I__2665 (
            .O(N__18208),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__2664 (
            .O(N__18203),
            .I(N__18199));
    InMux I__2663 (
            .O(N__18202),
            .I(N__18196));
    LocalMux I__2662 (
            .O(N__18199),
            .I(N__18192));
    LocalMux I__2661 (
            .O(N__18196),
            .I(N__18189));
    InMux I__2660 (
            .O(N__18195),
            .I(N__18186));
    Span4Mux_v I__2659 (
            .O(N__18192),
            .I(N__18183));
    Odrv4 I__2658 (
            .O(N__18189),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    LocalMux I__2657 (
            .O(N__18186),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    Odrv4 I__2656 (
            .O(N__18183),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    InMux I__2655 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__2654 (
            .O(N__18173),
            .I(N__18170));
    Odrv4 I__2653 (
            .O(N__18170),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO ));
    InMux I__2652 (
            .O(N__18167),
            .I(N__18164));
    LocalMux I__2651 (
            .O(N__18164),
            .I(N__18161));
    Odrv4 I__2650 (
            .O(N__18161),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO ));
    CascadeMux I__2649 (
            .O(N__18158),
            .I(N__18154));
    InMux I__2648 (
            .O(N__18157),
            .I(N__18151));
    InMux I__2647 (
            .O(N__18154),
            .I(N__18148));
    LocalMux I__2646 (
            .O(N__18151),
            .I(N__18145));
    LocalMux I__2645 (
            .O(N__18148),
            .I(N__18140));
    Span4Mux_h I__2644 (
            .O(N__18145),
            .I(N__18137));
    CascadeMux I__2643 (
            .O(N__18144),
            .I(N__18134));
    InMux I__2642 (
            .O(N__18143),
            .I(N__18130));
    Span12Mux_v I__2641 (
            .O(N__18140),
            .I(N__18127));
    Span4Mux_v I__2640 (
            .O(N__18137),
            .I(N__18124));
    InMux I__2639 (
            .O(N__18134),
            .I(N__18119));
    InMux I__2638 (
            .O(N__18133),
            .I(N__18119));
    LocalMux I__2637 (
            .O(N__18130),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    Odrv12 I__2636 (
            .O(N__18127),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    Odrv4 I__2635 (
            .O(N__18124),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    LocalMux I__2634 (
            .O(N__18119),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__2633 (
            .O(N__18110),
            .I(N__18105));
    InMux I__2632 (
            .O(N__18109),
            .I(N__18100));
    InMux I__2631 (
            .O(N__18108),
            .I(N__18100));
    LocalMux I__2630 (
            .O(N__18105),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__2629 (
            .O(N__18100),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__2628 (
            .O(N__18095),
            .I(N__18092));
    LocalMux I__2627 (
            .O(N__18092),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO ));
    CascadeMux I__2626 (
            .O(N__18089),
            .I(N__18086));
    InMux I__2625 (
            .O(N__18086),
            .I(N__18081));
    InMux I__2624 (
            .O(N__18085),
            .I(N__18076));
    InMux I__2623 (
            .O(N__18084),
            .I(N__18076));
    LocalMux I__2622 (
            .O(N__18081),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    LocalMux I__2621 (
            .O(N__18076),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__2620 (
            .O(N__18071),
            .I(N__18068));
    LocalMux I__2619 (
            .O(N__18068),
            .I(N__18065));
    Span4Mux_v I__2618 (
            .O(N__18065),
            .I(N__18060));
    InMux I__2617 (
            .O(N__18064),
            .I(N__18055));
    InMux I__2616 (
            .O(N__18063),
            .I(N__18055));
    Odrv4 I__2615 (
            .O(N__18060),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    LocalMux I__2614 (
            .O(N__18055),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    CascadeMux I__2613 (
            .O(N__18050),
            .I(N__18044));
    CascadeMux I__2612 (
            .O(N__18049),
            .I(N__18041));
    InMux I__2611 (
            .O(N__18048),
            .I(N__18036));
    InMux I__2610 (
            .O(N__18047),
            .I(N__18036));
    InMux I__2609 (
            .O(N__18044),
            .I(N__18033));
    InMux I__2608 (
            .O(N__18041),
            .I(N__18030));
    LocalMux I__2607 (
            .O(N__18036),
            .I(N__18027));
    LocalMux I__2606 (
            .O(N__18033),
            .I(N__18022));
    LocalMux I__2605 (
            .O(N__18030),
            .I(N__18022));
    Span4Mux_h I__2604 (
            .O(N__18027),
            .I(N__18019));
    Odrv4 I__2603 (
            .O(N__18022),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    Odrv4 I__2602 (
            .O(N__18019),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    InMux I__2601 (
            .O(N__18014),
            .I(N__18011));
    LocalMux I__2600 (
            .O(N__18011),
            .I(N__18006));
    InMux I__2599 (
            .O(N__18010),
            .I(N__18001));
    InMux I__2598 (
            .O(N__18009),
            .I(N__18001));
    Odrv4 I__2597 (
            .O(N__18006),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__2596 (
            .O(N__18001),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__2595 (
            .O(N__17996),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__2594 (
            .O(N__17993),
            .I(N__17990));
    LocalMux I__2593 (
            .O(N__17990),
            .I(N__17987));
    Span4Mux_h I__2592 (
            .O(N__17987),
            .I(N__17982));
    InMux I__2591 (
            .O(N__17986),
            .I(N__17977));
    InMux I__2590 (
            .O(N__17985),
            .I(N__17977));
    Odrv4 I__2589 (
            .O(N__17982),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    LocalMux I__2588 (
            .O(N__17977),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    CascadeMux I__2587 (
            .O(N__17972),
            .I(N__17968));
    CascadeMux I__2586 (
            .O(N__17971),
            .I(N__17963));
    InMux I__2585 (
            .O(N__17968),
            .I(N__17960));
    InMux I__2584 (
            .O(N__17967),
            .I(N__17955));
    InMux I__2583 (
            .O(N__17966),
            .I(N__17955));
    InMux I__2582 (
            .O(N__17963),
            .I(N__17952));
    LocalMux I__2581 (
            .O(N__17960),
            .I(N__17949));
    LocalMux I__2580 (
            .O(N__17955),
            .I(N__17946));
    LocalMux I__2579 (
            .O(N__17952),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv4 I__2578 (
            .O(N__17949),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv4 I__2577 (
            .O(N__17946),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    InMux I__2576 (
            .O(N__17939),
            .I(N__17935));
    CascadeMux I__2575 (
            .O(N__17938),
            .I(N__17932));
    LocalMux I__2574 (
            .O(N__17935),
            .I(N__17928));
    InMux I__2573 (
            .O(N__17932),
            .I(N__17923));
    InMux I__2572 (
            .O(N__17931),
            .I(N__17923));
    Odrv4 I__2571 (
            .O(N__17928),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__2570 (
            .O(N__17923),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    InMux I__2569 (
            .O(N__17918),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__2568 (
            .O(N__17915),
            .I(N__17912));
    LocalMux I__2567 (
            .O(N__17912),
            .I(N__17909));
    Span4Mux_v I__2566 (
            .O(N__17909),
            .I(N__17904));
    InMux I__2565 (
            .O(N__17908),
            .I(N__17899));
    InMux I__2564 (
            .O(N__17907),
            .I(N__17899));
    Odrv4 I__2563 (
            .O(N__17904),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    LocalMux I__2562 (
            .O(N__17899),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    CascadeMux I__2561 (
            .O(N__17894),
            .I(N__17889));
    CascadeMux I__2560 (
            .O(N__17893),
            .I(N__17885));
    CascadeMux I__2559 (
            .O(N__17892),
            .I(N__17882));
    InMux I__2558 (
            .O(N__17889),
            .I(N__17879));
    InMux I__2557 (
            .O(N__17888),
            .I(N__17874));
    InMux I__2556 (
            .O(N__17885),
            .I(N__17874));
    InMux I__2555 (
            .O(N__17882),
            .I(N__17871));
    LocalMux I__2554 (
            .O(N__17879),
            .I(N__17868));
    LocalMux I__2553 (
            .O(N__17874),
            .I(N__17865));
    LocalMux I__2552 (
            .O(N__17871),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv4 I__2551 (
            .O(N__17868),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv4 I__2550 (
            .O(N__17865),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__2549 (
            .O(N__17858),
            .I(N__17854));
    CascadeMux I__2548 (
            .O(N__17857),
            .I(N__17850));
    LocalMux I__2547 (
            .O(N__17854),
            .I(N__17847));
    InMux I__2546 (
            .O(N__17853),
            .I(N__17842));
    InMux I__2545 (
            .O(N__17850),
            .I(N__17842));
    Odrv4 I__2544 (
            .O(N__17847),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__2543 (
            .O(N__17842),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__2542 (
            .O(N__17837),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__2541 (
            .O(N__17834),
            .I(N__17831));
    LocalMux I__2540 (
            .O(N__17831),
            .I(N__17828));
    Span4Mux_v I__2539 (
            .O(N__17828),
            .I(N__17823));
    InMux I__2538 (
            .O(N__17827),
            .I(N__17818));
    InMux I__2537 (
            .O(N__17826),
            .I(N__17818));
    Odrv4 I__2536 (
            .O(N__17823),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    LocalMux I__2535 (
            .O(N__17818),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    CascadeMux I__2534 (
            .O(N__17813),
            .I(N__17809));
    CascadeMux I__2533 (
            .O(N__17812),
            .I(N__17804));
    InMux I__2532 (
            .O(N__17809),
            .I(N__17801));
    InMux I__2531 (
            .O(N__17808),
            .I(N__17796));
    InMux I__2530 (
            .O(N__17807),
            .I(N__17796));
    InMux I__2529 (
            .O(N__17804),
            .I(N__17793));
    LocalMux I__2528 (
            .O(N__17801),
            .I(N__17790));
    LocalMux I__2527 (
            .O(N__17796),
            .I(N__17787));
    LocalMux I__2526 (
            .O(N__17793),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    Odrv12 I__2525 (
            .O(N__17790),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    Odrv12 I__2524 (
            .O(N__17787),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    CascadeMux I__2523 (
            .O(N__17780),
            .I(N__17777));
    InMux I__2522 (
            .O(N__17777),
            .I(N__17773));
    InMux I__2521 (
            .O(N__17776),
            .I(N__17770));
    LocalMux I__2520 (
            .O(N__17773),
            .I(N__17767));
    LocalMux I__2519 (
            .O(N__17770),
            .I(N__17763));
    Span4Mux_h I__2518 (
            .O(N__17767),
            .I(N__17760));
    InMux I__2517 (
            .O(N__17766),
            .I(N__17757));
    Odrv4 I__2516 (
            .O(N__17763),
            .I(\pid_alt.error_i_acumm7lto12 ));
    Odrv4 I__2515 (
            .O(N__17760),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__2514 (
            .O(N__17757),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__2513 (
            .O(N__17750),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__2512 (
            .O(N__17747),
            .I(N__17741));
    InMux I__2511 (
            .O(N__17746),
            .I(N__17741));
    LocalMux I__2510 (
            .O(N__17741),
            .I(N__17737));
    InMux I__2509 (
            .O(N__17740),
            .I(N__17734));
    Span4Mux_v I__2508 (
            .O(N__17737),
            .I(N__17731));
    LocalMux I__2507 (
            .O(N__17734),
            .I(N__17728));
    Span4Mux_v I__2506 (
            .O(N__17731),
            .I(N__17725));
    Odrv4 I__2505 (
            .O(N__17728),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    Odrv4 I__2504 (
            .O(N__17725),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CascadeMux I__2503 (
            .O(N__17720),
            .I(N__17717));
    InMux I__2502 (
            .O(N__17717),
            .I(N__17714));
    LocalMux I__2501 (
            .O(N__17714),
            .I(N__17711));
    Span4Mux_h I__2500 (
            .O(N__17711),
            .I(N__17706));
    InMux I__2499 (
            .O(N__17710),
            .I(N__17703));
    InMux I__2498 (
            .O(N__17709),
            .I(N__17700));
    Span4Mux_v I__2497 (
            .O(N__17706),
            .I(N__17697));
    LocalMux I__2496 (
            .O(N__17703),
            .I(N__17692));
    LocalMux I__2495 (
            .O(N__17700),
            .I(N__17692));
    Odrv4 I__2494 (
            .O(N__17697),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    Odrv4 I__2493 (
            .O(N__17692),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__2492 (
            .O(N__17687),
            .I(N__17678));
    InMux I__2491 (
            .O(N__17686),
            .I(N__17678));
    InMux I__2490 (
            .O(N__17685),
            .I(N__17678));
    LocalMux I__2489 (
            .O(N__17678),
            .I(N__17675));
    Odrv4 I__2488 (
            .O(N__17675),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__2487 (
            .O(N__17672),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__2486 (
            .O(N__17669),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__2485 (
            .O(N__17666),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__2484 (
            .O(N__17663),
            .I(bfn_3_15_0_));
    InMux I__2483 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__2482 (
            .O(N__17657),
            .I(N__17652));
    InMux I__2481 (
            .O(N__17656),
            .I(N__17647));
    InMux I__2480 (
            .O(N__17655),
            .I(N__17647));
    Span4Mux_h I__2479 (
            .O(N__17652),
            .I(N__17644));
    LocalMux I__2478 (
            .O(N__17647),
            .I(N__17641));
    Odrv4 I__2477 (
            .O(N__17644),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    Odrv12 I__2476 (
            .O(N__17641),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    CascadeMux I__2475 (
            .O(N__17636),
            .I(N__17633));
    InMux I__2474 (
            .O(N__17633),
            .I(N__17630));
    LocalMux I__2473 (
            .O(N__17630),
            .I(N__17626));
    CascadeMux I__2472 (
            .O(N__17629),
            .I(N__17623));
    Span4Mux_v I__2471 (
            .O(N__17626),
            .I(N__17619));
    InMux I__2470 (
            .O(N__17623),
            .I(N__17614));
    InMux I__2469 (
            .O(N__17622),
            .I(N__17614));
    Odrv4 I__2468 (
            .O(N__17619),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    LocalMux I__2467 (
            .O(N__17614),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    InMux I__2466 (
            .O(N__17609),
            .I(N__17606));
    LocalMux I__2465 (
            .O(N__17606),
            .I(N__17603));
    Span4Mux_s3_h I__2464 (
            .O(N__17603),
            .I(N__17599));
    InMux I__2463 (
            .O(N__17602),
            .I(N__17596));
    Odrv4 I__2462 (
            .O(N__17599),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__2461 (
            .O(N__17596),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    InMux I__2460 (
            .O(N__17591),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__2459 (
            .O(N__17588),
            .I(N__17583));
    InMux I__2458 (
            .O(N__17587),
            .I(N__17578));
    InMux I__2457 (
            .O(N__17586),
            .I(N__17578));
    LocalMux I__2456 (
            .O(N__17583),
            .I(N__17575));
    LocalMux I__2455 (
            .O(N__17578),
            .I(N__17572));
    Odrv12 I__2454 (
            .O(N__17575),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    Odrv4 I__2453 (
            .O(N__17572),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    CascadeMux I__2452 (
            .O(N__17567),
            .I(N__17564));
    InMux I__2451 (
            .O(N__17564),
            .I(N__17561));
    LocalMux I__2450 (
            .O(N__17561),
            .I(N__17557));
    CascadeMux I__2449 (
            .O(N__17560),
            .I(N__17554));
    Span4Mux_h I__2448 (
            .O(N__17557),
            .I(N__17550));
    InMux I__2447 (
            .O(N__17554),
            .I(N__17545));
    InMux I__2446 (
            .O(N__17553),
            .I(N__17545));
    Odrv4 I__2445 (
            .O(N__17550),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    LocalMux I__2444 (
            .O(N__17545),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    InMux I__2443 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__2442 (
            .O(N__17537),
            .I(N__17534));
    Span4Mux_v I__2441 (
            .O(N__17534),
            .I(N__17530));
    InMux I__2440 (
            .O(N__17533),
            .I(N__17527));
    Odrv4 I__2439 (
            .O(N__17530),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    LocalMux I__2438 (
            .O(N__17527),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    InMux I__2437 (
            .O(N__17522),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__2436 (
            .O(N__17519),
            .I(N__17516));
    LocalMux I__2435 (
            .O(N__17516),
            .I(N__17513));
    Span4Mux_v I__2434 (
            .O(N__17513),
            .I(N__17508));
    InMux I__2433 (
            .O(N__17512),
            .I(N__17503));
    InMux I__2432 (
            .O(N__17511),
            .I(N__17503));
    Odrv4 I__2431 (
            .O(N__17508),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    LocalMux I__2430 (
            .O(N__17503),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    CascadeMux I__2429 (
            .O(N__17498),
            .I(N__17494));
    CascadeMux I__2428 (
            .O(N__17497),
            .I(N__17491));
    InMux I__2427 (
            .O(N__17494),
            .I(N__17487));
    InMux I__2426 (
            .O(N__17491),
            .I(N__17482));
    InMux I__2425 (
            .O(N__17490),
            .I(N__17482));
    LocalMux I__2424 (
            .O(N__17487),
            .I(N__17479));
    LocalMux I__2423 (
            .O(N__17482),
            .I(N__17476));
    Odrv4 I__2422 (
            .O(N__17479),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    Odrv4 I__2421 (
            .O(N__17476),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    CascadeMux I__2420 (
            .O(N__17471),
            .I(N__17467));
    CascadeMux I__2419 (
            .O(N__17470),
            .I(N__17461));
    InMux I__2418 (
            .O(N__17467),
            .I(N__17456));
    InMux I__2417 (
            .O(N__17466),
            .I(N__17456));
    InMux I__2416 (
            .O(N__17465),
            .I(N__17453));
    InMux I__2415 (
            .O(N__17464),
            .I(N__17450));
    InMux I__2414 (
            .O(N__17461),
            .I(N__17447));
    LocalMux I__2413 (
            .O(N__17456),
            .I(N__17442));
    LocalMux I__2412 (
            .O(N__17453),
            .I(N__17442));
    LocalMux I__2411 (
            .O(N__17450),
            .I(N__17437));
    LocalMux I__2410 (
            .O(N__17447),
            .I(N__17437));
    Span4Mux_s3_h I__2409 (
            .O(N__17442),
            .I(N__17433));
    Span4Mux_s3_h I__2408 (
            .O(N__17437),
            .I(N__17430));
    InMux I__2407 (
            .O(N__17436),
            .I(N__17427));
    Odrv4 I__2406 (
            .O(N__17433),
            .I(\pid_alt.error_i_acumm7lto4 ));
    Odrv4 I__2405 (
            .O(N__17430),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__2404 (
            .O(N__17427),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__2403 (
            .O(N__17420),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__2402 (
            .O(N__17417),
            .I(N__17412));
    InMux I__2401 (
            .O(N__17416),
            .I(N__17408));
    CascadeMux I__2400 (
            .O(N__17415),
            .I(N__17405));
    LocalMux I__2399 (
            .O(N__17412),
            .I(N__17402));
    InMux I__2398 (
            .O(N__17411),
            .I(N__17399));
    LocalMux I__2397 (
            .O(N__17408),
            .I(N__17396));
    InMux I__2396 (
            .O(N__17405),
            .I(N__17393));
    Span4Mux_v I__2395 (
            .O(N__17402),
            .I(N__17390));
    LocalMux I__2394 (
            .O(N__17399),
            .I(N__17385));
    Span12Mux_s8_v I__2393 (
            .O(N__17396),
            .I(N__17385));
    LocalMux I__2392 (
            .O(N__17393),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    Odrv4 I__2391 (
            .O(N__17390),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    Odrv12 I__2390 (
            .O(N__17385),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    CascadeMux I__2389 (
            .O(N__17378),
            .I(N__17374));
    InMux I__2388 (
            .O(N__17377),
            .I(N__17370));
    InMux I__2387 (
            .O(N__17374),
            .I(N__17367));
    InMux I__2386 (
            .O(N__17373),
            .I(N__17364));
    LocalMux I__2385 (
            .O(N__17370),
            .I(N__17361));
    LocalMux I__2384 (
            .O(N__17367),
            .I(N__17358));
    LocalMux I__2383 (
            .O(N__17364),
            .I(N__17355));
    Span4Mux_v I__2382 (
            .O(N__17361),
            .I(N__17352));
    Odrv12 I__2381 (
            .O(N__17358),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    Odrv12 I__2380 (
            .O(N__17355),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    Odrv4 I__2379 (
            .O(N__17352),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__2378 (
            .O(N__17345),
            .I(N__17340));
    InMux I__2377 (
            .O(N__17344),
            .I(N__17337));
    InMux I__2376 (
            .O(N__17343),
            .I(N__17334));
    LocalMux I__2375 (
            .O(N__17340),
            .I(N__17329));
    LocalMux I__2374 (
            .O(N__17337),
            .I(N__17329));
    LocalMux I__2373 (
            .O(N__17334),
            .I(N__17326));
    Span4Mux_v I__2372 (
            .O(N__17329),
            .I(N__17321));
    Span4Mux_s3_h I__2371 (
            .O(N__17326),
            .I(N__17318));
    InMux I__2370 (
            .O(N__17325),
            .I(N__17313));
    InMux I__2369 (
            .O(N__17324),
            .I(N__17313));
    Odrv4 I__2368 (
            .O(N__17321),
            .I(\pid_alt.error_i_acumm7lto5 ));
    Odrv4 I__2367 (
            .O(N__17318),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__2366 (
            .O(N__17313),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__2365 (
            .O(N__17306),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__2364 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__2363 (
            .O(N__17300),
            .I(N__17297));
    Span4Mux_s3_h I__2362 (
            .O(N__17297),
            .I(N__17292));
    InMux I__2361 (
            .O(N__17296),
            .I(N__17287));
    InMux I__2360 (
            .O(N__17295),
            .I(N__17287));
    Odrv4 I__2359 (
            .O(N__17292),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__2358 (
            .O(N__17287),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__2357 (
            .O(N__17282),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__2356 (
            .O(N__17279),
            .I(N__17276));
    LocalMux I__2355 (
            .O(N__17276),
            .I(N__17272));
    CascadeMux I__2354 (
            .O(N__17275),
            .I(N__17269));
    Span4Mux_v I__2353 (
            .O(N__17272),
            .I(N__17265));
    InMux I__2352 (
            .O(N__17269),
            .I(N__17260));
    InMux I__2351 (
            .O(N__17268),
            .I(N__17260));
    Odrv4 I__2350 (
            .O(N__17265),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__2349 (
            .O(N__17260),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    InMux I__2348 (
            .O(N__17255),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__2347 (
            .O(N__17252),
            .I(N__17249));
    LocalMux I__2346 (
            .O(N__17249),
            .I(N__17246));
    Span4Mux_v I__2345 (
            .O(N__17246),
            .I(N__17241));
    InMux I__2344 (
            .O(N__17245),
            .I(N__17236));
    InMux I__2343 (
            .O(N__17244),
            .I(N__17236));
    Odrv4 I__2342 (
            .O(N__17241),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    LocalMux I__2341 (
            .O(N__17236),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    CascadeMux I__2340 (
            .O(N__17231),
            .I(N__17227));
    CascadeMux I__2339 (
            .O(N__17230),
            .I(N__17222));
    InMux I__2338 (
            .O(N__17227),
            .I(N__17217));
    InMux I__2337 (
            .O(N__17226),
            .I(N__17217));
    CascadeMux I__2336 (
            .O(N__17225),
            .I(N__17214));
    InMux I__2335 (
            .O(N__17222),
            .I(N__17211));
    LocalMux I__2334 (
            .O(N__17217),
            .I(N__17208));
    InMux I__2333 (
            .O(N__17214),
            .I(N__17205));
    LocalMux I__2332 (
            .O(N__17211),
            .I(N__17202));
    Span4Mux_h I__2331 (
            .O(N__17208),
            .I(N__17199));
    LocalMux I__2330 (
            .O(N__17205),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    Odrv12 I__2329 (
            .O(N__17202),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    Odrv4 I__2328 (
            .O(N__17199),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    InMux I__2327 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__2326 (
            .O(N__17189),
            .I(N__17184));
    InMux I__2325 (
            .O(N__17188),
            .I(N__17179));
    InMux I__2324 (
            .O(N__17187),
            .I(N__17179));
    Odrv4 I__2323 (
            .O(N__17184),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__2322 (
            .O(N__17179),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    InMux I__2321 (
            .O(N__17174),
            .I(bfn_3_14_0_));
    InMux I__2320 (
            .O(N__17171),
            .I(N__17168));
    LocalMux I__2319 (
            .O(N__17168),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__2318 (
            .O(N__17165),
            .I(N__17162));
    LocalMux I__2317 (
            .O(N__17162),
            .I(drone_altitude_12));
    InMux I__2316 (
            .O(N__17159),
            .I(N__17156));
    LocalMux I__2315 (
            .O(N__17156),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__2314 (
            .O(N__17153),
            .I(N__17150));
    LocalMux I__2313 (
            .O(N__17150),
            .I(drone_altitude_13));
    InMux I__2312 (
            .O(N__17147),
            .I(N__17144));
    LocalMux I__2311 (
            .O(N__17144),
            .I(\pid_alt.error_axbZ0Z_14 ));
    CascadeMux I__2310 (
            .O(N__17141),
            .I(N__17138));
    InMux I__2309 (
            .O(N__17138),
            .I(N__17135));
    LocalMux I__2308 (
            .O(N__17135),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__2307 (
            .O(N__17132),
            .I(N__17129));
    LocalMux I__2306 (
            .O(N__17129),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__2305 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__2304 (
            .O(N__17123),
            .I(N__17120));
    Span4Mux_h I__2303 (
            .O(N__17120),
            .I(N__17115));
    InMux I__2302 (
            .O(N__17119),
            .I(N__17110));
    InMux I__2301 (
            .O(N__17118),
            .I(N__17110));
    Odrv4 I__2300 (
            .O(N__17115),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    LocalMux I__2299 (
            .O(N__17110),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    CascadeMux I__2298 (
            .O(N__17105),
            .I(N__17102));
    InMux I__2297 (
            .O(N__17102),
            .I(N__17097));
    InMux I__2296 (
            .O(N__17101),
            .I(N__17092));
    InMux I__2295 (
            .O(N__17100),
            .I(N__17092));
    LocalMux I__2294 (
            .O(N__17097),
            .I(N__17089));
    LocalMux I__2293 (
            .O(N__17092),
            .I(N__17086));
    Odrv4 I__2292 (
            .O(N__17089),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    Odrv12 I__2291 (
            .O(N__17086),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    CascadeMux I__2290 (
            .O(N__17081),
            .I(N__17078));
    InMux I__2289 (
            .O(N__17078),
            .I(N__17075));
    LocalMux I__2288 (
            .O(N__17075),
            .I(N__17072));
    Span4Mux_v I__2287 (
            .O(N__17072),
            .I(N__17069));
    Span4Mux_s1_h I__2286 (
            .O(N__17069),
            .I(N__17065));
    InMux I__2285 (
            .O(N__17068),
            .I(N__17062));
    Odrv4 I__2284 (
            .O(N__17065),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__2283 (
            .O(N__17062),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    InMux I__2282 (
            .O(N__17057),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    CascadeMux I__2281 (
            .O(N__17054),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    CascadeMux I__2280 (
            .O(N__17051),
            .I(N__17047));
    InMux I__2279 (
            .O(N__17050),
            .I(N__17044));
    InMux I__2278 (
            .O(N__17047),
            .I(N__17041));
    LocalMux I__2277 (
            .O(N__17044),
            .I(alt_command_0));
    LocalMux I__2276 (
            .O(N__17041),
            .I(alt_command_0));
    CascadeMux I__2275 (
            .O(N__17036),
            .I(N__17033));
    InMux I__2274 (
            .O(N__17033),
            .I(N__17030));
    LocalMux I__2273 (
            .O(N__17030),
            .I(drone_altitude_i_7));
    InMux I__2272 (
            .O(N__17027),
            .I(N__17024));
    LocalMux I__2271 (
            .O(N__17024),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    InMux I__2270 (
            .O(N__17021),
            .I(N__17018));
    LocalMux I__2269 (
            .O(N__17018),
            .I(drone_altitude_i_8));
    InMux I__2268 (
            .O(N__17015),
            .I(N__17012));
    LocalMux I__2267 (
            .O(N__17012),
            .I(drone_altitude_i_9));
    InMux I__2266 (
            .O(N__17009),
            .I(N__17006));
    LocalMux I__2265 (
            .O(N__17006),
            .I(drone_altitude_i_10));
    InMux I__2264 (
            .O(N__17003),
            .I(N__17000));
    LocalMux I__2263 (
            .O(N__17000),
            .I(drone_altitude_i_11));
    CascadeMux I__2262 (
            .O(N__16997),
            .I(N__16994));
    InMux I__2261 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__2260 (
            .O(N__16991),
            .I(\pid_alt.error_axbZ0Z_1 ));
    InMux I__2259 (
            .O(N__16988),
            .I(N__16985));
    LocalMux I__2258 (
            .O(N__16985),
            .I(drone_altitude_1));
    InMux I__2257 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__2256 (
            .O(N__16979),
            .I(N__16976));
    Span4Mux_s3_h I__2255 (
            .O(N__16976),
            .I(N__16973));
    Odrv4 I__2254 (
            .O(N__16973),
            .I(alt_kp_6));
    InMux I__2253 (
            .O(N__16970),
            .I(N__16967));
    LocalMux I__2252 (
            .O(N__16967),
            .I(N__16964));
    Span4Mux_s3_h I__2251 (
            .O(N__16964),
            .I(N__16961));
    Odrv4 I__2250 (
            .O(N__16961),
            .I(alt_kp_5));
    InMux I__2249 (
            .O(N__16958),
            .I(N__16955));
    LocalMux I__2248 (
            .O(N__16955),
            .I(N__16952));
    Span4Mux_s3_h I__2247 (
            .O(N__16952),
            .I(N__16949));
    Odrv4 I__2246 (
            .O(N__16949),
            .I(alt_kp_1));
    InMux I__2245 (
            .O(N__16946),
            .I(N__16943));
    LocalMux I__2244 (
            .O(N__16943),
            .I(N__16940));
    Odrv12 I__2243 (
            .O(N__16940),
            .I(alt_kp_0));
    InMux I__2242 (
            .O(N__16937),
            .I(N__16934));
    LocalMux I__2241 (
            .O(N__16934),
            .I(N__16931));
    Span4Mux_s3_h I__2240 (
            .O(N__16931),
            .I(N__16928));
    Odrv4 I__2239 (
            .O(N__16928),
            .I(drone_altitude_15));
    CascadeMux I__2238 (
            .O(N__16925),
            .I(N__16921));
    InMux I__2237 (
            .O(N__16924),
            .I(N__16918));
    InMux I__2236 (
            .O(N__16921),
            .I(N__16915));
    LocalMux I__2235 (
            .O(N__16918),
            .I(alt_command_2));
    LocalMux I__2234 (
            .O(N__16915),
            .I(alt_command_2));
    InMux I__2233 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__2232 (
            .O(N__16907),
            .I(N__16903));
    InMux I__2231 (
            .O(N__16906),
            .I(N__16900));
    Span4Mux_h I__2230 (
            .O(N__16903),
            .I(N__16897));
    LocalMux I__2229 (
            .O(N__16900),
            .I(alt_command_3));
    Odrv4 I__2228 (
            .O(N__16897),
            .I(alt_command_3));
    CascadeMux I__2227 (
            .O(N__16892),
            .I(N__16888));
    InMux I__2226 (
            .O(N__16891),
            .I(N__16885));
    InMux I__2225 (
            .O(N__16888),
            .I(N__16882));
    LocalMux I__2224 (
            .O(N__16885),
            .I(alt_command_1));
    LocalMux I__2223 (
            .O(N__16882),
            .I(alt_command_1));
    CascadeMux I__2222 (
            .O(N__16877),
            .I(\Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ));
    CascadeMux I__2221 (
            .O(N__16874),
            .I(N__16870));
    CascadeMux I__2220 (
            .O(N__16873),
            .I(N__16867));
    InMux I__2219 (
            .O(N__16870),
            .I(N__16859));
    InMux I__2218 (
            .O(N__16867),
            .I(N__16859));
    InMux I__2217 (
            .O(N__16866),
            .I(N__16859));
    LocalMux I__2216 (
            .O(N__16859),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    InMux I__2215 (
            .O(N__16856),
            .I(N__16853));
    LocalMux I__2214 (
            .O(N__16853),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ));
    CascadeMux I__2213 (
            .O(N__16850),
            .I(N__16847));
    InMux I__2212 (
            .O(N__16847),
            .I(N__16844));
    LocalMux I__2211 (
            .O(N__16844),
            .I(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ));
    InMux I__2210 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__2209 (
            .O(N__16838),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__2208 (
            .O(N__16835),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__2207 (
            .O(N__16832),
            .I(N__16829));
    LocalMux I__2206 (
            .O(N__16829),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__2205 (
            .O(N__16826),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__2204 (
            .O(N__16823),
            .I(N__16820));
    LocalMux I__2203 (
            .O(N__16820),
            .I(N__16817));
    Odrv4 I__2202 (
            .O(N__16817),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__2201 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__2200 (
            .O(N__16811),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__2199 (
            .O(N__16808),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__2198 (
            .O(N__16805),
            .I(bfn_2_30_0_));
    InMux I__2197 (
            .O(N__16802),
            .I(N__16799));
    LocalMux I__2196 (
            .O(N__16799),
            .I(N__16796));
    Odrv4 I__2195 (
            .O(N__16796),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__2194 (
            .O(N__16793),
            .I(N__16790));
    LocalMux I__2193 (
            .O(N__16790),
            .I(N__16787));
    Odrv4 I__2192 (
            .O(N__16787),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__2191 (
            .O(N__16784),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__2190 (
            .O(N__16781),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__2189 (
            .O(N__16778),
            .I(N__16775));
    LocalMux I__2188 (
            .O(N__16775),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__2187 (
            .O(N__16772),
            .I(N__16769));
    LocalMux I__2186 (
            .O(N__16769),
            .I(N__16766));
    Span4Mux_s3_h I__2185 (
            .O(N__16766),
            .I(N__16763));
    Odrv4 I__2184 (
            .O(N__16763),
            .I(alt_kp_3));
    InMux I__2183 (
            .O(N__16760),
            .I(N__16757));
    LocalMux I__2182 (
            .O(N__16757),
            .I(N__16754));
    Span4Mux_s3_v I__2181 (
            .O(N__16754),
            .I(N__16751));
    Odrv4 I__2180 (
            .O(N__16751),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__2179 (
            .O(N__16748),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__2178 (
            .O(N__16745),
            .I(N__16742));
    LocalMux I__2177 (
            .O(N__16742),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ));
    InMux I__2176 (
            .O(N__16739),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__2175 (
            .O(N__16736),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__2174 (
            .O(N__16733),
            .I(N__16730));
    LocalMux I__2173 (
            .O(N__16730),
            .I(N__16727));
    Odrv4 I__2172 (
            .O(N__16727),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__2171 (
            .O(N__16724),
            .I(bfn_2_29_0_));
    InMux I__2170 (
            .O(N__16721),
            .I(N__16718));
    LocalMux I__2169 (
            .O(N__16718),
            .I(N__16715));
    Span4Mux_s2_v I__2168 (
            .O(N__16715),
            .I(N__16712));
    Odrv4 I__2167 (
            .O(N__16712),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__2166 (
            .O(N__16709),
            .I(N__16706));
    LocalMux I__2165 (
            .O(N__16706),
            .I(N__16703));
    Odrv4 I__2164 (
            .O(N__16703),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__2163 (
            .O(N__16700),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__2162 (
            .O(N__16697),
            .I(N__16694));
    LocalMux I__2161 (
            .O(N__16694),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__2160 (
            .O(N__16691),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__2159 (
            .O(N__16688),
            .I(N__16685));
    LocalMux I__2158 (
            .O(N__16685),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__2157 (
            .O(N__16682),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__2156 (
            .O(N__16679),
            .I(N__16676));
    LocalMux I__2155 (
            .O(N__16676),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__2154 (
            .O(N__16673),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__2153 (
            .O(N__16670),
            .I(N__16667));
    LocalMux I__2152 (
            .O(N__16667),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__2151 (
            .O(N__16664),
            .I(N__16661));
    LocalMux I__2150 (
            .O(N__16661),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__2149 (
            .O(N__16658),
            .I(N__16655));
    LocalMux I__2148 (
            .O(N__16655),
            .I(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ));
    CascadeMux I__2147 (
            .O(N__16652),
            .I(N__16649));
    InMux I__2146 (
            .O(N__16649),
            .I(N__16646));
    LocalMux I__2145 (
            .O(N__16646),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__2144 (
            .O(N__16643),
            .I(N__16640));
    LocalMux I__2143 (
            .O(N__16640),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__2142 (
            .O(N__16637),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__2141 (
            .O(N__16634),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__2140 (
            .O(N__16631),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__2139 (
            .O(N__16628),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__2138 (
            .O(N__16625),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__2137 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__2136 (
            .O(N__16619),
            .I(N__16616));
    Span4Mux_s2_v I__2135 (
            .O(N__16616),
            .I(N__16613));
    Odrv4 I__2134 (
            .O(N__16613),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__2133 (
            .O(N__16610),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__2132 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__2131 (
            .O(N__16604),
            .I(N__16600));
    InMux I__2130 (
            .O(N__16603),
            .I(N__16597));
    Span4Mux_v I__2129 (
            .O(N__16600),
            .I(N__16592));
    LocalMux I__2128 (
            .O(N__16597),
            .I(N__16592));
    Span4Mux_v I__2127 (
            .O(N__16592),
            .I(N__16589));
    Odrv4 I__2126 (
            .O(N__16589),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    CascadeMux I__2125 (
            .O(N__16586),
            .I(N__16583));
    InMux I__2124 (
            .O(N__16583),
            .I(N__16580));
    LocalMux I__2123 (
            .O(N__16580),
            .I(N__16577));
    Odrv4 I__2122 (
            .O(N__16577),
            .I(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ));
    InMux I__2121 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__2120 (
            .O(N__16571),
            .I(N__16568));
    Span4Mux_s1_v I__2119 (
            .O(N__16568),
            .I(N__16565));
    Odrv4 I__2118 (
            .O(N__16565),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__2117 (
            .O(N__16562),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__2116 (
            .O(N__16559),
            .I(N__16556));
    LocalMux I__2115 (
            .O(N__16556),
            .I(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ));
    CascadeMux I__2114 (
            .O(N__16553),
            .I(N__16549));
    InMux I__2113 (
            .O(N__16552),
            .I(N__16546));
    InMux I__2112 (
            .O(N__16549),
            .I(N__16543));
    LocalMux I__2111 (
            .O(N__16546),
            .I(N__16538));
    LocalMux I__2110 (
            .O(N__16543),
            .I(N__16538));
    Span4Mux_v I__2109 (
            .O(N__16538),
            .I(N__16535));
    Odrv4 I__2108 (
            .O(N__16535),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    CascadeMux I__2107 (
            .O(N__16532),
            .I(N__16529));
    InMux I__2106 (
            .O(N__16529),
            .I(N__16526));
    LocalMux I__2105 (
            .O(N__16526),
            .I(N__16523));
    Odrv4 I__2104 (
            .O(N__16523),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__2103 (
            .O(N__16520),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__2102 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__2101 (
            .O(N__16514),
            .I(N__16511));
    Span4Mux_h I__2100 (
            .O(N__16511),
            .I(N__16508));
    Odrv4 I__2099 (
            .O(N__16508),
            .I(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ));
    CascadeMux I__2098 (
            .O(N__16505),
            .I(N__16502));
    InMux I__2097 (
            .O(N__16502),
            .I(N__16499));
    LocalMux I__2096 (
            .O(N__16499),
            .I(N__16496));
    Span4Mux_h I__2095 (
            .O(N__16496),
            .I(N__16493));
    Odrv4 I__2094 (
            .O(N__16493),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ));
    InMux I__2093 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__2092 (
            .O(N__16487),
            .I(N__16484));
    Span4Mux_s1_v I__2091 (
            .O(N__16484),
            .I(N__16481));
    Odrv4 I__2090 (
            .O(N__16481),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__2089 (
            .O(N__16478),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__2088 (
            .O(N__16475),
            .I(bfn_2_27_0_));
    CascadeMux I__2087 (
            .O(N__16472),
            .I(N__16469));
    InMux I__2086 (
            .O(N__16469),
            .I(N__16466));
    LocalMux I__2085 (
            .O(N__16466),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__2084 (
            .O(N__16463),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__2083 (
            .O(N__16460),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    CascadeMux I__2082 (
            .O(N__16457),
            .I(N__16454));
    InMux I__2081 (
            .O(N__16454),
            .I(N__16451));
    LocalMux I__2080 (
            .O(N__16451),
            .I(N__16448));
    Odrv4 I__2079 (
            .O(N__16448),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__2078 (
            .O(N__16445),
            .I(N__16442));
    LocalMux I__2077 (
            .O(N__16442),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__2076 (
            .O(N__16439),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__2075 (
            .O(N__16436),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__2074 (
            .O(N__16433),
            .I(N__16429));
    InMux I__2073 (
            .O(N__16432),
            .I(N__16426));
    LocalMux I__2072 (
            .O(N__16429),
            .I(N__16423));
    LocalMux I__2071 (
            .O(N__16426),
            .I(N__16420));
    Span4Mux_h I__2070 (
            .O(N__16423),
            .I(N__16417));
    Odrv4 I__2069 (
            .O(N__16420),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    Odrv4 I__2068 (
            .O(N__16417),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    CascadeMux I__2067 (
            .O(N__16412),
            .I(N__16409));
    InMux I__2066 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2065 (
            .O(N__16406),
            .I(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ));
    InMux I__2064 (
            .O(N__16403),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    CascadeMux I__2063 (
            .O(N__16400),
            .I(N__16397));
    InMux I__2062 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__2061 (
            .O(N__16394),
            .I(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ));
    InMux I__2060 (
            .O(N__16391),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    CascadeMux I__2059 (
            .O(N__16388),
            .I(N__16385));
    InMux I__2058 (
            .O(N__16385),
            .I(N__16382));
    LocalMux I__2057 (
            .O(N__16382),
            .I(N__16379));
    Odrv4 I__2056 (
            .O(N__16379),
            .I(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ));
    InMux I__2055 (
            .O(N__16376),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__2054 (
            .O(N__16373),
            .I(bfn_2_26_0_));
    CascadeMux I__2053 (
            .O(N__16370),
            .I(N__16367));
    InMux I__2052 (
            .O(N__16367),
            .I(N__16364));
    LocalMux I__2051 (
            .O(N__16364),
            .I(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ));
    CascadeMux I__2050 (
            .O(N__16361),
            .I(N__16358));
    InMux I__2049 (
            .O(N__16358),
            .I(N__16355));
    LocalMux I__2048 (
            .O(N__16355),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__2047 (
            .O(N__16352),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    CascadeMux I__2046 (
            .O(N__16349),
            .I(N__16346));
    InMux I__2045 (
            .O(N__16346),
            .I(N__16343));
    LocalMux I__2044 (
            .O(N__16343),
            .I(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ));
    InMux I__2043 (
            .O(N__16340),
            .I(N__16337));
    LocalMux I__2042 (
            .O(N__16337),
            .I(N__16334));
    Odrv4 I__2041 (
            .O(N__16334),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__2040 (
            .O(N__16331),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    CascadeMux I__2039 (
            .O(N__16328),
            .I(N__16325));
    InMux I__2038 (
            .O(N__16325),
            .I(N__16322));
    LocalMux I__2037 (
            .O(N__16322),
            .I(N__16319));
    Odrv12 I__2036 (
            .O(N__16319),
            .I(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ));
    CascadeMux I__2035 (
            .O(N__16316),
            .I(N__16313));
    InMux I__2034 (
            .O(N__16313),
            .I(N__16310));
    LocalMux I__2033 (
            .O(N__16310),
            .I(N__16307));
    Odrv4 I__2032 (
            .O(N__16307),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    CascadeMux I__2031 (
            .O(N__16304),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ));
    CascadeMux I__2030 (
            .O(N__16301),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    InMux I__2029 (
            .O(N__16298),
            .I(N__16295));
    LocalMux I__2028 (
            .O(N__16295),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    InMux I__2027 (
            .O(N__16292),
            .I(N__16289));
    LocalMux I__2026 (
            .O(N__16289),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13 ));
    InMux I__2025 (
            .O(N__16286),
            .I(N__16282));
    InMux I__2024 (
            .O(N__16285),
            .I(N__16279));
    LocalMux I__2023 (
            .O(N__16282),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    LocalMux I__2022 (
            .O(N__16279),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__2021 (
            .O(N__16274),
            .I(N__16270));
    InMux I__2020 (
            .O(N__16273),
            .I(N__16267));
    LocalMux I__2019 (
            .O(N__16270),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    LocalMux I__2018 (
            .O(N__16267),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    InMux I__2017 (
            .O(N__16262),
            .I(N__16259));
    LocalMux I__2016 (
            .O(N__16259),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5 ));
    InMux I__2015 (
            .O(N__16256),
            .I(N__16253));
    LocalMux I__2014 (
            .O(N__16253),
            .I(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ));
    InMux I__2013 (
            .O(N__16250),
            .I(N__16247));
    LocalMux I__2012 (
            .O(N__16247),
            .I(N__16244));
    Span4Mux_s3_v I__2011 (
            .O(N__16244),
            .I(N__16241));
    Odrv4 I__2010 (
            .O(N__16241),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__2009 (
            .O(N__16238),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__2008 (
            .O(N__16235),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    CascadeMux I__2007 (
            .O(N__16232),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    InMux I__2006 (
            .O(N__16229),
            .I(N__16226));
    LocalMux I__2005 (
            .O(N__16226),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    CascadeMux I__2004 (
            .O(N__16223),
            .I(\ppm_encoder_1.N_299_cascade_ ));
    InMux I__2003 (
            .O(N__16220),
            .I(N__16211));
    InMux I__2002 (
            .O(N__16219),
            .I(N__16211));
    InMux I__2001 (
            .O(N__16218),
            .I(N__16211));
    LocalMux I__2000 (
            .O(N__16211),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__1999 (
            .O(N__16208),
            .I(N__16199));
    InMux I__1998 (
            .O(N__16207),
            .I(N__16199));
    InMux I__1997 (
            .O(N__16206),
            .I(N__16199));
    LocalMux I__1996 (
            .O(N__16199),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__1995 (
            .O(N__16196),
            .I(N__16193));
    LocalMux I__1994 (
            .O(N__16193),
            .I(N__16190));
    Odrv4 I__1993 (
            .O(N__16190),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    CascadeMux I__1992 (
            .O(N__16187),
            .I(N__16184));
    InMux I__1991 (
            .O(N__16184),
            .I(N__16179));
    InMux I__1990 (
            .O(N__16183),
            .I(N__16176));
    InMux I__1989 (
            .O(N__16182),
            .I(N__16173));
    LocalMux I__1988 (
            .O(N__16179),
            .I(N__16168));
    LocalMux I__1987 (
            .O(N__16176),
            .I(N__16168));
    LocalMux I__1986 (
            .O(N__16173),
            .I(N__16165));
    Odrv4 I__1985 (
            .O(N__16168),
            .I(throttle_command_7));
    Odrv4 I__1984 (
            .O(N__16165),
            .I(throttle_command_7));
    InMux I__1983 (
            .O(N__16160),
            .I(N__16151));
    InMux I__1982 (
            .O(N__16159),
            .I(N__16151));
    InMux I__1981 (
            .O(N__16158),
            .I(N__16151));
    LocalMux I__1980 (
            .O(N__16151),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    CascadeMux I__1979 (
            .O(N__16148),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ));
    InMux I__1978 (
            .O(N__16145),
            .I(N__16142));
    LocalMux I__1977 (
            .O(N__16142),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    CascadeMux I__1976 (
            .O(N__16139),
            .I(\ppm_encoder_1.N_303_cascade_ ));
    InMux I__1975 (
            .O(N__16136),
            .I(N__16127));
    InMux I__1974 (
            .O(N__16135),
            .I(N__16127));
    InMux I__1973 (
            .O(N__16134),
            .I(N__16127));
    LocalMux I__1972 (
            .O(N__16127),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__1971 (
            .O(N__16124),
            .I(N__16115));
    InMux I__1970 (
            .O(N__16123),
            .I(N__16115));
    InMux I__1969 (
            .O(N__16122),
            .I(N__16115));
    LocalMux I__1968 (
            .O(N__16115),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__1967 (
            .O(N__16112),
            .I(N__16109));
    LocalMux I__1966 (
            .O(N__16109),
            .I(N__16104));
    InMux I__1965 (
            .O(N__16108),
            .I(N__16101));
    InMux I__1964 (
            .O(N__16107),
            .I(N__16098));
    Span4Mux_h I__1963 (
            .O(N__16104),
            .I(N__16095));
    LocalMux I__1962 (
            .O(N__16101),
            .I(N__16092));
    LocalMux I__1961 (
            .O(N__16098),
            .I(throttle_command_11));
    Odrv4 I__1960 (
            .O(N__16095),
            .I(throttle_command_11));
    Odrv12 I__1959 (
            .O(N__16092),
            .I(throttle_command_11));
    CascadeMux I__1958 (
            .O(N__16085),
            .I(N__16082));
    InMux I__1957 (
            .O(N__16082),
            .I(N__16079));
    LocalMux I__1956 (
            .O(N__16079),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__1955 (
            .O(N__16076),
            .I(N__16067));
    InMux I__1954 (
            .O(N__16075),
            .I(N__16067));
    InMux I__1953 (
            .O(N__16074),
            .I(N__16067));
    LocalMux I__1952 (
            .O(N__16067),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    InMux I__1951 (
            .O(N__16064),
            .I(N__16061));
    LocalMux I__1950 (
            .O(N__16061),
            .I(N__16058));
    Odrv4 I__1949 (
            .O(N__16058),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    InMux I__1948 (
            .O(N__16055),
            .I(N__16052));
    LocalMux I__1947 (
            .O(N__16052),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    CascadeMux I__1946 (
            .O(N__16049),
            .I(N__16046));
    InMux I__1945 (
            .O(N__16046),
            .I(N__16043));
    LocalMux I__1944 (
            .O(N__16043),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    InMux I__1943 (
            .O(N__16040),
            .I(N__16037));
    LocalMux I__1942 (
            .O(N__16037),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    InMux I__1941 (
            .O(N__16034),
            .I(N__16031));
    LocalMux I__1940 (
            .O(N__16031),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__1939 (
            .O(N__16028),
            .I(N__16025));
    LocalMux I__1938 (
            .O(N__16025),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    CascadeMux I__1937 (
            .O(N__16022),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_ ));
    CascadeMux I__1936 (
            .O(N__16019),
            .I(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_ ));
    InMux I__1935 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__1934 (
            .O(N__16013),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__1933 (
            .O(N__16010),
            .I(N__16007));
    LocalMux I__1932 (
            .O(N__16007),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__1931 (
            .O(N__16004),
            .I(N__16001));
    LocalMux I__1930 (
            .O(N__16001),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_3 ));
    CascadeMux I__1929 (
            .O(N__15998),
            .I(N__15995));
    InMux I__1928 (
            .O(N__15995),
            .I(N__15992));
    LocalMux I__1927 (
            .O(N__15992),
            .I(\pid_alt.source_pid_9_0_0_4 ));
    InMux I__1926 (
            .O(N__15989),
            .I(N__15986));
    LocalMux I__1925 (
            .O(N__15986),
            .I(N__15982));
    InMux I__1924 (
            .O(N__15985),
            .I(N__15979));
    Odrv4 I__1923 (
            .O(N__15982),
            .I(throttle_command_5));
    LocalMux I__1922 (
            .O(N__15979),
            .I(throttle_command_5));
    InMux I__1921 (
            .O(N__15974),
            .I(N__15971));
    LocalMux I__1920 (
            .O(N__15971),
            .I(N__15968));
    Span12Mux_v I__1919 (
            .O(N__15968),
            .I(N__15965));
    Odrv12 I__1918 (
            .O(N__15965),
            .I(\pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14 ));
    CascadeMux I__1917 (
            .O(N__15962),
            .I(N__15959));
    InMux I__1916 (
            .O(N__15959),
            .I(N__15956));
    LocalMux I__1915 (
            .O(N__15956),
            .I(N__15953));
    Span12Mux_h I__1914 (
            .O(N__15953),
            .I(N__15950));
    Span12Mux_v I__1913 (
            .O(N__15950),
            .I(N__15947));
    Odrv12 I__1912 (
            .O(N__15947),
            .I(\pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14 ));
    InMux I__1911 (
            .O(N__15944),
            .I(bfn_2_19_0_));
    InMux I__1910 (
            .O(N__15941),
            .I(N__15938));
    LocalMux I__1909 (
            .O(N__15938),
            .I(N__15935));
    Span12Mux_s3_h I__1908 (
            .O(N__15935),
            .I(N__15932));
    Span12Mux_v I__1907 (
            .O(N__15932),
            .I(N__15929));
    Odrv12 I__1906 (
            .O(N__15929),
            .I(\pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15 ));
    CascadeMux I__1905 (
            .O(N__15926),
            .I(N__15923));
    InMux I__1904 (
            .O(N__15923),
            .I(N__15920));
    LocalMux I__1903 (
            .O(N__15920),
            .I(N__15917));
    Span12Mux_v I__1902 (
            .O(N__15917),
            .I(N__15914));
    Odrv12 I__1901 (
            .O(N__15914),
            .I(\pid_alt.error_p_reg_esr_RNIKU581Z0Z_15 ));
    InMux I__1900 (
            .O(N__15911),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__1899 (
            .O(N__15908),
            .I(N__15905));
    LocalMux I__1898 (
            .O(N__15905),
            .I(N__15902));
    Span4Mux_v I__1897 (
            .O(N__15902),
            .I(N__15899));
    Odrv4 I__1896 (
            .O(N__15899),
            .I(\pid_alt.error_p_reg_esr_RNIO2681Z0Z_16 ));
    InMux I__1895 (
            .O(N__15896),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__1894 (
            .O(N__15893),
            .I(N__15890));
    LocalMux I__1893 (
            .O(N__15890),
            .I(N__15887));
    Span4Mux_h I__1892 (
            .O(N__15887),
            .I(N__15884));
    Span4Mux_v I__1891 (
            .O(N__15884),
            .I(N__15881));
    Odrv4 I__1890 (
            .O(N__15881),
            .I(\pid_alt.error_p_reg_esr_RNID23KZ0Z_17 ));
    CascadeMux I__1889 (
            .O(N__15878),
            .I(N__15875));
    InMux I__1888 (
            .O(N__15875),
            .I(N__15872));
    LocalMux I__1887 (
            .O(N__15872),
            .I(N__15869));
    Odrv4 I__1886 (
            .O(N__15869),
            .I(\pid_alt.error_p_reg_esr_RNIS6681Z0Z_17 ));
    InMux I__1885 (
            .O(N__15866),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    CascadeMux I__1884 (
            .O(N__15863),
            .I(N__15860));
    InMux I__1883 (
            .O(N__15860),
            .I(N__15857));
    LocalMux I__1882 (
            .O(N__15857),
            .I(N__15854));
    Odrv4 I__1881 (
            .O(N__15854),
            .I(\pid_alt.error_p_reg_esr_RNI0B681Z0Z_18 ));
    InMux I__1880 (
            .O(N__15851),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__1879 (
            .O(N__15848),
            .I(N__15845));
    LocalMux I__1878 (
            .O(N__15845),
            .I(N__15842));
    Span4Mux_v I__1877 (
            .O(N__15842),
            .I(N__15839));
    Odrv4 I__1876 (
            .O(N__15839),
            .I(\pid_alt.error_p_reg_esr_RNIIU781Z0Z_19 ));
    CascadeMux I__1875 (
            .O(N__15836),
            .I(N__15833));
    InMux I__1874 (
            .O(N__15833),
            .I(N__15830));
    LocalMux I__1873 (
            .O(N__15830),
            .I(N__15827));
    Span4Mux_v I__1872 (
            .O(N__15827),
            .I(N__15824));
    Span4Mux_v I__1871 (
            .O(N__15824),
            .I(N__15821));
    Odrv4 I__1870 (
            .O(N__15821),
            .I(\pid_alt.error_p_reg_esr_RNIH63KZ0Z_19 ));
    InMux I__1869 (
            .O(N__15818),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__1868 (
            .O(N__15815),
            .I(N__15812));
    LocalMux I__1867 (
            .O(N__15812),
            .I(N__15809));
    Odrv4 I__1866 (
            .O(N__15809),
            .I(\pid_alt.error_p_reg_esr_RNI2G981Z0Z_20 ));
    InMux I__1865 (
            .O(N__15806),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__1864 (
            .O(N__15803),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    InMux I__1863 (
            .O(N__15800),
            .I(bfn_2_18_0_));
    InMux I__1862 (
            .O(N__15797),
            .I(N__15794));
    LocalMux I__1861 (
            .O(N__15794),
            .I(N__15791));
    Odrv12 I__1860 (
            .O(N__15791),
            .I(\pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8 ));
    InMux I__1859 (
            .O(N__15788),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__1858 (
            .O(N__15785),
            .I(N__15782));
    LocalMux I__1857 (
            .O(N__15782),
            .I(N__15779));
    Odrv12 I__1856 (
            .O(N__15779),
            .I(\pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8 ));
    CascadeMux I__1855 (
            .O(N__15776),
            .I(N__15773));
    InMux I__1854 (
            .O(N__15773),
            .I(N__15770));
    LocalMux I__1853 (
            .O(N__15770),
            .I(N__15767));
    Span4Mux_v I__1852 (
            .O(N__15767),
            .I(N__15764));
    Span4Mux_v I__1851 (
            .O(N__15764),
            .I(N__15761));
    Odrv4 I__1850 (
            .O(N__15761),
            .I(\pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9 ));
    InMux I__1849 (
            .O(N__15758),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    CascadeMux I__1848 (
            .O(N__15755),
            .I(N__15751));
    InMux I__1847 (
            .O(N__15754),
            .I(N__15748));
    InMux I__1846 (
            .O(N__15751),
            .I(N__15745));
    LocalMux I__1845 (
            .O(N__15748),
            .I(N__15742));
    LocalMux I__1844 (
            .O(N__15745),
            .I(N__15739));
    Span4Mux_v I__1843 (
            .O(N__15742),
            .I(N__15736));
    Span4Mux_v I__1842 (
            .O(N__15739),
            .I(N__15733));
    Span4Mux_v I__1841 (
            .O(N__15736),
            .I(N__15730));
    Odrv4 I__1840 (
            .O(N__15733),
            .I(\pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9 ));
    Odrv4 I__1839 (
            .O(N__15730),
            .I(\pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9 ));
    CascadeMux I__1838 (
            .O(N__15725),
            .I(N__15722));
    InMux I__1837 (
            .O(N__15722),
            .I(N__15719));
    LocalMux I__1836 (
            .O(N__15719),
            .I(N__15716));
    Span4Mux_v I__1835 (
            .O(N__15716),
            .I(N__15713));
    Odrv4 I__1834 (
            .O(N__15713),
            .I(\pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10 ));
    InMux I__1833 (
            .O(N__15710),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__1832 (
            .O(N__15707),
            .I(N__15704));
    LocalMux I__1831 (
            .O(N__15704),
            .I(N__15701));
    Span4Mux_v I__1830 (
            .O(N__15701),
            .I(N__15697));
    InMux I__1829 (
            .O(N__15700),
            .I(N__15694));
    Span4Mux_v I__1828 (
            .O(N__15697),
            .I(N__15691));
    LocalMux I__1827 (
            .O(N__15694),
            .I(\pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10 ));
    Odrv4 I__1826 (
            .O(N__15691),
            .I(\pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10 ));
    CascadeMux I__1825 (
            .O(N__15686),
            .I(N__15683));
    InMux I__1824 (
            .O(N__15683),
            .I(N__15680));
    LocalMux I__1823 (
            .O(N__15680),
            .I(N__15677));
    Span4Mux_v I__1822 (
            .O(N__15677),
            .I(N__15674));
    Span4Mux_v I__1821 (
            .O(N__15674),
            .I(N__15671));
    Odrv4 I__1820 (
            .O(N__15671),
            .I(\pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11 ));
    InMux I__1819 (
            .O(N__15668),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__1818 (
            .O(N__15665),
            .I(N__15662));
    LocalMux I__1817 (
            .O(N__15662),
            .I(N__15659));
    Span4Mux_h I__1816 (
            .O(N__15659),
            .I(N__15656));
    Span4Mux_v I__1815 (
            .O(N__15656),
            .I(N__15653));
    Odrv4 I__1814 (
            .O(N__15653),
            .I(\pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12 ));
    CascadeMux I__1813 (
            .O(N__15650),
            .I(N__15647));
    InMux I__1812 (
            .O(N__15647),
            .I(N__15644));
    LocalMux I__1811 (
            .O(N__15644),
            .I(N__15641));
    Span4Mux_v I__1810 (
            .O(N__15641),
            .I(N__15638));
    Odrv4 I__1809 (
            .O(N__15638),
            .I(\pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11 ));
    InMux I__1808 (
            .O(N__15635),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__1807 (
            .O(N__15632),
            .I(N__15629));
    LocalMux I__1806 (
            .O(N__15629),
            .I(N__15626));
    Span4Mux_v I__1805 (
            .O(N__15626),
            .I(N__15623));
    Span4Mux_v I__1804 (
            .O(N__15623),
            .I(N__15620));
    Span4Mux_v I__1803 (
            .O(N__15620),
            .I(N__15617));
    Odrv4 I__1802 (
            .O(N__15617),
            .I(\pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13 ));
    CascadeMux I__1801 (
            .O(N__15614),
            .I(N__15610));
    CascadeMux I__1800 (
            .O(N__15613),
            .I(N__15607));
    InMux I__1799 (
            .O(N__15610),
            .I(N__15604));
    InMux I__1798 (
            .O(N__15607),
            .I(N__15601));
    LocalMux I__1797 (
            .O(N__15604),
            .I(N__15598));
    LocalMux I__1796 (
            .O(N__15601),
            .I(N__15595));
    Span4Mux_h I__1795 (
            .O(N__15598),
            .I(N__15592));
    Span4Mux_v I__1794 (
            .O(N__15595),
            .I(N__15587));
    Span4Mux_v I__1793 (
            .O(N__15592),
            .I(N__15587));
    Odrv4 I__1792 (
            .O(N__15587),
            .I(\pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12 ));
    InMux I__1791 (
            .O(N__15584),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__1790 (
            .O(N__15581),
            .I(N__15578));
    LocalMux I__1789 (
            .O(N__15578),
            .I(N__15575));
    Span4Mux_v I__1788 (
            .O(N__15575),
            .I(N__15572));
    Span4Mux_v I__1787 (
            .O(N__15572),
            .I(N__15569));
    Odrv4 I__1786 (
            .O(N__15569),
            .I(\pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14 ));
    CascadeMux I__1785 (
            .O(N__15566),
            .I(N__15563));
    InMux I__1784 (
            .O(N__15563),
            .I(N__15560));
    LocalMux I__1783 (
            .O(N__15560),
            .I(N__15557));
    Span4Mux_v I__1782 (
            .O(N__15557),
            .I(N__15554));
    Span4Mux_v I__1781 (
            .O(N__15554),
            .I(N__15551));
    Span4Mux_v I__1780 (
            .O(N__15551),
            .I(N__15548));
    Odrv4 I__1779 (
            .O(N__15548),
            .I(\pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13 ));
    InMux I__1778 (
            .O(N__15545),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    CascadeMux I__1777 (
            .O(N__15542),
            .I(N__15539));
    InMux I__1776 (
            .O(N__15539),
            .I(N__15536));
    LocalMux I__1775 (
            .O(N__15536),
            .I(N__15532));
    InMux I__1774 (
            .O(N__15535),
            .I(N__15529));
    Span4Mux_h I__1773 (
            .O(N__15532),
            .I(N__15524));
    LocalMux I__1772 (
            .O(N__15529),
            .I(N__15524));
    Span4Mux_v I__1771 (
            .O(N__15524),
            .I(N__15521));
    Span4Mux_v I__1770 (
            .O(N__15521),
            .I(N__15518));
    Span4Mux_v I__1769 (
            .O(N__15518),
            .I(N__15515));
    Odrv4 I__1768 (
            .O(N__15515),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__1767 (
            .O(N__15512),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__1766 (
            .O(N__15509),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__1765 (
            .O(N__15506),
            .I(N__15503));
    LocalMux I__1764 (
            .O(N__15503),
            .I(\pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1 ));
    CascadeMux I__1763 (
            .O(N__15500),
            .I(N__15497));
    InMux I__1762 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__1761 (
            .O(N__15494),
            .I(\pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2 ));
    InMux I__1760 (
            .O(N__15491),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    CascadeMux I__1759 (
            .O(N__15488),
            .I(N__15485));
    InMux I__1758 (
            .O(N__15485),
            .I(N__15481));
    InMux I__1757 (
            .O(N__15484),
            .I(N__15478));
    LocalMux I__1756 (
            .O(N__15481),
            .I(\pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2 ));
    LocalMux I__1755 (
            .O(N__15478),
            .I(\pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2 ));
    CascadeMux I__1754 (
            .O(N__15473),
            .I(N__15470));
    InMux I__1753 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__1752 (
            .O(N__15467),
            .I(N__15464));
    Odrv4 I__1751 (
            .O(N__15464),
            .I(\pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3 ));
    InMux I__1750 (
            .O(N__15461),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    InMux I__1749 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__1748 (
            .O(N__15455),
            .I(N__15452));
    Odrv4 I__1747 (
            .O(N__15452),
            .I(\pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3 ));
    CascadeMux I__1746 (
            .O(N__15449),
            .I(N__15446));
    InMux I__1745 (
            .O(N__15446),
            .I(N__15443));
    LocalMux I__1744 (
            .O(N__15443),
            .I(N__15440));
    Span4Mux_h I__1743 (
            .O(N__15440),
            .I(N__15437));
    Odrv4 I__1742 (
            .O(N__15437),
            .I(\pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4 ));
    InMux I__1741 (
            .O(N__15434),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__1740 (
            .O(N__15431),
            .I(N__15428));
    LocalMux I__1739 (
            .O(N__15428),
            .I(N__15425));
    Span4Mux_v I__1738 (
            .O(N__15425),
            .I(N__15422));
    Span4Mux_v I__1737 (
            .O(N__15422),
            .I(N__15419));
    Odrv4 I__1736 (
            .O(N__15419),
            .I(\pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5 ));
    CascadeMux I__1735 (
            .O(N__15416),
            .I(N__15413));
    InMux I__1734 (
            .O(N__15413),
            .I(N__15410));
    LocalMux I__1733 (
            .O(N__15410),
            .I(N__15406));
    CascadeMux I__1732 (
            .O(N__15409),
            .I(N__15403));
    Span4Mux_v I__1731 (
            .O(N__15406),
            .I(N__15400));
    InMux I__1730 (
            .O(N__15403),
            .I(N__15397));
    Span4Mux_v I__1729 (
            .O(N__15400),
            .I(N__15394));
    LocalMux I__1728 (
            .O(N__15397),
            .I(N__15391));
    Odrv4 I__1727 (
            .O(N__15394),
            .I(\pid_alt.error_p_reg_esr_RNI91H61Z0Z_4 ));
    Odrv4 I__1726 (
            .O(N__15391),
            .I(\pid_alt.error_p_reg_esr_RNI91H61Z0Z_4 ));
    InMux I__1725 (
            .O(N__15386),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__1724 (
            .O(N__15383),
            .I(N__15380));
    LocalMux I__1723 (
            .O(N__15380),
            .I(N__15377));
    Odrv4 I__1722 (
            .O(N__15377),
            .I(\pid_alt.error_p_reg_esr_RNI36J71Z0Z_5 ));
    CascadeMux I__1721 (
            .O(N__15374),
            .I(N__15371));
    InMux I__1720 (
            .O(N__15371),
            .I(N__15368));
    LocalMux I__1719 (
            .O(N__15368),
            .I(\pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6 ));
    InMux I__1718 (
            .O(N__15365),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__1717 (
            .O(N__15362),
            .I(N__15359));
    LocalMux I__1716 (
            .O(N__15359),
            .I(N__15355));
    InMux I__1715 (
            .O(N__15358),
            .I(N__15352));
    Span4Mux_s2_h I__1714 (
            .O(N__15355),
            .I(N__15349));
    LocalMux I__1713 (
            .O(N__15352),
            .I(N__15346));
    Span4Mux_v I__1712 (
            .O(N__15349),
            .I(N__15342));
    Span4Mux_s2_h I__1711 (
            .O(N__15346),
            .I(N__15339));
    InMux I__1710 (
            .O(N__15345),
            .I(N__15336));
    Odrv4 I__1709 (
            .O(N__15342),
            .I(drone_altitude_0));
    Odrv4 I__1708 (
            .O(N__15339),
            .I(drone_altitude_0));
    LocalMux I__1707 (
            .O(N__15336),
            .I(drone_altitude_0));
    InMux I__1706 (
            .O(N__15329),
            .I(N__15314));
    InMux I__1705 (
            .O(N__15328),
            .I(N__15314));
    InMux I__1704 (
            .O(N__15327),
            .I(N__15314));
    InMux I__1703 (
            .O(N__15326),
            .I(N__15314));
    InMux I__1702 (
            .O(N__15325),
            .I(N__15314));
    LocalMux I__1701 (
            .O(N__15314),
            .I(N__15310));
    InMux I__1700 (
            .O(N__15313),
            .I(N__15307));
    Span4Mux_s3_h I__1699 (
            .O(N__15310),
            .I(N__15301));
    LocalMux I__1698 (
            .O(N__15307),
            .I(N__15298));
    InMux I__1697 (
            .O(N__15306),
            .I(N__15293));
    InMux I__1696 (
            .O(N__15305),
            .I(N__15293));
    InMux I__1695 (
            .O(N__15304),
            .I(N__15290));
    Odrv4 I__1694 (
            .O(N__15301),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ));
    Odrv12 I__1693 (
            .O(N__15298),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ));
    LocalMux I__1692 (
            .O(N__15293),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ));
    LocalMux I__1691 (
            .O(N__15290),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ));
    InMux I__1690 (
            .O(N__15281),
            .I(N__15278));
    LocalMux I__1689 (
            .O(N__15278),
            .I(\pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14 ));
    CascadeMux I__1688 (
            .O(N__15275),
            .I(\pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_ ));
    CascadeMux I__1687 (
            .O(N__15272),
            .I(\pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_ ));
    InMux I__1686 (
            .O(N__15269),
            .I(N__15265));
    InMux I__1685 (
            .O(N__15268),
            .I(N__15262));
    LocalMux I__1684 (
            .O(N__15265),
            .I(N__15255));
    LocalMux I__1683 (
            .O(N__15262),
            .I(N__15255));
    InMux I__1682 (
            .O(N__15261),
            .I(N__15250));
    InMux I__1681 (
            .O(N__15260),
            .I(N__15250));
    Odrv4 I__1680 (
            .O(N__15255),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__1679 (
            .O(N__15250),
            .I(\pid_alt.N_9_0 ));
    InMux I__1678 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__1677 (
            .O(N__15242),
            .I(N__15239));
    Odrv4 I__1676 (
            .O(N__15239),
            .I(\pid_alt.m21_e_9 ));
    CascadeMux I__1675 (
            .O(N__15236),
            .I(\pid_alt.N_9_0_cascade_ ));
    InMux I__1674 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__1673 (
            .O(N__15230),
            .I(N__15227));
    Odrv4 I__1672 (
            .O(N__15227),
            .I(\pid_alt.m21_e_10 ));
    CascadeMux I__1671 (
            .O(N__15224),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_ ));
    SRMux I__1670 (
            .O(N__15221),
            .I(N__15218));
    LocalMux I__1669 (
            .O(N__15218),
            .I(N__15213));
    SRMux I__1668 (
            .O(N__15217),
            .I(N__15209));
    SRMux I__1667 (
            .O(N__15216),
            .I(N__15205));
    Span4Mux_v I__1666 (
            .O(N__15213),
            .I(N__15202));
    SRMux I__1665 (
            .O(N__15212),
            .I(N__15199));
    LocalMux I__1664 (
            .O(N__15209),
            .I(N__15196));
    SRMux I__1663 (
            .O(N__15208),
            .I(N__15193));
    LocalMux I__1662 (
            .O(N__15205),
            .I(N__15190));
    Span4Mux_v I__1661 (
            .O(N__15202),
            .I(N__15185));
    LocalMux I__1660 (
            .O(N__15199),
            .I(N__15185));
    Span4Mux_v I__1659 (
            .O(N__15196),
            .I(N__15180));
    LocalMux I__1658 (
            .O(N__15193),
            .I(N__15180));
    Odrv4 I__1657 (
            .O(N__15190),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__1656 (
            .O(N__15185),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__1655 (
            .O(N__15180),
            .I(\pid_alt.un1_reset_1_0_i ));
    CascadeMux I__1654 (
            .O(N__15173),
            .I(\pid_alt.un1_reset_1_0_i_cascade_ ));
    CEMux I__1653 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__1652 (
            .O(N__15167),
            .I(N__15163));
    CEMux I__1651 (
            .O(N__15166),
            .I(N__15160));
    Span4Mux_v I__1650 (
            .O(N__15163),
            .I(N__15154));
    LocalMux I__1649 (
            .O(N__15160),
            .I(N__15154));
    CEMux I__1648 (
            .O(N__15159),
            .I(N__15151));
    Span4Mux_h I__1647 (
            .O(N__15154),
            .I(N__15148));
    LocalMux I__1646 (
            .O(N__15151),
            .I(N__15143));
    Span4Mux_s1_h I__1645 (
            .O(N__15148),
            .I(N__15143));
    Odrv4 I__1644 (
            .O(N__15143),
            .I(\pid_alt.N_60_i_0 ));
    InMux I__1643 (
            .O(N__15140),
            .I(\scaler_2.un3_source_data_0_cry_1 ));
    InMux I__1642 (
            .O(N__15137),
            .I(\scaler_2.un3_source_data_0_cry_2 ));
    InMux I__1641 (
            .O(N__15134),
            .I(\scaler_2.un3_source_data_0_cry_3 ));
    InMux I__1640 (
            .O(N__15131),
            .I(\scaler_2.un3_source_data_0_cry_4 ));
    InMux I__1639 (
            .O(N__15128),
            .I(\scaler_2.un3_source_data_0_cry_5 ));
    InMux I__1638 (
            .O(N__15125),
            .I(\scaler_2.un3_source_data_0_cry_6 ));
    InMux I__1637 (
            .O(N__15122),
            .I(bfn_2_15_0_));
    InMux I__1636 (
            .O(N__15119),
            .I(\scaler_2.un3_source_data_0_cry_8 ));
    CascadeMux I__1635 (
            .O(N__15116),
            .I(N__15113));
    InMux I__1634 (
            .O(N__15113),
            .I(N__15110));
    LocalMux I__1633 (
            .O(N__15110),
            .I(N__15106));
    InMux I__1632 (
            .O(N__15109),
            .I(N__15103));
    Span4Mux_s3_h I__1631 (
            .O(N__15106),
            .I(N__15100));
    LocalMux I__1630 (
            .O(N__15103),
            .I(\pid_alt.drone_altitude_i_0 ));
    Odrv4 I__1629 (
            .O(N__15100),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__1628 (
            .O(N__15095),
            .I(N__15089));
    InMux I__1627 (
            .O(N__15094),
            .I(N__15089));
    LocalMux I__1626 (
            .O(N__15089),
            .I(N__15086));
    Span4Mux_s2_h I__1625 (
            .O(N__15086),
            .I(N__15083));
    Odrv4 I__1624 (
            .O(N__15083),
            .I(\pid_alt.m35_e_2 ));
    CascadeMux I__1623 (
            .O(N__15080),
            .I(\pid_alt.m35_e_2_cascade_ ));
    InMux I__1622 (
            .O(N__15077),
            .I(N__15074));
    LocalMux I__1621 (
            .O(N__15074),
            .I(N__15071));
    Span4Mux_v I__1620 (
            .O(N__15071),
            .I(N__15068));
    Odrv4 I__1619 (
            .O(N__15068),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5 ));
    CascadeMux I__1618 (
            .O(N__15065),
            .I(N__15061));
    CascadeMux I__1617 (
            .O(N__15064),
            .I(N__15058));
    InMux I__1616 (
            .O(N__15061),
            .I(N__15053));
    InMux I__1615 (
            .O(N__15058),
            .I(N__15053));
    LocalMux I__1614 (
            .O(N__15053),
            .I(N__15050));
    Span4Mux_v I__1613 (
            .O(N__15050),
            .I(N__15046));
    InMux I__1612 (
            .O(N__15049),
            .I(N__15043));
    Odrv4 I__1611 (
            .O(N__15046),
            .I(\pid_alt.m35_e_3 ));
    LocalMux I__1610 (
            .O(N__15043),
            .I(\pid_alt.m35_e_3 ));
    CascadeMux I__1609 (
            .O(N__15038),
            .I(\pid_alt.m21_e_2_cascade_ ));
    CascadeMux I__1608 (
            .O(N__15035),
            .I(\pid_alt.m21_e_0_cascade_ ));
    InMux I__1607 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__1606 (
            .O(N__15029),
            .I(\pid_alt.m21_e_8 ));
    InMux I__1605 (
            .O(N__15026),
            .I(\scaler_2.un3_source_data_0_cry_0 ));
    InMux I__1604 (
            .O(N__15023),
            .I(N__15020));
    LocalMux I__1603 (
            .O(N__15020),
            .I(N__15016));
    InMux I__1602 (
            .O(N__15019),
            .I(N__15013));
    Span4Mux_v I__1601 (
            .O(N__15016),
            .I(N__15010));
    LocalMux I__1600 (
            .O(N__15013),
            .I(N__15007));
    Span4Mux_v I__1599 (
            .O(N__15010),
            .I(N__15002));
    Span4Mux_s1_h I__1598 (
            .O(N__15007),
            .I(N__15002));
    Odrv4 I__1597 (
            .O(N__15002),
            .I(\pid_alt.error_8 ));
    InMux I__1596 (
            .O(N__14999),
            .I(bfn_2_12_0_));
    InMux I__1595 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__1594 (
            .O(N__14993),
            .I(N__14989));
    InMux I__1593 (
            .O(N__14992),
            .I(N__14986));
    Span4Mux_v I__1592 (
            .O(N__14989),
            .I(N__14983));
    LocalMux I__1591 (
            .O(N__14986),
            .I(N__14980));
    Span4Mux_v I__1590 (
            .O(N__14983),
            .I(N__14975));
    Span4Mux_s1_h I__1589 (
            .O(N__14980),
            .I(N__14975));
    Odrv4 I__1588 (
            .O(N__14975),
            .I(\pid_alt.error_9 ));
    InMux I__1587 (
            .O(N__14972),
            .I(\pid_alt.error_cry_8 ));
    InMux I__1586 (
            .O(N__14969),
            .I(N__14966));
    LocalMux I__1585 (
            .O(N__14966),
            .I(N__14962));
    InMux I__1584 (
            .O(N__14965),
            .I(N__14959));
    Span4Mux_v I__1583 (
            .O(N__14962),
            .I(N__14956));
    LocalMux I__1582 (
            .O(N__14959),
            .I(N__14953));
    Span4Mux_v I__1581 (
            .O(N__14956),
            .I(N__14948));
    Span4Mux_s1_h I__1580 (
            .O(N__14953),
            .I(N__14948));
    Odrv4 I__1579 (
            .O(N__14948),
            .I(\pid_alt.error_10 ));
    InMux I__1578 (
            .O(N__14945),
            .I(\pid_alt.error_cry_9 ));
    InMux I__1577 (
            .O(N__14942),
            .I(N__14939));
    LocalMux I__1576 (
            .O(N__14939),
            .I(N__14936));
    Span4Mux_v I__1575 (
            .O(N__14936),
            .I(N__14932));
    InMux I__1574 (
            .O(N__14935),
            .I(N__14929));
    Span4Mux_v I__1573 (
            .O(N__14932),
            .I(N__14924));
    LocalMux I__1572 (
            .O(N__14929),
            .I(N__14924));
    Span4Mux_s1_h I__1571 (
            .O(N__14924),
            .I(N__14921));
    Odrv4 I__1570 (
            .O(N__14921),
            .I(\pid_alt.error_11 ));
    InMux I__1569 (
            .O(N__14918),
            .I(\pid_alt.error_cry_10 ));
    InMux I__1568 (
            .O(N__14915),
            .I(N__14912));
    LocalMux I__1567 (
            .O(N__14912),
            .I(N__14909));
    Span4Mux_v I__1566 (
            .O(N__14909),
            .I(N__14905));
    InMux I__1565 (
            .O(N__14908),
            .I(N__14902));
    Span4Mux_v I__1564 (
            .O(N__14905),
            .I(N__14897));
    LocalMux I__1563 (
            .O(N__14902),
            .I(N__14897));
    Odrv4 I__1562 (
            .O(N__14897),
            .I(\pid_alt.error_12 ));
    InMux I__1561 (
            .O(N__14894),
            .I(\pid_alt.error_cry_11 ));
    InMux I__1560 (
            .O(N__14891),
            .I(N__14888));
    LocalMux I__1559 (
            .O(N__14888),
            .I(N__14885));
    Span4Mux_v I__1558 (
            .O(N__14885),
            .I(N__14881));
    InMux I__1557 (
            .O(N__14884),
            .I(N__14878));
    Span4Mux_v I__1556 (
            .O(N__14881),
            .I(N__14873));
    LocalMux I__1555 (
            .O(N__14878),
            .I(N__14873));
    Odrv4 I__1554 (
            .O(N__14873),
            .I(\pid_alt.error_13 ));
    InMux I__1553 (
            .O(N__14870),
            .I(\pid_alt.error_cry_12 ));
    InMux I__1552 (
            .O(N__14867),
            .I(N__14864));
    LocalMux I__1551 (
            .O(N__14864),
            .I(N__14861));
    Span4Mux_v I__1550 (
            .O(N__14861),
            .I(N__14857));
    InMux I__1549 (
            .O(N__14860),
            .I(N__14854));
    Span4Mux_v I__1548 (
            .O(N__14857),
            .I(N__14849));
    LocalMux I__1547 (
            .O(N__14854),
            .I(N__14849));
    Odrv4 I__1546 (
            .O(N__14849),
            .I(\pid_alt.error_14 ));
    InMux I__1545 (
            .O(N__14846),
            .I(\pid_alt.error_cry_13 ));
    InMux I__1544 (
            .O(N__14843),
            .I(\pid_alt.error_cry_14 ));
    InMux I__1543 (
            .O(N__14840),
            .I(N__14837));
    LocalMux I__1542 (
            .O(N__14837),
            .I(N__14834));
    Span4Mux_v I__1541 (
            .O(N__14834),
            .I(N__14830));
    InMux I__1540 (
            .O(N__14833),
            .I(N__14827));
    Span4Mux_v I__1539 (
            .O(N__14830),
            .I(N__14822));
    LocalMux I__1538 (
            .O(N__14827),
            .I(N__14822));
    Odrv4 I__1537 (
            .O(N__14822),
            .I(\pid_alt.error_15 ));
    InMux I__1536 (
            .O(N__14819),
            .I(N__14813));
    InMux I__1535 (
            .O(N__14818),
            .I(N__14813));
    LocalMux I__1534 (
            .O(N__14813),
            .I(N__14810));
    Span4Mux_v I__1533 (
            .O(N__14810),
            .I(N__14807));
    Odrv4 I__1532 (
            .O(N__14807),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    InMux I__1531 (
            .O(N__14804),
            .I(N__14800));
    InMux I__1530 (
            .O(N__14803),
            .I(N__14797));
    LocalMux I__1529 (
            .O(N__14800),
            .I(N__14794));
    LocalMux I__1528 (
            .O(N__14797),
            .I(N__14791));
    Span4Mux_s2_h I__1527 (
            .O(N__14794),
            .I(N__14788));
    Span4Mux_s3_h I__1526 (
            .O(N__14791),
            .I(N__14785));
    Odrv4 I__1525 (
            .O(N__14788),
            .I(\pid_alt.error_1 ));
    Odrv4 I__1524 (
            .O(N__14785),
            .I(\pid_alt.error_1 ));
    InMux I__1523 (
            .O(N__14780),
            .I(\pid_alt.error_cry_0 ));
    InMux I__1522 (
            .O(N__14777),
            .I(N__14773));
    InMux I__1521 (
            .O(N__14776),
            .I(N__14770));
    LocalMux I__1520 (
            .O(N__14773),
            .I(N__14767));
    LocalMux I__1519 (
            .O(N__14770),
            .I(N__14764));
    Span4Mux_s3_h I__1518 (
            .O(N__14767),
            .I(N__14761));
    Span4Mux_s2_h I__1517 (
            .O(N__14764),
            .I(N__14758));
    Odrv4 I__1516 (
            .O(N__14761),
            .I(\pid_alt.error_2 ));
    Odrv4 I__1515 (
            .O(N__14758),
            .I(\pid_alt.error_2 ));
    InMux I__1514 (
            .O(N__14753),
            .I(\pid_alt.error_cry_1 ));
    InMux I__1513 (
            .O(N__14750),
            .I(N__14746));
    InMux I__1512 (
            .O(N__14749),
            .I(N__14743));
    LocalMux I__1511 (
            .O(N__14746),
            .I(N__14740));
    LocalMux I__1510 (
            .O(N__14743),
            .I(N__14737));
    Span4Mux_s2_h I__1509 (
            .O(N__14740),
            .I(N__14734));
    Span4Mux_s2_h I__1508 (
            .O(N__14737),
            .I(N__14731));
    Odrv4 I__1507 (
            .O(N__14734),
            .I(\pid_alt.error_3 ));
    Odrv4 I__1506 (
            .O(N__14731),
            .I(\pid_alt.error_3 ));
    InMux I__1505 (
            .O(N__14726),
            .I(\pid_alt.error_cry_2 ));
    InMux I__1504 (
            .O(N__14723),
            .I(N__14719));
    InMux I__1503 (
            .O(N__14722),
            .I(N__14716));
    LocalMux I__1502 (
            .O(N__14719),
            .I(N__14713));
    LocalMux I__1501 (
            .O(N__14716),
            .I(N__14710));
    Span4Mux_v I__1500 (
            .O(N__14713),
            .I(N__14707));
    Span4Mux_s3_h I__1499 (
            .O(N__14710),
            .I(N__14704));
    Span4Mux_s0_h I__1498 (
            .O(N__14707),
            .I(N__14701));
    Odrv4 I__1497 (
            .O(N__14704),
            .I(\pid_alt.error_4 ));
    Odrv4 I__1496 (
            .O(N__14701),
            .I(\pid_alt.error_4 ));
    InMux I__1495 (
            .O(N__14696),
            .I(\pid_alt.error_cry_3 ));
    InMux I__1494 (
            .O(N__14693),
            .I(N__14689));
    InMux I__1493 (
            .O(N__14692),
            .I(N__14686));
    LocalMux I__1492 (
            .O(N__14689),
            .I(N__14683));
    LocalMux I__1491 (
            .O(N__14686),
            .I(N__14680));
    Span4Mux_s2_h I__1490 (
            .O(N__14683),
            .I(N__14677));
    Span4Mux_v I__1489 (
            .O(N__14680),
            .I(N__14674));
    Odrv4 I__1488 (
            .O(N__14677),
            .I(\pid_alt.error_5 ));
    Odrv4 I__1487 (
            .O(N__14674),
            .I(\pid_alt.error_5 ));
    InMux I__1486 (
            .O(N__14669),
            .I(\pid_alt.error_cry_4 ));
    InMux I__1485 (
            .O(N__14666),
            .I(N__14663));
    LocalMux I__1484 (
            .O(N__14663),
            .I(N__14659));
    InMux I__1483 (
            .O(N__14662),
            .I(N__14656));
    Span4Mux_s1_h I__1482 (
            .O(N__14659),
            .I(N__14653));
    LocalMux I__1481 (
            .O(N__14656),
            .I(N__14650));
    Span4Mux_v I__1480 (
            .O(N__14653),
            .I(N__14647));
    Span4Mux_s2_h I__1479 (
            .O(N__14650),
            .I(N__14644));
    Odrv4 I__1478 (
            .O(N__14647),
            .I(\pid_alt.error_6 ));
    Odrv4 I__1477 (
            .O(N__14644),
            .I(\pid_alt.error_6 ));
    InMux I__1476 (
            .O(N__14639),
            .I(\pid_alt.error_cry_5 ));
    InMux I__1475 (
            .O(N__14636),
            .I(N__14633));
    LocalMux I__1474 (
            .O(N__14633),
            .I(N__14629));
    InMux I__1473 (
            .O(N__14632),
            .I(N__14626));
    Span4Mux_s1_h I__1472 (
            .O(N__14629),
            .I(N__14623));
    LocalMux I__1471 (
            .O(N__14626),
            .I(N__14620));
    Span4Mux_v I__1470 (
            .O(N__14623),
            .I(N__14617));
    Span4Mux_s2_h I__1469 (
            .O(N__14620),
            .I(N__14614));
    Odrv4 I__1468 (
            .O(N__14617),
            .I(\pid_alt.error_7 ));
    Odrv4 I__1467 (
            .O(N__14614),
            .I(\pid_alt.error_7 ));
    InMux I__1466 (
            .O(N__14609),
            .I(\pid_alt.error_cry_6 ));
    InMux I__1465 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__1464 (
            .O(N__14603),
            .I(N__14600));
    Span4Mux_v I__1463 (
            .O(N__14600),
            .I(N__14597));
    Span4Mux_s1_h I__1462 (
            .O(N__14597),
            .I(N__14594));
    Odrv4 I__1461 (
            .O(N__14594),
            .I(alt_ki_2));
    InMux I__1460 (
            .O(N__14591),
            .I(N__14588));
    LocalMux I__1459 (
            .O(N__14588),
            .I(N__14585));
    Span4Mux_s3_h I__1458 (
            .O(N__14585),
            .I(N__14582));
    Odrv4 I__1457 (
            .O(N__14582),
            .I(alt_ki_3));
    InMux I__1456 (
            .O(N__14579),
            .I(N__14576));
    LocalMux I__1455 (
            .O(N__14576),
            .I(N__14573));
    Span4Mux_s3_h I__1454 (
            .O(N__14573),
            .I(N__14570));
    Odrv4 I__1453 (
            .O(N__14570),
            .I(alt_ki_5));
    InMux I__1452 (
            .O(N__14567),
            .I(N__14564));
    LocalMux I__1451 (
            .O(N__14564),
            .I(N__14561));
    Span4Mux_v I__1450 (
            .O(N__14561),
            .I(N__14558));
    Odrv4 I__1449 (
            .O(N__14558),
            .I(alt_ki_6));
    InMux I__1448 (
            .O(N__14555),
            .I(N__14552));
    LocalMux I__1447 (
            .O(N__14552),
            .I(N__14549));
    Span4Mux_h I__1446 (
            .O(N__14549),
            .I(N__14546));
    Odrv4 I__1445 (
            .O(N__14546),
            .I(\pid_alt.O_12 ));
    InMux I__1444 (
            .O(N__14543),
            .I(N__14537));
    InMux I__1443 (
            .O(N__14542),
            .I(N__14537));
    LocalMux I__1442 (
            .O(N__14537),
            .I(N__14534));
    Span4Mux_v I__1441 (
            .O(N__14534),
            .I(N__14531));
    Odrv4 I__1440 (
            .O(N__14531),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    CascadeMux I__1439 (
            .O(N__14528),
            .I(\pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_ ));
    InMux I__1438 (
            .O(N__14525),
            .I(N__14522));
    LocalMux I__1437 (
            .O(N__14522),
            .I(N__14519));
    Span4Mux_h I__1436 (
            .O(N__14519),
            .I(N__14516));
    Odrv4 I__1435 (
            .O(N__14516),
            .I(\pid_alt.O_13 ));
    InMux I__1434 (
            .O(N__14513),
            .I(N__14510));
    LocalMux I__1433 (
            .O(N__14510),
            .I(N__14507));
    Span4Mux_v I__1432 (
            .O(N__14507),
            .I(N__14504));
    Odrv4 I__1431 (
            .O(N__14504),
            .I(\pid_alt.O_0_8 ));
    InMux I__1430 (
            .O(N__14501),
            .I(N__14495));
    InMux I__1429 (
            .O(N__14500),
            .I(N__14495));
    LocalMux I__1428 (
            .O(N__14495),
            .I(N__14492));
    Sp12to4 I__1427 (
            .O(N__14492),
            .I(N__14489));
    Span12Mux_v I__1426 (
            .O(N__14489),
            .I(N__14486));
    Odrv12 I__1425 (
            .O(N__14486),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    InMux I__1424 (
            .O(N__14483),
            .I(N__14480));
    LocalMux I__1423 (
            .O(N__14480),
            .I(N__14477));
    Span4Mux_s3_h I__1422 (
            .O(N__14477),
            .I(N__14474));
    Odrv4 I__1421 (
            .O(N__14474),
            .I(alt_kp_2));
    InMux I__1420 (
            .O(N__14471),
            .I(N__14468));
    LocalMux I__1419 (
            .O(N__14468),
            .I(N__14465));
    Span4Mux_s2_h I__1418 (
            .O(N__14465),
            .I(N__14462));
    Odrv4 I__1417 (
            .O(N__14462),
            .I(alt_ki_4));
    InMux I__1416 (
            .O(N__14459),
            .I(N__14456));
    LocalMux I__1415 (
            .O(N__14456),
            .I(N__14453));
    Span12Mux_s2_h I__1414 (
            .O(N__14453),
            .I(N__14450));
    Odrv12 I__1413 (
            .O(N__14450),
            .I(alt_ki_1));
    CascadeMux I__1412 (
            .O(N__14447),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ));
    CascadeMux I__1411 (
            .O(N__14444),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ));
    InMux I__1410 (
            .O(N__14441),
            .I(N__14438));
    LocalMux I__1409 (
            .O(N__14438),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9 ));
    InMux I__1408 (
            .O(N__14435),
            .I(N__14430));
    InMux I__1407 (
            .O(N__14434),
            .I(N__14425));
    InMux I__1406 (
            .O(N__14433),
            .I(N__14425));
    LocalMux I__1405 (
            .O(N__14430),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__1404 (
            .O(N__14425),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__1403 (
            .O(N__14420),
            .I(N__14417));
    LocalMux I__1402 (
            .O(N__14417),
            .I(N__14414));
    Odrv12 I__1401 (
            .O(N__14414),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__1400 (
            .O(N__14411),
            .I(N__14408));
    LocalMux I__1399 (
            .O(N__14408),
            .I(N__14403));
    InMux I__1398 (
            .O(N__14407),
            .I(N__14400));
    InMux I__1397 (
            .O(N__14406),
            .I(N__14397));
    Span4Mux_v I__1396 (
            .O(N__14403),
            .I(N__14392));
    LocalMux I__1395 (
            .O(N__14400),
            .I(N__14392));
    LocalMux I__1394 (
            .O(N__14397),
            .I(throttle_command_9));
    Odrv4 I__1393 (
            .O(N__14392),
            .I(throttle_command_9));
    CascadeMux I__1392 (
            .O(N__14387),
            .I(N__14384));
    InMux I__1391 (
            .O(N__14384),
            .I(N__14379));
    InMux I__1390 (
            .O(N__14383),
            .I(N__14374));
    InMux I__1389 (
            .O(N__14382),
            .I(N__14374));
    LocalMux I__1388 (
            .O(N__14379),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    LocalMux I__1387 (
            .O(N__14374),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__1386 (
            .O(N__14369),
            .I(N__14364));
    InMux I__1385 (
            .O(N__14368),
            .I(N__14359));
    InMux I__1384 (
            .O(N__14367),
            .I(N__14359));
    LocalMux I__1383 (
            .O(N__14364),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    LocalMux I__1382 (
            .O(N__14359),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    CascadeMux I__1381 (
            .O(N__14354),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ));
    InMux I__1380 (
            .O(N__14351),
            .I(N__14348));
    LocalMux I__1379 (
            .O(N__14348),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10 ));
    InMux I__1378 (
            .O(N__14345),
            .I(N__14341));
    InMux I__1377 (
            .O(N__14344),
            .I(N__14338));
    LocalMux I__1376 (
            .O(N__14341),
            .I(N__14335));
    LocalMux I__1375 (
            .O(N__14338),
            .I(N__14332));
    Odrv4 I__1374 (
            .O(N__14335),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    Odrv4 I__1373 (
            .O(N__14332),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__1372 (
            .O(N__14327),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ));
    InMux I__1371 (
            .O(N__14324),
            .I(N__14321));
    LocalMux I__1370 (
            .O(N__14321),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    CascadeMux I__1369 (
            .O(N__14318),
            .I(\ppm_encoder_1.un1_init_pulses_10_0_cascade_ ));
    CascadeMux I__1368 (
            .O(N__14315),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ));
    InMux I__1367 (
            .O(N__14312),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    CascadeMux I__1366 (
            .O(N__14309),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ));
    CascadeMux I__1365 (
            .O(N__14306),
            .I(N__14301));
    InMux I__1364 (
            .O(N__14305),
            .I(N__14298));
    InMux I__1363 (
            .O(N__14304),
            .I(N__14295));
    InMux I__1362 (
            .O(N__14301),
            .I(N__14292));
    LocalMux I__1361 (
            .O(N__14298),
            .I(N__14287));
    LocalMux I__1360 (
            .O(N__14295),
            .I(N__14287));
    LocalMux I__1359 (
            .O(N__14292),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__1358 (
            .O(N__14287),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__1357 (
            .O(N__14282),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    InMux I__1356 (
            .O(N__14279),
            .I(N__14276));
    LocalMux I__1355 (
            .O(N__14276),
            .I(N__14273));
    Span4Mux_v I__1354 (
            .O(N__14273),
            .I(N__14270));
    Odrv4 I__1353 (
            .O(N__14270),
            .I(scaler_2_data_5));
    InMux I__1352 (
            .O(N__14267),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__1351 (
            .O(N__14264),
            .I(N__14259));
    InMux I__1350 (
            .O(N__14263),
            .I(N__14256));
    InMux I__1349 (
            .O(N__14262),
            .I(N__14253));
    LocalMux I__1348 (
            .O(N__14259),
            .I(N__14250));
    LocalMux I__1347 (
            .O(N__14256),
            .I(throttle_command_6));
    LocalMux I__1346 (
            .O(N__14253),
            .I(throttle_command_6));
    Odrv4 I__1345 (
            .O(N__14250),
            .I(throttle_command_6));
    InMux I__1344 (
            .O(N__14243),
            .I(N__14240));
    LocalMux I__1343 (
            .O(N__14240),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    InMux I__1342 (
            .O(N__14237),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__1341 (
            .O(N__14234),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__1340 (
            .O(N__14231),
            .I(bfn_1_23_0_));
    InMux I__1339 (
            .O(N__14228),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__1338 (
            .O(N__14225),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__1337 (
            .O(N__14222),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__1336 (
            .O(N__14219),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__1335 (
            .O(N__14216),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__1334 (
            .O(N__14213),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__1333 (
            .O(N__14210),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__1332 (
            .O(N__14207),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__1331 (
            .O(N__14204),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__1330 (
            .O(N__14201),
            .I(N__14198));
    LocalMux I__1329 (
            .O(N__14198),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__1328 (
            .O(N__14195),
            .I(N__14192));
    LocalMux I__1327 (
            .O(N__14192),
            .I(N__14188));
    InMux I__1326 (
            .O(N__14191),
            .I(N__14185));
    Odrv12 I__1325 (
            .O(N__14188),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    LocalMux I__1324 (
            .O(N__14185),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    CascadeMux I__1323 (
            .O(N__14180),
            .I(\pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_ ));
    CascadeMux I__1322 (
            .O(N__14177),
            .I(N__14174));
    InMux I__1321 (
            .O(N__14174),
            .I(N__14169));
    InMux I__1320 (
            .O(N__14173),
            .I(N__14166));
    InMux I__1319 (
            .O(N__14172),
            .I(N__14163));
    LocalMux I__1318 (
            .O(N__14169),
            .I(N__14158));
    LocalMux I__1317 (
            .O(N__14166),
            .I(N__14158));
    LocalMux I__1316 (
            .O(N__14163),
            .I(N__14155));
    Span12Mux_v I__1315 (
            .O(N__14158),
            .I(N__14152));
    Span4Mux_v I__1314 (
            .O(N__14155),
            .I(N__14149));
    Odrv12 I__1313 (
            .O(N__14152),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    Odrv4 I__1312 (
            .O(N__14149),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    InMux I__1311 (
            .O(N__14144),
            .I(N__14141));
    LocalMux I__1310 (
            .O(N__14141),
            .I(N__14138));
    Span12Mux_v I__1309 (
            .O(N__14138),
            .I(N__14135));
    Odrv12 I__1308 (
            .O(N__14135),
            .I(alt_ki_0));
    CascadeMux I__1307 (
            .O(N__14132),
            .I(\pid_alt.N_37_cascade_ ));
    InMux I__1306 (
            .O(N__14129),
            .I(N__14122));
    InMux I__1305 (
            .O(N__14128),
            .I(N__14117));
    InMux I__1304 (
            .O(N__14127),
            .I(N__14117));
    InMux I__1303 (
            .O(N__14126),
            .I(N__14114));
    InMux I__1302 (
            .O(N__14125),
            .I(N__14111));
    LocalMux I__1301 (
            .O(N__14122),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__1300 (
            .O(N__14117),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__1299 (
            .O(N__14114),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__1298 (
            .O(N__14111),
            .I(\pid_alt.N_62_mux ));
    InMux I__1297 (
            .O(N__14102),
            .I(N__14097));
    InMux I__1296 (
            .O(N__14101),
            .I(N__14092));
    InMux I__1295 (
            .O(N__14100),
            .I(N__14092));
    LocalMux I__1294 (
            .O(N__14097),
            .I(\pid_alt.N_37 ));
    LocalMux I__1293 (
            .O(N__14092),
            .I(\pid_alt.N_37 ));
    InMux I__1292 (
            .O(N__14087),
            .I(N__14081));
    InMux I__1291 (
            .O(N__14086),
            .I(N__14081));
    LocalMux I__1290 (
            .O(N__14081),
            .I(N__14078));
    Odrv12 I__1289 (
            .O(N__14078),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    CascadeMux I__1288 (
            .O(N__14075),
            .I(\pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_ ));
    InMux I__1287 (
            .O(N__14072),
            .I(N__14066));
    InMux I__1286 (
            .O(N__14071),
            .I(N__14066));
    LocalMux I__1285 (
            .O(N__14066),
            .I(N__14063));
    Span4Mux_v I__1284 (
            .O(N__14063),
            .I(N__14060));
    Sp12to4 I__1283 (
            .O(N__14060),
            .I(N__14057));
    Odrv12 I__1282 (
            .O(N__14057),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    CascadeMux I__1281 (
            .O(N__14054),
            .I(N__14051));
    InMux I__1280 (
            .O(N__14051),
            .I(N__14048));
    LocalMux I__1279 (
            .O(N__14048),
            .I(N__14045));
    Sp12to4 I__1278 (
            .O(N__14045),
            .I(N__14040));
    InMux I__1277 (
            .O(N__14044),
            .I(N__14035));
    InMux I__1276 (
            .O(N__14043),
            .I(N__14035));
    Span12Mux_v I__1275 (
            .O(N__14040),
            .I(N__14030));
    LocalMux I__1274 (
            .O(N__14035),
            .I(N__14030));
    Odrv12 I__1273 (
            .O(N__14030),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    CascadeMux I__1272 (
            .O(N__14027),
            .I(\pid_alt.N_62_mux_cascade_ ));
    CascadeMux I__1271 (
            .O(N__14024),
            .I(\pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_ ));
    InMux I__1270 (
            .O(N__14021),
            .I(N__14015));
    InMux I__1269 (
            .O(N__14020),
            .I(N__14015));
    LocalMux I__1268 (
            .O(N__14015),
            .I(N__14012));
    Span4Mux_v I__1267 (
            .O(N__14012),
            .I(N__14009));
    Span4Mux_v I__1266 (
            .O(N__14009),
            .I(N__14006));
    Odrv4 I__1265 (
            .O(N__14006),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__1264 (
            .O(N__14003),
            .I(N__14000));
    LocalMux I__1263 (
            .O(N__14000),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5 ));
    InMux I__1262 (
            .O(N__13997),
            .I(N__13994));
    LocalMux I__1261 (
            .O(N__13994),
            .I(N__13991));
    Odrv4 I__1260 (
            .O(N__13991),
            .I(\pid_alt.O_9 ));
    InMux I__1259 (
            .O(N__13988),
            .I(N__13985));
    LocalMux I__1258 (
            .O(N__13985),
            .I(N__13982));
    Odrv4 I__1257 (
            .O(N__13982),
            .I(\pid_alt.O_8 ));
    CascadeMux I__1256 (
            .O(N__13979),
            .I(\pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_ ));
    InMux I__1255 (
            .O(N__13976),
            .I(N__13973));
    LocalMux I__1254 (
            .O(N__13973),
            .I(\pid_alt.O_16 ));
    InMux I__1253 (
            .O(N__13970),
            .I(N__13964));
    InMux I__1252 (
            .O(N__13969),
            .I(N__13964));
    LocalMux I__1251 (
            .O(N__13964),
            .I(N__13961));
    Span4Mux_v I__1250 (
            .O(N__13961),
            .I(N__13958));
    Odrv4 I__1249 (
            .O(N__13958),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__1248 (
            .O(N__13955),
            .I(N__13952));
    LocalMux I__1247 (
            .O(N__13952),
            .I(\pid_alt.O_14 ));
    InMux I__1246 (
            .O(N__13949),
            .I(N__13943));
    InMux I__1245 (
            .O(N__13948),
            .I(N__13943));
    LocalMux I__1244 (
            .O(N__13943),
            .I(N__13940));
    Odrv12 I__1243 (
            .O(N__13940),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__1242 (
            .O(N__13937),
            .I(N__13934));
    LocalMux I__1241 (
            .O(N__13934),
            .I(N__13931));
    Span4Mux_h I__1240 (
            .O(N__13931),
            .I(N__13928));
    Odrv4 I__1239 (
            .O(N__13928),
            .I(\pid_alt.O_5 ));
    InMux I__1238 (
            .O(N__13925),
            .I(N__13922));
    LocalMux I__1237 (
            .O(N__13922),
            .I(N__13919));
    Span4Mux_h I__1236 (
            .O(N__13919),
            .I(N__13916));
    Odrv4 I__1235 (
            .O(N__13916),
            .I(\pid_alt.O_7 ));
    InMux I__1234 (
            .O(N__13913),
            .I(N__13910));
    LocalMux I__1233 (
            .O(N__13910),
            .I(N__13907));
    Odrv4 I__1232 (
            .O(N__13907),
            .I(\pid_alt.O_19 ));
    InMux I__1231 (
            .O(N__13904),
            .I(N__13901));
    LocalMux I__1230 (
            .O(N__13901),
            .I(N__13898));
    Odrv4 I__1229 (
            .O(N__13898),
            .I(\pid_alt.O_20 ));
    InMux I__1228 (
            .O(N__13895),
            .I(N__13892));
    LocalMux I__1227 (
            .O(N__13892),
            .I(N__13889));
    Odrv4 I__1226 (
            .O(N__13889),
            .I(\pid_alt.O_21 ));
    InMux I__1225 (
            .O(N__13886),
            .I(N__13883));
    LocalMux I__1224 (
            .O(N__13883),
            .I(N__13880));
    Odrv4 I__1223 (
            .O(N__13880),
            .I(\pid_alt.O_22 ));
    InMux I__1222 (
            .O(N__13877),
            .I(N__13874));
    LocalMux I__1221 (
            .O(N__13874),
            .I(\pid_alt.O_6 ));
    InMux I__1220 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__1219 (
            .O(N__13868),
            .I(N__13865));
    Odrv4 I__1218 (
            .O(N__13865),
            .I(\pid_alt.O_24 ));
    InMux I__1217 (
            .O(N__13862),
            .I(N__13859));
    LocalMux I__1216 (
            .O(N__13859),
            .I(\pid_alt.O_15 ));
    CascadeMux I__1215 (
            .O(N__13856),
            .I(N__13853));
    InMux I__1214 (
            .O(N__13853),
            .I(N__13847));
    InMux I__1213 (
            .O(N__13852),
            .I(N__13847));
    LocalMux I__1212 (
            .O(N__13847),
            .I(N__13844));
    Span4Mux_v I__1211 (
            .O(N__13844),
            .I(N__13841));
    Odrv4 I__1210 (
            .O(N__13841),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    CascadeMux I__1209 (
            .O(N__13838),
            .I(\pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_ ));
    InMux I__1208 (
            .O(N__13835),
            .I(N__13829));
    InMux I__1207 (
            .O(N__13834),
            .I(N__13829));
    LocalMux I__1206 (
            .O(N__13829),
            .I(N__13826));
    Odrv12 I__1205 (
            .O(N__13826),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__1204 (
            .O(N__13823),
            .I(N__13820));
    LocalMux I__1203 (
            .O(N__13820),
            .I(N__13817));
    Span4Mux_h I__1202 (
            .O(N__13817),
            .I(N__13814));
    Odrv4 I__1201 (
            .O(N__13814),
            .I(\pid_alt.O_18 ));
    InMux I__1200 (
            .O(N__13811),
            .I(N__13804));
    InMux I__1199 (
            .O(N__13810),
            .I(N__13804));
    InMux I__1198 (
            .O(N__13809),
            .I(N__13801));
    LocalMux I__1197 (
            .O(N__13804),
            .I(N__13798));
    LocalMux I__1196 (
            .O(N__13801),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    Odrv4 I__1195 (
            .O(N__13798),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    InMux I__1194 (
            .O(N__13793),
            .I(N__13790));
    LocalMux I__1193 (
            .O(N__13790),
            .I(N__13787));
    Span4Mux_h I__1192 (
            .O(N__13787),
            .I(N__13784));
    Odrv4 I__1191 (
            .O(N__13784),
            .I(\pid_alt.O_23 ));
    InMux I__1190 (
            .O(N__13781),
            .I(N__13778));
    LocalMux I__1189 (
            .O(N__13778),
            .I(\pid_alt.O_4 ));
    InMux I__1188 (
            .O(N__13775),
            .I(N__13772));
    LocalMux I__1187 (
            .O(N__13772),
            .I(N__13769));
    Odrv4 I__1186 (
            .O(N__13769),
            .I(\pid_alt.O_17 ));
    InMux I__1185 (
            .O(N__13766),
            .I(N__13763));
    LocalMux I__1184 (
            .O(N__13763),
            .I(\pid_alt.O_0_13 ));
    InMux I__1183 (
            .O(N__13760),
            .I(N__13757));
    LocalMux I__1182 (
            .O(N__13757),
            .I(N__13754));
    Odrv4 I__1181 (
            .O(N__13754),
            .I(\pid_alt.O_0_24 ));
    InMux I__1180 (
            .O(N__13751),
            .I(N__13748));
    LocalMux I__1179 (
            .O(N__13748),
            .I(\pid_alt.O_0_19 ));
    InMux I__1178 (
            .O(N__13745),
            .I(N__13742));
    LocalMux I__1177 (
            .O(N__13742),
            .I(\pid_alt.O_0_20 ));
    InMux I__1176 (
            .O(N__13739),
            .I(N__13736));
    LocalMux I__1175 (
            .O(N__13736),
            .I(\pid_alt.O_0_18 ));
    InMux I__1174 (
            .O(N__13733),
            .I(N__13730));
    LocalMux I__1173 (
            .O(N__13730),
            .I(\pid_alt.O_0_9 ));
    CascadeMux I__1172 (
            .O(N__13727),
            .I(N__13722));
    InMux I__1171 (
            .O(N__13726),
            .I(N__13719));
    InMux I__1170 (
            .O(N__13725),
            .I(N__13714));
    InMux I__1169 (
            .O(N__13722),
            .I(N__13714));
    LocalMux I__1168 (
            .O(N__13719),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    LocalMux I__1167 (
            .O(N__13714),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__1166 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__1165 (
            .O(N__13706),
            .I(N__13703));
    Odrv4 I__1164 (
            .O(N__13703),
            .I(\pid_alt.O_0_17 ));
    InMux I__1163 (
            .O(N__13700),
            .I(N__13697));
    LocalMux I__1162 (
            .O(N__13697),
            .I(\pid_alt.O_0_15 ));
    InMux I__1161 (
            .O(N__13694),
            .I(N__13691));
    LocalMux I__1160 (
            .O(N__13691),
            .I(N__13688));
    Odrv4 I__1159 (
            .O(N__13688),
            .I(\pid_alt.O_0_16 ));
    InMux I__1158 (
            .O(N__13685),
            .I(N__13682));
    LocalMux I__1157 (
            .O(N__13682),
            .I(\pid_alt.O_0_5 ));
    InMux I__1156 (
            .O(N__13679),
            .I(N__13676));
    LocalMux I__1155 (
            .O(N__13676),
            .I(N__13673));
    Odrv4 I__1154 (
            .O(N__13673),
            .I(\pid_alt.O_0_22 ));
    InMux I__1153 (
            .O(N__13670),
            .I(N__13667));
    LocalMux I__1152 (
            .O(N__13667),
            .I(\pid_alt.O_0_4 ));
    InMux I__1151 (
            .O(N__13664),
            .I(N__13661));
    LocalMux I__1150 (
            .O(N__13661),
            .I(\pid_alt.O_0_10 ));
    InMux I__1149 (
            .O(N__13658),
            .I(N__13655));
    LocalMux I__1148 (
            .O(N__13655),
            .I(\pid_alt.O_0_23 ));
    InMux I__1147 (
            .O(N__13652),
            .I(N__13649));
    LocalMux I__1146 (
            .O(N__13649),
            .I(\pid_alt.O_0_11 ));
    InMux I__1145 (
            .O(N__13646),
            .I(N__13643));
    LocalMux I__1144 (
            .O(N__13643),
            .I(N__13640));
    Odrv4 I__1143 (
            .O(N__13640),
            .I(\pid_alt.O_0_6 ));
    InMux I__1142 (
            .O(N__13637),
            .I(N__13634));
    LocalMux I__1141 (
            .O(N__13634),
            .I(N__13631));
    Odrv4 I__1140 (
            .O(N__13631),
            .I(\pid_alt.O_0_14 ));
    InMux I__1139 (
            .O(N__13628),
            .I(N__13625));
    LocalMux I__1138 (
            .O(N__13625),
            .I(N__13622));
    Odrv4 I__1137 (
            .O(N__13622),
            .I(\pid_alt.O_0_12 ));
    InMux I__1136 (
            .O(N__13619),
            .I(N__13616));
    LocalMux I__1135 (
            .O(N__13616),
            .I(N__13613));
    Odrv4 I__1134 (
            .O(N__13613),
            .I(\pid_alt.O_0_21 ));
    InMux I__1133 (
            .O(N__13610),
            .I(N__13607));
    LocalMux I__1132 (
            .O(N__13607),
            .I(\pid_alt.O_0_7 ));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\scaler_3.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(\scaler_3.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\scaler_2.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(\scaler_2.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_5_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_29_0_));
    defparam IN_MUX_bfv_5_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_5_30_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_13 ),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_3_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_22_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_13 ),
            .carryinitout(bfn_3_22_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_2_27_0_));
    defparam IN_MUX_bfv_2_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_28_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_5_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_28_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_5_28_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_11_16_0_));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__26141),
            .GLOBALBUFFEROUTPUT(N_423_g));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__35079),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__21494),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_422_0_g ));
    ICE_GB debug_CH3_20A_c_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__36377),
            .GLOBALBUFFEROUTPUT(debug_CH3_20A_c_0_g));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34076),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__25313),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_320_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_2_LC_1_3_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13646),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36167),
            .ce(N__20312),
            .sr(N__21582));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_4_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13637),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36166),
            .ce(N__20311),
            .sr(N__21581));
    defparam \pid_alt.error_p_reg_esr_8_LC_1_4_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13628),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36166),
            .ce(N__20311),
            .sr(N__21581));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_4_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13619),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36166),
            .ce(N__20311),
            .sr(N__21581));
    defparam \pid_alt.error_p_reg_esr_3_LC_1_4_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13610),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36166),
            .ce(N__20311),
            .sr(N__21581));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_5_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13709),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_5_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13700),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13694),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_1_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13685),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13679),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_0_LC_1_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13670),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36165),
            .ce(N__20310),
            .sr(N__21580));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13664),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13658),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13652),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13766),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13760),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13751),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_6_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13745),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_6_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13739),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36163),
            .ce(N__20308),
            .sr(N__21578));
    defparam \pid_alt.error_p_reg_esr_RNIC74E2_5_LC_1_7_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIC74E2_5_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIC74E2_5_LC_1_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIC74E2_5_LC_1_7_0  (
            .in0(N__17377),
            .in1(N__17416),
            .in2(N__15416),
            .in3(N__14191),
            .lcout(\pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_5_LC_1_7_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13733),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36161),
            .ce(N__20307),
            .sr(N__21577));
    defparam \pid_alt.error_p_reg_esr_RNIGQ581_14_LC_1_7_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIGQ581_14_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIGQ581_14_LC_1_7_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIGQ581_14_LC_1_7_4  (
            .in0(N__13809),
            .in1(N__18370),
            .in2(N__13727),
            .in3(N__18143),
            .lcout(\pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI9U2K_15_LC_1_7_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI9U2K_15_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI9U2K_15_LC_1_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI9U2K_15_LC_1_7_6  (
            .in0(N__13725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18371),
            .lcout(\pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIKU581_15_LC_1_7_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIKU581_15_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIKU581_15_LC_1_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIKU581_15_LC_1_7_7  (
            .in0(N__13726),
            .in1(N__18489),
            .in2(N__18381),
            .in3(N__18525),
            .lcout(\pid_alt.error_p_reg_esr_RNIKU581Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI6JDH1_13_LC_1_8_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI6JDH1_13_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI6JDH1_13_LC_1_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI6JDH1_13_LC_1_8_2  (
            .in0(N__13834),
            .in1(N__17710),
            .in2(N__15613),
            .in3(N__17746),
            .lcout(\pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_0_14_LC_1_8_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_0_14_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_0_14_LC_1_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI7S2K_0_14_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__18133),
            .in2(_gnd_net_),
            .in3(N__13810),
            .lcout(\pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14 ),
            .ltout(\pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI0R7B1_13_LC_1_8_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI0R7B1_13_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI0R7B1_13_LC_1_8_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI0R7B1_13_LC_1_8_5  (
            .in0(N__17747),
            .in1(N__17709),
            .in2(N__13838),
            .in3(N__13835),
            .lcout(\pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_8_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13823),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36157),
            .ce(N__20306),
            .sr(N__21576));
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_14_LC_1_8_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_14_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI7S2K_14_LC_1_8_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI7S2K_14_LC_1_8_7  (
            .in0(N__13811),
            .in1(_gnd_net_),
            .in2(N__18144),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIH63K_19_LC_1_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIH63K_19_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIH63K_19_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIH63K_19_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__18585),
            .in2(_gnd_net_),
            .in3(N__14172),
            .lcout(\pid_alt.error_p_reg_esr_RNIH63KZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_9_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13793),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36154),
            .ce(N__20305),
            .sr(N__21575));
    defparam \pid_alt.error_i_reg_esr_0_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13781),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13775),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13913),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13904),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13895),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13886),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_2_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13877),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13871),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36151),
            .ce(N__20304),
            .sr(N__21574));
    defparam \pid_alt.error_p_reg_esr_RNIHVGK1_11_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIHVGK1_11_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIHVGK1_11_LC_1_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIHVGK1_11_LC_1_11_0  (
            .in0(N__15700),
            .in1(N__13852),
            .in2(N__17893),
            .in3(N__17907),
            .lcout(\pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13862),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36147),
            .ce(N__20302),
            .sr(N__21572));
    defparam \pid_alt.error_p_reg_esr_RNIAH8Q_11_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIAH8Q_11_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIAH8Q_11_LC_1_11_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIAH8Q_11_LC_1_11_3  (
            .in0(N__17908),
            .in1(_gnd_net_),
            .in2(N__13856),
            .in3(N__17888),
            .lcout(\pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11 ),
            .ltout(\pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIN5HK1_12_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIN5HK1_12_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIN5HK1_12_LC_1_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIN5HK1_12_LC_1_11_4  (
            .in0(N__13969),
            .in1(N__17807),
            .in2(N__13979),
            .in3(N__17826),
            .lcout(\pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13976),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36147),
            .ce(N__20302),
            .sr(N__21572));
    defparam \pid_alt.error_p_reg_esr_RNIDK8Q_12_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIDK8Q_12_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIDK8Q_12_LC_1_11_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIDK8Q_12_LC_1_11_6  (
            .in0(N__13970),
            .in1(N__17808),
            .in2(_gnd_net_),
            .in3(N__17827),
            .lcout(\pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIM0S12_10_LC_1_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIM0S12_10_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIM0S12_10_LC_1_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIM0S12_10_LC_1_12_0  (
            .in0(N__17966),
            .in1(N__17985),
            .in2(N__15755),
            .in3(N__13948),
            .lcout(\pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13955),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36144),
            .ce(N__20301),
            .sr(N__21571));
    defparam \pid_alt.error_p_reg_esr_RNI7E8Q_10_LC_1_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI7E8Q_10_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI7E8Q_10_LC_1_12_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI7E8Q_10_LC_1_12_2  (
            .in0(N__17967),
            .in1(N__13949),
            .in2(_gnd_net_),
            .in3(N__17986),
            .lcout(\pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIO2681_16_LC_1_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIO2681_16_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIO2681_16_LC_1_12_4 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIO2681_16_LC_1_12_4  (
            .in0(N__18860),
            .in1(N__14044),
            .in2(N__18498),
            .in3(N__18539),
            .lcout(\pid_alt.error_p_reg_esr_RNIO2681Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNID23K_17_LC_1_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNID23K_17_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNID23K_17_LC_1_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNID23K_17_LC_1_12_6  (
            .in0(N__18861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14043),
            .lcout(\pid_alt.error_p_reg_esr_RNID23KZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13937),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36140),
            .ce(N__20299),
            .sr(N__21569));
    defparam \pid_alt.error_i_reg_esr_3_LC_1_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13925),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36140),
            .ce(N__20299),
            .sr(N__21569));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13997),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36140),
            .ce(N__20299),
            .sr(N__21569));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13988),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36140),
            .ce(N__20299),
            .sr(N__21569));
    defparam \pid_alt.error_i_acumm_10_LC_1_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_1_14_0 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_1_14_0  (
            .in0(N__15325),
            .in1(N__23950),
            .in2(N__17971),
            .in3(N__17939),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_11_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_1_14_1 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_1_14_1  (
            .in0(N__23947),
            .in1(N__15328),
            .in2(N__17892),
            .in3(N__17858),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_6_LC_1_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_1_14_2 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_1_14_2  (
            .in0(N__15326),
            .in1(N__23951),
            .in2(N__20397),
            .in3(N__17303),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_9_LC_1_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_1_14_3 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_1_14_3  (
            .in0(N__23949),
            .in1(N__15329),
            .in2(N__18050),
            .in3(N__18014),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_8_LC_1_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_1_14_4 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_1_14_4  (
            .in0(N__15327),
            .in1(N__23952),
            .in2(N__17225),
            .in3(N__17192),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_12_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_1_14_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_1_14_6  (
            .in0(N__17776),
            .in1(N__15269),
            .in2(N__17812),
            .in3(N__23953),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_5_LC_1_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_1_14_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_1_14_7  (
            .in0(N__23948),
            .in1(N__17344),
            .in2(N__17415),
            .in3(N__14125),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36135),
            .ce(),
            .sr(N__15216));
    defparam \pid_alt.error_i_acumm_esr_3_LC_1_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_1_15_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_1_15_0  (
            .in0(N__14126),
            .in1(N__14102),
            .in2(N__17470),
            .in3(N__17540),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36131),
            .ce(N__15170),
            .sr(N__15217));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6M6T3_10_LC_1_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6M6T3_10_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6M6T3_10_LC_1_15_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI6M6T3_10_LC_1_15_1  (
            .in0(N__15095),
            .in1(N__15261),
            .in2(N__15065),
            .in3(N__15305),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(\pid_alt.N_62_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_4_LC_1_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_1_15_2 .LUT_INIT=16'b1111111100011101;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_1_15_2  (
            .in0(N__15306),
            .in1(N__17345),
            .in2(N__14027),
            .in3(N__17464),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36131),
            .ce(N__15170),
            .sr(N__15217));
    defparam \pid_alt.error_p_reg_esr_RNI6UG61_3_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI6UG61_3_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI6UG61_3_LC_1_15_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI6UG61_3_LC_1_15_3  (
            .in0(N__17587),
            .in1(_gnd_net_),
            .in2(N__17560),
            .in3(N__14021),
            .lcout(\pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3 ),
            .ltout(\pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIFV1D2_4_LC_1_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIFV1D2_4_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIFV1D2_4_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIFV1D2_4_LC_1_15_4  (
            .in0(N__14500),
            .in1(N__17490),
            .in2(N__14024),
            .in3(N__17511),
            .lcout(\pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI91H61_4_LC_1_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI91H61_4_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI91H61_4_LC_1_15_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI91H61_4_LC_1_15_5  (
            .in0(N__17512),
            .in1(_gnd_net_),
            .in2(N__17497),
            .in3(N__14501),
            .lcout(\pid_alt.error_p_reg_esr_RNI91H61Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI9P1D2_3_LC_1_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI9P1D2_3_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI9P1D2_3_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI9P1D2_3_LC_1_15_6  (
            .in0(N__14020),
            .in1(N__17553),
            .in2(N__15488),
            .in3(N__17586),
            .lcout(\pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0_5_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0_5_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0_5_LC_1_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0_5_LC_1_15_7  (
            .in0(N__15094),
            .in1(N__17343),
            .in2(N__15064),
            .in3(N__15260),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_1_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_1_16_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_1_16_0  (
            .in0(N__17466),
            .in1(N__14128),
            .in2(N__17081),
            .in3(N__14100),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36125),
            .ce(N__15159),
            .sr(N__15212));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNISKMM7_5_LC_1_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNISKMM7_5_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNISKMM7_5_LC_1_16_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNISKMM7_5_LC_1_16_1  (
            .in0(N__15077),
            .in1(N__14003),
            .in2(_gnd_net_),
            .in3(N__15304),
            .lcout(\pid_alt.N_37 ),
            .ltout(\pid_alt.N_37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_1_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_1_16_2 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_1_16_2  (
            .in0(N__18202),
            .in1(N__14127),
            .in2(N__14132),
            .in3(N__17465),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36125),
            .ce(N__15159),
            .sr(N__15212));
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_0_1_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_0_1_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_0_1_LC_1_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI0OG61_0_1_LC_1_16_3  (
            .in0(N__17118),
            .in1(N__14086),
            .in2(_gnd_net_),
            .in3(N__17100),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_2_LC_1_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_1_16_4 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_1_16_4  (
            .in0(N__14129),
            .in1(N__14101),
            .in2(N__17471),
            .in3(N__17609),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36125),
            .ce(N__15159),
            .sr(N__15212));
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_1_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_1_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI0OG61_1_LC_1_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI0OG61_1_LC_1_16_5  (
            .in0(N__17119),
            .in1(N__14087),
            .in2(_gnd_net_),
            .in3(N__17101),
            .lcout(\pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1 ),
            .ltout(\pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3J1D2_2_LC_1_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3J1D2_2_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3J1D2_2_LC_1_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3J1D2_2_LC_1_16_6  (
            .in0(N__14071),
            .in1(N__17622),
            .in2(N__14075),
            .in3(N__17655),
            .lcout(\pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3RG61_2_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3RG61_2_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3RG61_2_LC_1_16_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3RG61_2_LC_1_16_7  (
            .in0(N__17656),
            .in1(_gnd_net_),
            .in2(N__17629),
            .in3(N__14072),
            .lcout(\pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI2G981_20_LC_1_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI2G981_20_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI2G981_20_LC_1_17_0 .LUT_INIT=16'b0111011101111000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI2G981_20_LC_1_17_0  (
            .in0(N__20789),
            .in1(N__20844),
            .in2(N__20799),
            .in3(N__20846),
            .lcout(\pid_alt.error_p_reg_esr_RNI2G981Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIS6681_17_LC_1_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIS6681_17_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIS6681_17_LC_1_17_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIS6681_17_LC_1_17_1  (
            .in0(N__18870),
            .in1(N__20581),
            .in2(N__14054),
            .in3(N__20620),
            .lcout(\pid_alt.error_p_reg_esr_RNIS6681Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIIU781_19_LC_1_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIIU781_19_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIIU781_19_LC_1_17_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIIU781_19_LC_1_17_2  (
            .in0(N__20788),
            .in1(N__18597),
            .in2(N__14177),
            .in3(N__20845),
            .lcout(\pid_alt.error_p_reg_esr_RNIIU781Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI36J71_5_LC_1_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI36J71_5_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI36J71_5_LC_1_17_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI36J71_5_LC_1_17_3  (
            .in0(N__14195),
            .in1(N__17373),
            .in2(_gnd_net_),
            .in3(N__17411),
            .lcout(\pid_alt.error_p_reg_esr_RNI36J71Z0Z_5 ),
            .ltout(\pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI9F6F2_6_LC_1_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI9F6F2_6_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI9F6F2_6_LC_1_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI9F6F2_6_LC_1_17_4  (
            .in0(N__20434),
            .in1(N__20458),
            .in2(N__14180),
            .in3(N__20390),
            .lcout(\pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI0B681_18_LC_1_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI0B681_18_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI0B681_18_LC_1_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI0B681_18_LC_1_17_6  (
            .in0(N__20621),
            .in1(N__14173),
            .in2(N__20585),
            .in3(N__18596),
            .lcout(\pid_alt.error_p_reg_esr_RNI0B681Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_18_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__31493),
            .in2(_gnd_net_),
            .in3(N__21625),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36115),
            .ce(N__28049),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_5_LC_1_19_3 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_5_LC_1_19_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_5_LC_1_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.source_data_1_esr_5_LC_1_19_3  (
            .in0(N__23780),
            .in1(N__23818),
            .in2(_gnd_net_),
            .in3(N__21041),
            .lcout(scaler_2_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36109),
            .ce(N__29572),
            .sr(N__36739));
    defparam \pid_alt.source_pid_1_10_LC_1_20_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_1_20_0 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \pid_alt.source_pid_1_10_LC_1_20_0  (
            .in0(N__18659),
            .in1(N__18802),
            .in2(N__21415),
            .in3(N__23939),
            .lcout(throttle_command_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(),
            .sr(N__19260));
    defparam \pid_alt.source_pid_1_11_LC_1_20_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_1_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_1_20_1 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \pid_alt.source_pid_1_11_LC_1_20_1  (
            .in0(N__18803),
            .in1(N__18761),
            .in2(N__23954),
            .in3(N__16107),
            .lcout(throttle_command_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(),
            .sr(N__19260));
    defparam \pid_alt.source_pid_1_7_LC_1_20_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_1_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_1_20_4 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \pid_alt.source_pid_1_7_LC_1_20_4  (
            .in0(N__18641),
            .in1(N__18805),
            .in2(N__16187),
            .in3(N__23940),
            .lcout(throttle_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(),
            .sr(N__19260));
    defparam \pid_alt.source_pid_1_6_LC_1_20_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_1_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_1_20_5 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \pid_alt.source_pid_1_6_LC_1_20_5  (
            .in0(N__18804),
            .in1(N__18710),
            .in2(N__23955),
            .in3(N__14263),
            .lcout(throttle_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(),
            .sr(N__19260));
    defparam \pid_alt.source_pid_1_9_LC_1_20_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_1_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_1_20_7 .LUT_INIT=16'b1110111001001110;
    LogicCell40 \pid_alt.source_pid_1_9_LC_1_20_7  (
            .in0(N__23932),
            .in1(N__14406),
            .in2(N__18809),
            .in3(N__18737),
            .lcout(throttle_command_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36103),
            .ce(),
            .sr(N__19260));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_1_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_1_21_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_14_LC_1_21_0  (
            .in0(N__24300),
            .in1(N__23089),
            .in2(_gnd_net_),
            .in3(N__30099),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_1_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_1_21_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_1_21_2  (
            .in0(N__29426),
            .in1(N__14345),
            .in2(_gnd_net_),
            .in3(N__24407),
            .lcout(\ppm_encoder_1.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_5_LC_1_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_1_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_1_21_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_1_21_3  (
            .in0(N__24972),
            .in1(N__15989),
            .in2(N__14306),
            .in3(N__14201),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36096),
            .ce(),
            .sr(N__36750));
    defparam \ppm_encoder_1.throttle_6_LC_1_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_1_21_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_1_21_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_1_21_4  (
            .in0(N__14243),
            .in1(N__14262),
            .in2(N__29329),
            .in3(N__24973),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36096),
            .ce(),
            .sr(N__36750));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_1_22_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_1_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(N__24526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_1_22_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_1_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(N__25069),
            .in2(N__28567),
            .in3(N__14213),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_1_22_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_1_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(N__21322),
            .in2(_gnd_net_),
            .in3(N__14210),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_1_22_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_1_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__25021),
            .in2(N__28568),
            .in3(N__14207),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_1_22_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(N__21811),
            .in2(_gnd_net_),
            .in3(N__14204),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_1_22_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(N__15985),
            .in2(_gnd_net_),
            .in3(N__14267),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_1_22_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_1_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(N__14264),
            .in2(N__28569),
            .in3(N__14237),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_1_22_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_1_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(N__16182),
            .in2(_gnd_net_),
            .in3(N__14234),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_1_23_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_1_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(N__21922),
            .in2(_gnd_net_),
            .in3(N__14231),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_1_23_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(N__14407),
            .in2(_gnd_net_),
            .in3(N__14228),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_1_23_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_1_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__21411),
            .in2(_gnd_net_),
            .in3(N__14225),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_1_23_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_1_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_1_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(N__16108),
            .in2(_gnd_net_),
            .in3(N__14222),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_1_23_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(N__21685),
            .in2(_gnd_net_),
            .in3(N__14219),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_1_23_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_1_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(N__21370),
            .in2(N__28535),
            .in3(N__14216),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_1_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14312),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36081),
            .ce(N__27302),
            .sr(N__36757));
    defparam CONSTANT_ONE_LUT4_LC_1_23_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_23_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_23_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_1_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_1_24_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_1_24_0  (
            .in0(N__14304),
            .in1(N__27319),
            .in2(N__22361),
            .in3(N__22262),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_1_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_1_24_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_1_24_1  (
            .in0(N__16432),
            .in1(_gnd_net_),
            .in2(N__14309),
            .in3(N__16262),
            .lcout(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_1_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_1_24_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_1_24_3  (
            .in0(N__14305),
            .in1(N__16274),
            .in2(_gnd_net_),
            .in3(N__22500),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_1_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_1_24_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(N__29237),
            .in2(N__14282),
            .in3(N__16286),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_5_LC_1_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_5_LC_1_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_5_LC_1_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_5_LC_1_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14279),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36072),
            .ce(N__27294),
            .sr(N__36759));
    defparam \ppm_encoder_1.elevator_esr_5_LC_1_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_5_LC_1_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_5_LC_1_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_5_LC_1_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29588),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36072),
            .ce(N__27294),
            .sr(N__36759));
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_1_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_1_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_1_24_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_1_24_7  (
            .in0(N__24403),
            .in1(N__19052),
            .in2(N__22125),
            .in3(N__22026),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_1_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_1_25_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNIU0DH2_10_LC_1_25_0  (
            .in0(N__24160),
            .in1(N__24103),
            .in2(N__22130),
            .in3(N__22030),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_1_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_1_25_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI5GRT5_10_LC_1_25_1  (
            .in0(_gnd_net_),
            .in1(N__19616),
            .in2(N__14354),
            .in3(N__14351),
            .lcout(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_1_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_1_25_2 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIE2JI2_10_LC_1_25_2  (
            .in0(N__22606),
            .in1(N__25456),
            .in2(N__22264),
            .in3(N__22353),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_1_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_1_25_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_1_25_3  (
            .in0(N__22354),
            .in1(N__14344),
            .in2(N__25784),
            .in3(N__22256),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_1_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_1_25_4 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_1_25_4  (
            .in0(N__16552),
            .in1(_gnd_net_),
            .in2(N__14327),
            .in3(N__14324),
            .lcout(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_1_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_1_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_1_25_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIN3352_0_LC_1_25_5  (
            .in0(_gnd_net_),
            .in1(N__24514),
            .in2(N__19838),
            .in3(N__22252),
            .lcout(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_1_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_1_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_1_25_6 .LUT_INIT=16'b0110001101100011;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_1_25_6  (
            .in0(N__24515),
            .in1(N__19833),
            .in2(N__22265),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_1_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_1_25_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_1_25_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_1_25_7  (
            .in0(N__23230),
            .in1(N__19664),
            .in2(N__14318),
            .in3(N__20121),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36062),
            .ce(),
            .sr(N__36762));
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_1_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_1_26_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNIEMVN2_9_LC_1_26_0  (
            .in0(N__14433),
            .in1(N__23421),
            .in2(N__22031),
            .in3(N__22129),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_1_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_1_26_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNITSI96_9_LC_1_26_1  (
            .in0(N__19577),
            .in1(_gnd_net_),
            .in2(N__14315),
            .in3(N__14441),
            .lcout(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_1_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_1_26_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIU7KK2_9_LC_1_26_2  (
            .in0(N__14382),
            .in1(N__14367),
            .in2(N__22360),
            .in3(N__22260),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_1_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_1_26_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_1_26_3  (
            .in0(N__29483),
            .in1(N__14383),
            .in2(_gnd_net_),
            .in3(N__14434),
            .lcout(\ppm_encoder_1.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_9_LC_1_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_1_26_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_1_26_4 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_1_26_4  (
            .in0(N__24991),
            .in1(N__14435),
            .in2(N__24467),
            .in3(N__28907),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36055),
            .ce(),
            .sr(N__36766));
    defparam \ppm_encoder_1.throttle_9_LC_1_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_1_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_1_26_5 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_1_26_5  (
            .in0(N__24996),
            .in1(N__14420),
            .in2(N__14387),
            .in3(N__14411),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36055),
            .ce(),
            .sr(N__36766));
    defparam \ppm_encoder_1.aileron_9_LC_1_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_1_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_1_26_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_1_26_6  (
            .in0(N__19091),
            .in1(N__20915),
            .in2(N__25001),
            .in3(N__23422),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36055),
            .ce(),
            .sr(N__36766));
    defparam \ppm_encoder_1.rudder_9_LC_1_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_1_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_1_26_7 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_1_26_7  (
            .in0(N__14368),
            .in1(N__24992),
            .in2(N__25559),
            .in3(N__26477),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36055),
            .ce(),
            .sr(N__36766));
    defparam \ppm_encoder_1.init_pulses_9_LC_1_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_1_27_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_1_27_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_1_27_0  (
            .in0(N__20108),
            .in1(N__23237),
            .in2(N__16361),
            .in3(N__16709),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36048),
            .ce(),
            .sr(N__36769));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_1_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_1_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_1_27_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_1_27_1  (
            .in0(N__19596),
            .in1(N__23059),
            .in2(_gnd_net_),
            .in3(N__30048),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_1_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_1_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_1_27_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_1_27_3  (
            .in0(N__19597),
            .in1(N__27957),
            .in2(N__30583),
            .in3(N__14369),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_1_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_1_27_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_1_27_4  (
            .in0(N__30047),
            .in1(_gnd_net_),
            .in2(N__23085),
            .in3(N__20008),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_1_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_1_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_1_27_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_1_27_5  (
            .in0(N__20007),
            .in1(N__23055),
            .in2(_gnd_net_),
            .in3(N__30046),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_1_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_1_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_1_27_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_1_27_6  (
            .in0(N__27956),
            .in1(N__20009),
            .in2(N__27326),
            .in3(N__30575),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_1_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_1_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_1_27_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_1_27_7  (
            .in0(N__24259),
            .in1(N__23060),
            .in2(_gnd_net_),
            .in3(N__30049),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_1_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_1_28_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_1_28_0  (
            .in0(N__23288),
            .in1(N__24580),
            .in2(N__30089),
            .in3(N__19945),
            .lcout(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_1_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_1_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_1_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_1_28_1  (
            .in0(_gnd_net_),
            .in1(N__23284),
            .in2(_gnd_net_),
            .in3(N__30051),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_1_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_1_28_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_1_28_2  (
            .in0(N__30052),
            .in1(_gnd_net_),
            .in2(N__23296),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_1_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_1_28_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_1_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30050),
            .lcout(\ppm_encoder_1.N_1014_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_17_LC_1_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_1_28_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_1_28_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_1_28_6  (
            .in0(N__23236),
            .in1(N__20083),
            .in2(N__16472),
            .in3(N__16793),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36041),
            .ce(),
            .sr(N__36771));
    defparam \ppm_encoder_1.init_pulses_14_LC_1_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_1_28_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_1_28_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_1_28_7  (
            .in0(N__20082),
            .in1(N__23235),
            .in2(N__16532),
            .in3(N__16832),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36041),
            .ce(),
            .sr(N__36771));
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_1_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_1_29_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_1_29_0  (
            .in0(N__25298),
            .in1(N__22417),
            .in2(N__22505),
            .in3(N__25362),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_1_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_1_29_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_1_29_1  (
            .in0(N__25397),
            .in1(_gnd_net_),
            .in2(N__14447),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_1_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_1_29_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_1_29_2 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_1_29_2  (
            .in0(N__23212),
            .in1(N__16643),
            .in2(N__14444),
            .in3(N__16250),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36032),
            .ce(),
            .sr(N__36772));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_1_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_1_29_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_1_29_3  (
            .in0(N__23361),
            .in1(N__23051),
            .in2(_gnd_net_),
            .in3(N__30044),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_1_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_1_29_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_1_29_4  (
            .in0(N__30045),
            .in1(_gnd_net_),
            .in2(N__23084),
            .in3(N__23362),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_1_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_1_29_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_1_29_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_1_29_5  (
            .in0(N__20071),
            .in1(N__16697),
            .in2(N__23231),
            .in3(N__16340),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36032),
            .ce(),
            .sr(N__36772));
    defparam \ppm_encoder_1.init_pulses_11_LC_1_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_1_29_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_1_29_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_1_29_6  (
            .in0(N__23211),
            .in1(N__20072),
            .in2(N__16316),
            .in3(N__16688),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36032),
            .ce(),
            .sr(N__36772));
    defparam \ppm_encoder_1.init_pulses_12_LC_1_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_1_29_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_1_29_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_1_29_7  (
            .in0(N__20073),
            .in1(N__16679),
            .in2(N__23232),
            .in3(N__16622),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36032),
            .ce(),
            .sr(N__36772));
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_1_30_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_1_30_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_1_30_0  (
            .in0(N__19946),
            .in1(N__23075),
            .in2(N__30101),
            .in3(N__30153),
            .lcout(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_1_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_1_30_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_1_30_1  (
            .in0(N__30154),
            .in1(N__23063),
            .in2(_gnd_net_),
            .in3(N__30092),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_1_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_1_30_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_1_30_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_1_30_2  (
            .in0(N__20101),
            .in1(N__16814),
            .in2(N__23234),
            .in3(N__16490),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36022),
            .ce(),
            .sr(N__36773));
    defparam \ppm_encoder_1.init_pulses_18_LC_1_30_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_1_30_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_1_30_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_1_30_4  (
            .in0(N__16778),
            .in1(N__20084),
            .in2(N__16457),
            .in3(N__23227),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36022),
            .ce(),
            .sr(N__36773));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_1_30_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_1_30_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_1_30_5  (
            .in0(_gnd_net_),
            .in1(N__23062),
            .in2(_gnd_net_),
            .in3(N__30091),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_1_30_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_1_30_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_1_30_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_1_30_6  (
            .in0(N__20100),
            .in1(N__16841),
            .in2(N__23233),
            .in3(N__16574),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36022),
            .ce(),
            .sr(N__36773));
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_1_30_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_1_30_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_1_30_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISFRP_13_LC_1_30_7  (
            .in0(N__24573),
            .in1(N__23061),
            .in2(_gnd_net_),
            .in3(N__30090),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_4_LC_2_5_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_2_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14513),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36164),
            .ce(N__20309),
            .sr(N__21579));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_7_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_7_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__30869),
            .in2(_gnd_net_),
            .in3(N__21633),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36158),
            .ce(N__25756),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_7_LC_2_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_2_8_0 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_2_8_0  (
            .in0(N__17279),
            .in1(N__15313),
            .in2(N__20222),
            .in3(N__23957),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36155),
            .ce(),
            .sr(N__15221));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_9_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_2_9_0  (
            .in0(N__31689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21629),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__31829),
            .in2(_gnd_net_),
            .in3(N__21626),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_9_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_2_9_3  (
            .in0(N__21627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30868),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_9_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__31220),
            .in2(_gnd_net_),
            .in3(N__21628),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_9_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_2_9_5  (
            .in0(N__21630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30745),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__31369),
            .in2(_gnd_net_),
            .in3(N__21631),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36152),
            .ce(N__28045),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNILR6F2_8_LC_2_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNILR6F2_8_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNILR6F2_8_LC_2_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNILR6F2_8_LC_2_10_0  (
            .in0(N__14543),
            .in1(N__17226),
            .in2(N__20191),
            .in3(N__17244),
            .lcout(\pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_2_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14555),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36148),
            .ce(N__20303),
            .sr(N__21573));
    defparam \pid_alt.error_p_reg_esr_RNICFJ71_8_LC_2_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNICFJ71_8_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNICFJ71_8_LC_2_10_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNICFJ71_8_LC_2_10_3  (
            .in0(N__17245),
            .in1(_gnd_net_),
            .in2(N__17231),
            .in3(N__14542),
            .lcout(\pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8 ),
            .ltout(\pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIR17F2_9_LC_2_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIR17F2_9_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIR17F2_9_LC_2_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIR17F2_9_LC_2_10_4  (
            .in0(N__14818),
            .in1(N__18047),
            .in2(N__14528),
            .in3(N__18063),
            .lcout(\pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_9_LC_2_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_2_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14525),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36148),
            .ce(N__20303),
            .sr(N__21573));
    defparam \pid_alt.error_p_reg_esr_RNIFIJ71_9_LC_2_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIFIJ71_9_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIFIJ71_9_LC_2_10_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIFIJ71_9_LC_2_10_6  (
            .in0(N__14819),
            .in1(N__18048),
            .in2(_gnd_net_),
            .in3(N__18064),
            .lcout(\pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_LC_2_11_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15116),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_11_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_2_11_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16997),
            .in3(N__14780),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_11_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17141),
            .in3(N__14753),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_11_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_2_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__14726),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_11_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__23495),
            .in2(N__17051),
            .in3(N__14696),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_11_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__23480),
            .in2(N__16892),
            .in3(N__14669),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_11_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__23465),
            .in2(N__16925),
            .in3(N__14639),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_11_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__16910),
            .in2(N__17036),
            .in3(N__14609),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_12_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_2_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__17021),
            .in2(N__23456),
            .in3(N__14999),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_12_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__17015),
            .in2(N__23591),
            .in3(N__14972),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_12_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__17009),
            .in2(N__23579),
            .in3(N__14945),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_12_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__17003),
            .in2(N__23567),
            .in3(N__14918),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_12_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_2_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__17171),
            .in2(_gnd_net_),
            .in3(N__14894),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_12_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_2_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__17159),
            .in2(_gnd_net_),
            .in3(N__14870),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_12_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_2_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__17147),
            .in2(_gnd_net_),
            .in3(N__14846),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_2_12_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__16937),
            .in2(_gnd_net_),
            .in3(N__14843),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_13_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_13_0  (
            .in0(N__17296),
            .in1(_gnd_net_),
            .in2(N__17275),
            .in3(_gnd_net_),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(\pid_alt.m35_e_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_5_LC_2_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_5_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_5_LC_2_13_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_5_LC_2_13_1  (
            .in0(N__17325),
            .in1(N__15049),
            .in2(N__15080),
            .in3(N__15268),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_2_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_2_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_2_13_2  (
            .in0(N__17188),
            .in1(N__17853),
            .in2(N__17938),
            .in3(N__18010),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_2_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_2_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__17931),
            .in2(_gnd_net_),
            .in3(N__17766),
            .lcout(),
            .ltout(\pid_alt.m21_e_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI56PT1_1_LC_2_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI56PT1_1_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI56PT1_1_LC_2_13_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI56PT1_1_LC_2_13_4  (
            .in0(N__17068),
            .in1(N__18203),
            .in2(N__15038),
            .in3(N__15032),
            .lcout(\pid_alt.m21_e_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_2_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_2_13_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_2_13_5  (
            .in0(N__17602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17533),
            .lcout(),
            .ltout(\pid_alt.m21_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_2_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_2_13_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_2_13_6  (
            .in0(N__17268),
            .in1(N__17324),
            .in2(N__15035),
            .in3(N__17436),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_2_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_2_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_2_13_7  (
            .in0(N__18009),
            .in1(N__17187),
            .in2(N__17857),
            .in3(N__17295),
            .lcout(\pid_alt.m21_e_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_14_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__23769),
            .in2(N__23817),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_2_14_1 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20738),
            .in2(N__23549),
            .in3(N__15026),
            .lcout(\scaler_2.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_0 ),
            .carryout(\scaler_2.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_2_14_2 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20729),
            .in2(N__23537),
            .in3(N__15140),
            .lcout(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_1 ),
            .carryout(\scaler_2.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_2_14_3 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__20720),
            .in2(N__23525),
            .in3(N__15137),
            .lcout(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_2 ),
            .carryout(\scaler_2.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_2_14_4 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__23513),
            .in2(N__20711),
            .in3(N__15134),
            .lcout(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_3 ),
            .carryout(\scaler_2.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_2_14_5 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__23669),
            .in2(N__20699),
            .in3(N__15131),
            .lcout(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_4 ),
            .carryout(\scaler_2.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_2_14_6 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__23660),
            .in2(N__20687),
            .in3(N__15128),
            .lcout(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_5 ),
            .carryout(\scaler_2.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_2_14_7 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_2_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__21062),
            .in2(_gnd_net_),
            .in3(N__15125),
            .lcout(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_6 ),
            .carryout(\scaler_2.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_2_15_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_2_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__21080),
            .in2(N__28690),
            .in3(N__15122),
            .lcout(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_15_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15119),
            .lcout(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_inv_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_2_15_2  (
            .in0(N__15109),
            .in1(N__28659),
            .in2(_gnd_net_),
            .in3(N__15345),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_15_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26125),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36126),
            .ce(N__25703),
            .sr(N__36717));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI24S01_12_LC_2_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI24S01_12_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI24S01_12_LC_2_16_0 .LUT_INIT=16'b1010111011101110;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI24S01_12_LC_2_16_0  (
            .in0(N__18320),
            .in1(N__15281),
            .in2(N__17780),
            .in3(N__17686),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_RNISOGT_14_LC_2_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_RNISOGT_14_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_RNISOGT_14_LC_2_16_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_RNISOGT_14_LC_2_16_1  (
            .in0(N__18413),
            .in1(N__18085),
            .in2(N__18559),
            .in3(N__18109),
            .lcout(\pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14 ),
            .ltout(\pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_13_LC_2_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_2_16_2 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__18318),
            .in2(N__15275),
            .in3(N__17687),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36121),
            .ce(N__15166),
            .sr(N__15208));
    defparam \pid_alt.error_i_acumm_prereg_RNINGKC_14_LC_2_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_RNINGKC_14_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_RNINGKC_14_LC_2_16_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_RNINGKC_14_LC_2_16_3  (
            .in0(N__18552),
            .in1(N__18084),
            .in2(_gnd_net_),
            .in3(N__18108),
            .lcout(),
            .ltout(\pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBMOV_13_LC_2_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBMOV_13_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBMOV_13_LC_2_16_4 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIBMOV_13_LC_2_16_4  (
            .in0(N__18319),
            .in1(N__17685),
            .in2(N__15272),
            .in3(N__18412),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(\pid_alt.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75_21_LC_2_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75_21_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75_21_LC_2_16_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75_21_LC_2_16_5  (
            .in0(N__18317),
            .in1(N__15245),
            .in2(N__15236),
            .in3(N__15233),
            .lcout(),
            .ltout(\pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNI2P1V5_1_LC_2_16_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNI2P1V5_1_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNI2P1V5_1_LC_2_16_6 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \pid_alt.state_RNI2P1V5_1_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__23912),
            .in2(N__15224),
            .in3(N__35080),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(\pid_alt.un1_reset_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNINE9D6_1_LC_2_16_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNINE9D6_1_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNINE9D6_1_LC_2_16_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_alt.state_RNINE9D6_1_LC_2_16_7  (
            .in0(N__23913),
            .in1(_gnd_net_),
            .in2(N__15173),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_60_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_2_17_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_2_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__15535),
            .in2(N__15542),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_2_17_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_2_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_2_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__18264),
            .in2(N__18248),
            .in3(N__15512),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.un1_pid_prereg_0_cry_0_THRU_LUT4_0_LC_2_17_2 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_0_cry_0_THRU_LUT4_0_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_0_cry_0_THRU_LUT4_0_LC_2_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_pid_prereg_0_cry_0_THRU_LUT4_0_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__21130),
            .in2(_gnd_net_),
            .in3(N__15509),
            .lcout(\pid_alt.un1_pid_prereg_0_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_2_LC_2_17_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_2_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_2_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__15506),
            .in2(N__15500),
            .in3(N__15491),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.pid_prereg_esr_3_LC_2_17_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__15484),
            .in2(N__15473),
            .in3(N__15461),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.pid_prereg_esr_4_LC_2_17_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_2_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__15458),
            .in2(N__15449),
            .in3(N__15434),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.pid_prereg_esr_5_LC_2_17_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_2_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_2_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__15431),
            .in2(N__15409),
            .in3(N__15386),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.pid_prereg_esr_6_LC_2_17_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_2_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_2_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__15383),
            .in2(N__15374),
            .in3(N__15365),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__36116),
            .ce(N__18297),
            .sr(N__36726));
    defparam \pid_alt.pid_prereg_esr_7_LC_2_18_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_2_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_2_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__20339),
            .in2(N__20360),
            .in3(N__15800),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_8_LC_2_18_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_2_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__15797),
            .in2(N__20192),
            .in3(N__15788),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_9_LC_2_18_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_2_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__15785),
            .in2(N__15776),
            .in3(N__15758),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_10_LC_2_18_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_2_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_2_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__15754),
            .in2(N__15725),
            .in3(N__15710),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_11_LC_2_18_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_2_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__15707),
            .in2(N__15686),
            .in3(N__15668),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_12_LC_2_18_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_2_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__15665),
            .in2(N__15650),
            .in3(N__15635),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_13_LC_2_18_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_2_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_2_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__15632),
            .in2(N__15614),
            .in3(N__15584),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_14_LC_2_18_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_2_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__15581),
            .in2(N__15566),
            .in3(N__15545),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__36110),
            .ce(N__18298),
            .sr(N__36729));
    defparam \pid_alt.pid_prereg_esr_15_LC_2_19_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_2_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__15974),
            .in2(N__15962),
            .in3(N__15944),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_16_LC_2_19_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_2_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__15941),
            .in2(N__15926),
            .in3(N__15911),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_17_LC_2_19_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_2_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__15908),
            .in2(N__18461),
            .in3(N__15896),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_18_LC_2_19_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_2_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_2_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__15893),
            .in2(N__15878),
            .in3(N__15866),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_19_LC_2_19_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_2_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__20552),
            .in2(N__15863),
            .in3(N__15851),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_20_LC_2_19_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_2_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__15848),
            .in2(N__15836),
            .in3(N__15818),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_21_LC_2_19_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_2_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_2_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__15815),
            .in2(N__20756),
            .in3(N__15806),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_22_LC_2_19_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_22_LC_2_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_2_19_7 .LUT_INIT=16'b0001000111101110;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_2_19_7  (
            .in0(N__20882),
            .in1(N__20810),
            .in2(_gnd_net_),
            .in3(N__15803),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36104),
            .ce(N__18299),
            .sr(N__36735));
    defparam \pid_alt.pid_prereg_esr_RNI8OUM_14_LC_2_20_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI8OUM_14_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI8OUM_14_LC_2_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI8OUM_14_LC_2_20_0  (
            .in0(N__16064),
            .in1(N__16055),
            .in2(N__16049),
            .in3(N__16040),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIQORD1_15_LC_2_20_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIQORD1_15_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIQORD1_15_LC_2_20_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIQORD1_15_LC_2_20_1  (
            .in0(N__16034),
            .in1(N__16028),
            .in2(N__16022),
            .in3(N__16004),
            .lcout(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15 ),
            .ltout(\pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_2_20_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_2_20_2 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \pid_alt.source_pid_1_esr_RNO_0_4_LC_2_20_2  (
            .in0(N__19398),
            .in1(N__19488),
            .in2(N__16019),
            .in3(N__19165),
            .lcout(\pid_alt.source_pid_9_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIBIEB_17_LC_2_20_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIBIEB_17_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIBIEB_17_LC_2_20_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIBIEB_17_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__16016),
            .in2(_gnd_net_),
            .in3(N__16010),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_13_LC_2_20_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_2_20_6 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(N__19330),
            .in2(N__19414),
            .in3(N__19005),
            .lcout(throttle_command_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36097),
            .ce(N__19284),
            .sr(N__19249));
    defparam \pid_alt.source_pid_1_esr_12_LC_2_20_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_2_20_7 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_2_20_7  (
            .in0(N__19197),
            .in1(N__19402),
            .in2(N__19010),
            .in3(N__19335),
            .lcout(throttle_command_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36097),
            .ce(N__19284),
            .sr(N__19249));
    defparam \pid_alt.source_pid_1_esr_1_LC_2_21_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_1_LC_2_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_1_LC_2_21_2 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_1_LC_2_21_2  (
            .in0(N__19331),
            .in1(N__19448),
            .in2(N__19425),
            .in3(N__21104),
            .lcout(throttle_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36090),
            .ce(N__19285),
            .sr(N__19256));
    defparam \pid_alt.source_pid_1_esr_4_LC_2_21_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_2_21_4 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_2_21_4  (
            .in0(N__19332),
            .in1(N__18952),
            .in2(N__15998),
            .in3(N__19490),
            .lcout(throttle_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36090),
            .ce(N__19285),
            .sr(N__19256));
    defparam \pid_alt.source_pid_1_esr_5_LC_2_21_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_2_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_2_21_5 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_2_21_5  (
            .in0(N__18953),
            .in1(N__19419),
            .in2(N__19223),
            .in3(N__19334),
            .lcout(throttle_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36090),
            .ce(N__19285),
            .sr(N__19256));
    defparam \pid_alt.source_pid_1_esr_0_LC_2_21_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_0_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_0_LC_2_21_7 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_0_LC_2_21_7  (
            .in0(N__19447),
            .in1(N__19415),
            .in2(N__18680),
            .in3(N__19333),
            .lcout(throttle_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36090),
            .ce(N__19285),
            .sr(N__19256));
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_2_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_2_22_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIG4JI2_11_LC_2_22_0  (
            .in0(N__16074),
            .in1(N__21475),
            .in2(N__22358),
            .in3(N__22263),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_2_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_2_22_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIALRT5_11_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(N__22628),
            .in2(N__16148),
            .in3(N__16145),
            .lcout(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_2_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_2_22_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI03DH2_11_LC_2_22_2  (
            .in0(N__16122),
            .in1(N__16134),
            .in2(N__22123),
            .in3(N__22001),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_2_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_2_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_2_22_3  (
            .in0(N__29490),
            .in1(N__16075),
            .in2(_gnd_net_),
            .in3(N__16123),
            .lcout(),
            .ltout(\ppm_encoder_1.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_2_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_2_22_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_2_22_4  (
            .in0(_gnd_net_),
            .in1(N__29268),
            .in2(N__16139),
            .in3(N__16135),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_2_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_2_22_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_2_22_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_2_22_5  (
            .in0(N__16136),
            .in1(N__24970),
            .in2(N__21260),
            .in3(N__19070),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36082),
            .ce(),
            .sr(N__36751));
    defparam \ppm_encoder_1.elevator_11_LC_2_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_2_22_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_2_22_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_2_22_6  (
            .in0(N__16124),
            .in1(N__29738),
            .in2(N__24997),
            .in3(N__24440),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36082),
            .ce(),
            .sr(N__36751));
    defparam \ppm_encoder_1.throttle_11_LC_2_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_2_22_7 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_2_22_7  (
            .in0(N__16112),
            .in1(N__16076),
            .in2(N__16085),
            .in3(N__24971),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36082),
            .ce(),
            .sr(N__36751));
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0  (
            .in0(N__16158),
            .in1(N__22314),
            .in2(N__21445),
            .in3(N__22261),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__19712),
            .in2(N__16232),
            .in3(N__16229),
            .lcout(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2  (
            .in0(N__16206),
            .in1(N__16218),
            .in2(N__22106),
            .in3(N__21999),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3  (
            .in0(N__29462),
            .in1(N__16159),
            .in2(_gnd_net_),
            .in3(N__16207),
            .lcout(),
            .ltout(\ppm_encoder_1.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_2_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_2_23_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_2_23_4  (
            .in0(N__29262),
            .in1(_gnd_net_),
            .in2(N__16223),
            .in3(N__16219),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_2_23_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_2_23_5  (
            .in0(N__16220),
            .in1(N__18908),
            .in2(N__24998),
            .in3(N__20978),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36073),
            .ce(),
            .sr(N__36754));
    defparam \ppm_encoder_1.elevator_7_LC_2_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_2_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_2_23_6 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_2_23_6  (
            .in0(N__16208),
            .in1(N__24080),
            .in2(N__28988),
            .in3(N__24980),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36073),
            .ce(),
            .sr(N__36754));
    defparam \ppm_encoder_1.throttle_7_LC_2_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_2_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_2_23_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_2_23_7  (
            .in0(N__16196),
            .in1(N__16183),
            .in2(N__24999),
            .in3(N__16160),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36073),
            .ce(),
            .sr(N__36754));
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_2_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_2_24_0 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \ppm_encoder_1.elevator_RNI47DH2_13_LC_2_24_0  (
            .in0(N__21998),
            .in1(N__24335),
            .in2(N__29534),
            .in3(N__22082),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_2_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_2_24_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIKVRT5_13_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__16607),
            .in2(N__16304),
            .in3(N__16292),
            .lcout(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_2_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_2_24_2 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \ppm_encoder_1.elevator_RNI8GVN2_6_LC_2_24_2  (
            .in0(N__21996),
            .in1(N__29302),
            .in2(N__29123),
            .in3(N__22078),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_2_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_2_24_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIO1KK2_6_LC_2_24_3  (
            .in0(N__29325),
            .in1(N__24607),
            .in2(N__22342),
            .in3(N__22224),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_2_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_2_24_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEDI96_6_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__19862),
            .in2(N__16301),
            .in3(N__16298),
            .lcout(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_2_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_2_24_5 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIK8JI2_13_LC_2_24_5  (
            .in0(N__23693),
            .in1(N__24560),
            .in2(N__22341),
            .in3(N__22223),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_2_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_2_24_7 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_2_24_7  (
            .in0(N__16285),
            .in1(N__16273),
            .in2(N__22105),
            .in3(N__21997),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_2_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_2_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIVO123_0_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__16256),
            .in2(N__19837),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_2_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_2_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(N__19126),
            .in2(N__19100),
            .in3(N__16238),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_2_25_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_2_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_2_25_2  (
            .in0(_gnd_net_),
            .in1(N__19562),
            .in2(N__19502),
            .in3(N__16235),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_2_25_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_2_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_2_25_3  (
            .in0(_gnd_net_),
            .in1(N__19652),
            .in2(N__19640),
            .in3(N__16439),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_2_25_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_2_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_2_25_4  (
            .in0(_gnd_net_),
            .in1(N__19526),
            .in2(N__20168),
            .in3(N__16436),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_2_25_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_2_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_2_25_5  (
            .in0(_gnd_net_),
            .in1(N__16433),
            .in2(N__16412),
            .in3(N__16403),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_2_25_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_2_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_2_25_6  (
            .in0(_gnd_net_),
            .in1(N__19861),
            .in2(N__16400),
            .in3(N__16391),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_2_25_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_2_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_2_25_7  (
            .in0(_gnd_net_),
            .in1(N__19708),
            .in2(N__16388),
            .in3(N__16376),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_2_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_2_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_2_26_0  (
            .in0(_gnd_net_),
            .in1(N__22159),
            .in2(N__22145),
            .in3(N__16373),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_2_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_2_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_2_26_1  (
            .in0(_gnd_net_),
            .in1(N__19576),
            .in2(N__16370),
            .in3(N__16352),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_2_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_2_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_2_26_2  (
            .in0(_gnd_net_),
            .in1(N__19609),
            .in2(N__16349),
            .in3(N__16331),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_2_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_2_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_2_26_3  (
            .in0(_gnd_net_),
            .in1(N__22627),
            .in2(N__16328),
            .in3(N__16625),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_2_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_2_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_2_26_4  (
            .in0(_gnd_net_),
            .in1(N__21781),
            .in2(N__21767),
            .in3(N__16610),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_2_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_2_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_2_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_2_26_5  (
            .in0(_gnd_net_),
            .in1(N__16603),
            .in2(N__16586),
            .in3(N__16562),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_2_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_2_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_2_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_2_26_6  (
            .in0(_gnd_net_),
            .in1(N__16559),
            .in2(N__16553),
            .in3(N__16520),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_2_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_2_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(N__16517),
            .in2(N__16505),
            .in3(N__16478),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_2_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_2_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_2_27_0  (
            .in0(_gnd_net_),
            .in1(N__16664),
            .in2(_gnd_net_),
            .in3(N__16475),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_2_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_2_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_2_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_2_27_1  (
            .in0(_gnd_net_),
            .in1(N__16445),
            .in2(_gnd_net_),
            .in3(N__16463),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_2_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_2_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_2_27_2  (
            .in0(_gnd_net_),
            .in1(N__16670),
            .in2(_gnd_net_),
            .in3(N__16460),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_2_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_2_27_3 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_2_27_3  (
            .in0(N__30342),
            .in1(_gnd_net_),
            .in2(N__30097),
            .in3(N__22985),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_2_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_2_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_2_27_4 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_2_27_4  (
            .in0(N__19922),
            .in1(N__30304),
            .in2(N__23045),
            .in3(N__30072),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_2_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_2_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_2_27_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_2_27_5  (
            .in0(N__30394),
            .in1(_gnd_net_),
            .in2(N__30096),
            .in3(N__22983),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_27_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_27_6  (
            .in0(N__22984),
            .in1(N__30065),
            .in2(_gnd_net_),
            .in3(N__30343),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_7  (
            .in0(N__23292),
            .in1(N__24374),
            .in2(N__30098),
            .in3(N__19921),
            .lcout(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_2_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_2_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_2_28_0  (
            .in0(_gnd_net_),
            .in1(N__16658),
            .in2(N__22655),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_28_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_2_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_2_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_2_28_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_2_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16652),
            .in3(N__16637),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_2_28_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_2_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_2_28_2  (
            .in0(_gnd_net_),
            .in1(N__19631),
            .in2(N__19973),
            .in3(N__16634),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_2_28_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_2_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_2_28_3  (
            .in0(_gnd_net_),
            .in1(N__19742),
            .in2(_gnd_net_),
            .in3(N__16631),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_2_28_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_2_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_2_28_4  (
            .in0(_gnd_net_),
            .in1(N__20144),
            .in2(_gnd_net_),
            .in3(N__16628),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_2_28_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_2_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_2_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_2_28_5  (
            .in0(_gnd_net_),
            .in1(N__16760),
            .in2(_gnd_net_),
            .in3(N__16748),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_2_28_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_2_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_2_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_2_28_6  (
            .in0(_gnd_net_),
            .in1(N__16745),
            .in2(N__19892),
            .in3(N__16739),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_2_28_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_2_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_2_28_7  (
            .in0(_gnd_net_),
            .in1(N__19718),
            .in2(_gnd_net_),
            .in3(N__16736),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_2_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_2_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_2_29_0  (
            .in0(_gnd_net_),
            .in1(N__16733),
            .in2(_gnd_net_),
            .in3(N__16724),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_2_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_2_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_2_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_2_29_1  (
            .in0(_gnd_net_),
            .in1(N__16721),
            .in2(_gnd_net_),
            .in3(N__16700),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_2_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_2_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_2_29_2  (
            .in0(_gnd_net_),
            .in1(N__19541),
            .in2(_gnd_net_),
            .in3(N__16691),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_2_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_2_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_2_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_2_29_3  (
            .in0(_gnd_net_),
            .in1(N__23306),
            .in2(_gnd_net_),
            .in3(N__16682),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_2_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_2_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_2_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_2_29_4  (
            .in0(_gnd_net_),
            .in1(N__19979),
            .in2(_gnd_net_),
            .in3(N__16673),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_2_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_2_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__16856),
            .in2(N__16850),
            .in3(N__16835),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_2_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_2_29_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_2_29_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19991),
            .in3(N__16826),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_2_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_2_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_2_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_2_29_7  (
            .in0(_gnd_net_),
            .in1(N__16823),
            .in2(_gnd_net_),
            .in3(N__16808),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_2_30_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_2_30_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_2_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_2_30_0  (
            .in0(_gnd_net_),
            .in1(N__22871),
            .in2(_gnd_net_),
            .in3(N__16805),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_2_30_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_2_30_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_2_30_1  (
            .in0(_gnd_net_),
            .in1(N__16802),
            .in2(_gnd_net_),
            .in3(N__16784),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_2_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_2_30_2 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_2_30_2  (
            .in0(N__30294),
            .in1(N__23088),
            .in2(N__30100),
            .in3(N__16781),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_2_30_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_2_30_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_2_30_5 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_2_30_5  (
            .in0(N__30076),
            .in1(N__29388),
            .in2(N__29279),
            .in3(N__36912),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36017),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_3_5_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_3_5_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_3_5_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_3_5_0  (
            .in0(_gnd_net_),
            .in1(N__31222),
            .in2(_gnd_net_),
            .in3(N__21637),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36162),
            .ce(N__25757),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_5_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_5_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_5_1  (
            .in0(N__21638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31373),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36162),
            .ce(N__25757),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_5_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_5_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_5_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_5_6  (
            .in0(_gnd_net_),
            .in1(N__30749),
            .in2(_gnd_net_),
            .in3(N__21635),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36162),
            .ce(N__25757),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_5_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_5_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_5_7  (
            .in0(N__21636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31841),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36162),
            .ce(N__25757),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_6_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_6_2  (
            .in0(_gnd_net_),
            .in1(N__31499),
            .in2(_gnd_net_),
            .in3(N__21632),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36159),
            .ce(N__25754),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_3_9_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_3_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26183),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36149),
            .ce(N__25652),
            .sr(N__36693));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_10_0 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_3_10_0  (
            .in0(N__30846),
            .in1(N__25843),
            .in2(N__16874),
            .in3(N__16924),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36145),
            .ce(),
            .sr(N__36695));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_10_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_3_10_1  (
            .in0(N__25844),
            .in1(N__16866),
            .in2(N__31221),
            .in3(N__16906),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36145),
            .ce(),
            .sr(N__36695));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_10_2 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_3_10_2  (
            .in0(N__31840),
            .in1(N__25842),
            .in2(N__16873),
            .in3(N__16891),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36145),
            .ce(),
            .sr(N__36695));
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3  (
            .in0(N__31210),
            .in1(N__30845),
            .in2(_gnd_net_),
            .in3(N__31839),
            .lcout(),
            .ltout(\Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_10_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_3_10_4  (
            .in0(N__31360),
            .in1(N__31654),
            .in2(N__16877),
            .in3(N__28070),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_10_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_3_10_5  (
            .in0(N__25841),
            .in1(N__31498),
            .in2(N__17054),
            .in3(N__17050),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36145),
            .ce(),
            .sr(N__36695));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_3_11_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_3_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17027),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_3_11_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_3_11_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_3_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26179),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36141),
            .ce(N__25709),
            .sr(N__36701));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_3_11_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_3_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20657),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_3_11_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_3_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20669),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_3_11_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_3_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20663),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20675),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_1_LC_3_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_3_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16988),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_3_11_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_3_11_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_3_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_3_11_7  (
            .in0(N__26090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36141),
            .ce(N__25709),
            .sr(N__36701));
    defparam \pid_alt.error_axb_12_LC_3_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_3_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17165),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_3_12_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_3_12_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_3_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25963),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36136),
            .ce(N__25648),
            .sr(N__36705));
    defparam \pid_alt.error_axb_13_LC_3_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_3_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17153),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_3_12_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_3_12_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_3_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26261),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36136),
            .ce(N__25648),
            .sr(N__36705));
    defparam \pid_alt.error_axb_14_LC_3_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_3_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20651),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_2_LC_3_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_3_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20645),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_3_LC_3_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_3_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_3_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20639),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_LC_3_13_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_LC_3_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__18271),
            .in2(N__18240),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_13_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__17126),
            .in2(N__17105),
            .in3(N__17057),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_13_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__17660),
            .in2(N__17636),
            .in3(N__17591),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_13_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(N__17588),
            .in2(N__17567),
            .in3(N__17522),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__17519),
            .in2(N__17498),
            .in3(N__17420),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__17417),
            .in2(N__17378),
            .in3(N__17306),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(N__20398),
            .in2(N__20435),
            .in3(N__17282),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__20223),
            .in2(N__20249),
            .in3(N__17255),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(N__36132),
            .ce(N__18294),
            .sr(N__36707));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_14_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__17252),
            .in2(N__17230),
            .in3(N__17174),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_14_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__18071),
            .in2(N__18049),
            .in3(N__17996),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_14_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__17993),
            .in2(N__17972),
            .in3(N__17918),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_14_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__17915),
            .in2(N__17894),
            .in3(N__17837),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_14_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__17834),
            .in2(N__17813),
            .in3(N__17750),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_14_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__17740),
            .in2(N__17720),
            .in3(N__17672),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(N__36127),
            .ce(N__18295),
            .sr(N__36711));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_LUT4_0_LC_3_14_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_LUT4_0_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_LUT4_0_LC_3_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_LUT4_0_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__18157),
            .in2(_gnd_net_),
            .in3(N__17669),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_LUT4_0_LC_3_14_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_LUT4_0_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_LUT4_0_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_LUT4_0_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18388),
            .in3(N__17666),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_LUT4_0_LC_3_15_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_LUT4_0_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_LUT4_0_LC_3_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_LUT4_0_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__18509),
            .in2(_gnd_net_),
            .in3(N__17663),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_LUT4_0_LC_3_15_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_LUT4_0_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_LUT4_0_LC_3_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_LUT4_0_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__18877),
            .in2(_gnd_net_),
            .in3(N__18335),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_LUT4_0_LC_3_15_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_LUT4_0_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_LUT4_0_LC_3_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_LUT4_0_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__20629),
            .in2(_gnd_net_),
            .in3(N__18332),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_LUT4_0_LC_3_15_3 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_LUT4_0_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_LUT4_0_LC_3_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_LUT4_0_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__18604),
            .in2(_gnd_net_),
            .in3(N__18329),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_LUT4_0_LC_3_15_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_LUT4_0_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_LUT4_0_LC_3_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_LUT4_0_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__20873),
            .in2(_gnd_net_),
            .in3(N__18326),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_3_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_3_15_5  (
            .in0(N__20874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18323),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36122),
            .ce(N__18296),
            .sr(N__36713));
    defparam \pid_alt.error_i_acumm_prereg_0_LC_3_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_0_LC_3_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_0_LC_3_16_0 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_0_LC_3_16_0  (
            .in0(N__18275),
            .in1(N__34163),
            .in2(N__18247),
            .in3(N__18195),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36117),
            .ce(),
            .sr(N__36718));
    defparam \pid_alt.error_i_acumm_prereg_20_LC_3_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_20_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_20_LC_3_16_1 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_20_LC_3_16_1  (
            .in0(N__34162),
            .in1(N__18176),
            .in2(N__20881),
            .in3(N__18427),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36117),
            .ce(),
            .sr(N__36718));
    defparam \pid_alt.error_i_acumm_prereg_14_LC_3_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_14_LC_3_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_14_LC_3_16_2 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_14_LC_3_16_2  (
            .in0(N__18167),
            .in1(N__34164),
            .in2(N__18158),
            .in3(N__18110),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36117),
            .ce(),
            .sr(N__36718));
    defparam \pid_alt.error_i_acumm_prereg_16_LC_3_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_16_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_16_LC_3_16_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_16_LC_3_16_3  (
            .in0(N__34161),
            .in1(N__18095),
            .in2(N__18089),
            .in3(N__18508),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36117),
            .ce(),
            .sr(N__36718));
    defparam \pid_alt.error_i_acumm_prereg_19_LC_3_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_19_LC_3_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_19_LC_3_16_4 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_19_LC_3_16_4  (
            .in0(N__18611),
            .in1(N__34165),
            .in2(N__18560),
            .in3(N__18566),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36117),
            .ce(),
            .sr(N__36718));
    defparam \pid_alt.error_p_reg_esr_RNIB03K_16_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIB03K_16_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIB03K_16_LC_3_16_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIB03K_16_LC_3_16_5  (
            .in0(N__18538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18507),
            .lcout(\pid_alt.error_p_reg_esr_RNIB03KZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_16_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_16_6  (
            .in0(N__29494),
            .in1(N__29275),
            .in2(_gnd_net_),
            .in3(N__22421),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_3_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_3_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_3_16_7  (
            .in0(N__29274),
            .in1(N__18446),
            .in2(_gnd_net_),
            .in3(N__19051),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_3_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_3_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_3_17_0  (
            .in0(N__26003),
            .in1(N__25962),
            .in2(N__26230),
            .in3(N__26082),
            .lcout(\dron_frame_decoder_1.N_194_4 ),
            .ltout(\dron_frame_decoder_1.N_194_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_3_17_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_3_17_1  (
            .in0(N__24028),
            .in1(_gnd_net_),
            .in2(N__18431),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_RNI58SG_15_LC_3_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_RNI58SG_15_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_RNI58SG_15_LC_3_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_RNI58SG_15_LC_3_17_3  (
            .in0(N__18817),
            .in1(N__18835),
            .in2(N__18428),
            .in3(N__18343),
            .lcout(\pid_alt.m7_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_15_LC_3_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_15_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_15_LC_3_17_4 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_15_LC_3_17_4  (
            .in0(N__18344),
            .in1(N__18404),
            .in2(N__18395),
            .in3(N__34160),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36111),
            .ce(),
            .sr(N__36723));
    defparam \pid_alt.error_i_acumm_prereg_17_LC_3_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_17_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_17_LC_3_17_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_17_LC_3_17_5  (
            .in0(N__34158),
            .in1(N__18890),
            .in2(N__18881),
            .in3(N__18836),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36111),
            .ce(),
            .sr(N__36723));
    defparam \pid_alt.error_i_acumm_prereg_18_LC_3_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_18_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_18_LC_3_17_6 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_18_LC_3_17_6  (
            .in0(N__18827),
            .in1(N__34159),
            .in2(N__20633),
            .in3(N__18818),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36111),
            .ce(),
            .sr(N__36723));
    defparam \pid_alt.pid_prereg_esr_RNIC62V1_12_LC_3_18_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIC62V1_12_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIC62V1_12_LC_3_18_1 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIC62V1_12_LC_3_18_1  (
            .in0(N__18994),
            .in1(N__19188),
            .in2(N__19413),
            .in3(N__19336),
            .lcout(\pid_alt.source_pid_9_0_tz_6 ),
            .ltout(\pid_alt.source_pid_9_0_tz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_8_LC_3_18_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_3_18_2 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \pid_alt.source_pid_1_8_LC_3_18_2  (
            .in0(N__21909),
            .in1(N__18775),
            .in2(N__18782),
            .in3(N__23886),
            .lcout(throttle_command_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36105),
            .ce(),
            .sr(N__19261));
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_3_18_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_3_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_3_18_4  (
            .in0(N__18753),
            .in1(N__18774),
            .in2(N__18705),
            .in3(N__18729),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_3_19_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI8H141_10_LC_3_19_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI8H141_10_LC_3_19_2  (
            .in0(N__18779),
            .in1(N__18754),
            .in2(N__18736),
            .in3(N__18654),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_3_19_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_3_19_3 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__18636),
            .in2(N__18713),
            .in3(N__18706),
            .lcout(\pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHBUI1_0_LC_3_19_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHBUI1_0_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHBUI1_0_LC_3_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHBUI1_0_LC_3_19_4  (
            .in0(N__21096),
            .in1(N__19360),
            .in2(N__19030),
            .in3(N__18676),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_3_19_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_3_19_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_3_19_5  (
            .in0(N__18655),
            .in1(N__18637),
            .in2(N__18623),
            .in3(N__23868),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI845S4_4_LC_3_19_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI845S4_4_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI845S4_4_LC_3_19_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI845S4_4_LC_3_19_6  (
            .in0(N__19481),
            .in1(N__18938),
            .in2(N__18941),
            .in3(N__19164),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_3_20_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_3_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_3_20_1  (
            .in0(N__19000),
            .in1(N__23869),
            .in2(N__19169),
            .in3(N__19480),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIJ1OF6_4_LC_3_20_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIJ1OF6_4_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIJ1OF6_4_LC_3_20_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIJ1OF6_4_LC_3_20_2  (
            .in0(N__19322),
            .in1(N__18937),
            .in2(N__18926),
            .in3(N__18964),
            .lcout(),
            .ltout(\pid_alt.N_92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIM9UC7_22_LC_3_20_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIM9UC7_22_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIM9UC7_22_LC_3_20_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIM9UC7_22_LC_3_20_3  (
            .in0(N__19394),
            .in1(N__23870),
            .in2(N__18923),
            .in3(N__35081),
            .lcout(),
            .ltout(\pid_alt.un1_reset_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI9BMSD_13_LC_3_20_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI9BMSD_13_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI9BMSD_13_LC_3_20_4 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI9BMSD_13_LC_3_20_4  (
            .in0(N__19323),
            .in1(N__19001),
            .in2(N__18920),
            .in3(N__18917),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(\pid_alt.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIU0UAE_1_LC_3_20_5 .C_ON=1'b0;
    defparam \pid_alt.state_RNIU0UAE_1_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIU0UAE_1_LC_3_20_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIU0UAE_1_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18911),
            .in3(N__23871),
            .lcout(\pid_alt.N_60_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_3_21_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_3_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_c_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__24652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_3_21_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_3_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__20974),
            .in2(_gnd_net_),
            .in3(N__18896),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_3_21_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_3_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__21871),
            .in2(_gnd_net_),
            .in3(N__18893),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_3_21_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_3_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__20908),
            .in2(_gnd_net_),
            .in3(N__19076),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_3_21_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_3_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__24199),
            .in2(_gnd_net_),
            .in3(N__19073),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_3_21_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_3_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(N__21256),
            .in2(_gnd_net_),
            .in3(N__19064),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_3_21_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_3_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__21742),
            .in2(_gnd_net_),
            .in3(N__19061),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_3_21_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_3_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__24133),
            .in2(N__28602),
            .in3(N__19058),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_3_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_3_22_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_3_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_3_22_0  (
            .in0(_gnd_net_),
            .in1(N__21164),
            .in2(_gnd_net_),
            .in3(N__19055),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36074),
            .ce(N__27301),
            .sr(N__36744));
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_4_LC_3_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_4_LC_3_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23741),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36074),
            .ce(N__27301),
            .sr(N__36744));
    defparam \pid_alt.source_pid_1_esr_3_LC_3_23_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_3_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_3_LC_3_23_1 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_3_LC_3_23_1  (
            .in0(N__19441),
            .in1(N__19031),
            .in2(N__19430),
            .in3(N__19343),
            .lcout(throttle_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36063),
            .ce(N__19286),
            .sr(N__19262));
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_3_23_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_3_23_3 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG2382_12_LC_3_23_3  (
            .in0(N__19199),
            .in1(N__19009),
            .in2(_gnd_net_),
            .in3(N__18968),
            .lcout(\pid_alt.N_88 ),
            .ltout(\pid_alt.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_3_23_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_3_23_4 .LUT_INIT=16'b1111001011110010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_3_23_4  (
            .in0(N__19154),
            .in1(N__19489),
            .in2(N__19451),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_90 ),
            .ltout(\pid_alt.N_90_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_2_LC_3_23_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_2_LC_3_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_2_LC_3_23_5 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_2_LC_3_23_5  (
            .in0(N__19426),
            .in1(N__19364),
            .in2(N__19346),
            .in3(N__19342),
            .lcout(throttle_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36063),
            .ce(N__19286),
            .sr(N__19262));
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_3_23_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_3_23_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__19222),
            .in2(_gnd_net_),
            .in3(N__19198),
            .lcout(\pid_alt.N_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_3_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_3_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_3_23_7  (
            .in0(N__25267),
            .in1(N__22482),
            .in2(N__22406),
            .in3(N__30024),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_3_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_3_24_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_3_24_0  (
            .in0(N__22543),
            .in1(N__22527),
            .in2(N__30025),
            .in3(N__22407),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_3_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_3_24_1 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_3_24_1  (
            .in0(N__22002),
            .in1(N__22433),
            .in2(N__19133),
            .in3(N__29928),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_3_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_3_24_2 .LUT_INIT=16'b1010111100001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIALN65_1_LC_3_24_2  (
            .in0(N__25058),
            .in1(N__19130),
            .in2(N__19103),
            .in3(N__22222),
            .lcout(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_3  (
            .in0(N__19774),
            .in1(N__26677),
            .in2(N__22016),
            .in3(N__22095),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_3_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_3_24_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_3_24_4  (
            .in0(N__20164),
            .in1(_gnd_net_),
            .in2(N__19529),
            .in3(N__19514),
            .lcout(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_3_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_3_24_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_3_24_5  (
            .in0(N__22450),
            .in1(N__22576),
            .in2(N__22529),
            .in3(N__22542),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_3_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_3_24_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_3_24_6  (
            .in0(N__29927),
            .in1(_gnd_net_),
            .in2(N__19520),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_3_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_3_24_7 .LUT_INIT=16'b1011101100001011;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_3_24_7  (
            .in0(N__21844),
            .in1(N__22202),
            .in2(N__19517),
            .in3(N__26641),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_3_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_3_25_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_3_25_0  (
            .in0(N__22481),
            .in1(N__25266),
            .in2(N__22405),
            .in3(N__29879),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_3_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_3_25_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \ppm_encoder_1.throttle_RNIR7352_2_LC_3_25_1  (
            .in0(N__20533),
            .in1(N__22771),
            .in2(N__19508),
            .in3(N__19917),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_3_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_3_25_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5V123_2_LC_3_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19505),
            .in3(N__19552),
            .lcout(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_3_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_3_25_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_3_25_3  (
            .in0(N__29880),
            .in1(N__25185),
            .in2(_gnd_net_),
            .in3(N__22948),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_3_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_3_25_4 .LUT_INIT=16'b1001011010100101;
    LogicCell40 \ppm_encoder_1.throttle_RNIT9352_3_LC_3_25_4  (
            .in0(N__25186),
            .in1(N__24769),
            .in2(N__19935),
            .in3(N__22249),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_3_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_3_25_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI82223_3_LC_3_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19493),
            .in3(N__19651),
            .lcout(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_3_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_3_25_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_12_LC_3_25_6  (
            .in0(N__22950),
            .in1(N__27838),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_3_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_3_25_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_3_25_7  (
            .in0(N__29881),
            .in1(N__24258),
            .in2(_gnd_net_),
            .in3(N__22949),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_3_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_3_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__23253),
            .in2(_gnd_net_),
            .in3(N__29885),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_3_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_3_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__22575),
            .in2(_gnd_net_),
            .in3(N__25215),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_3_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_3_26_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19619),
            .in3(N__29883),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_3_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_3_26_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_3_26_3  (
            .in0(N__29888),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__22947),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_3_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_3_26_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_3_26_4  (
            .in0(N__22945),
            .in1(N__19598),
            .in2(_gnd_net_),
            .in3(N__29886),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_3_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_3_26_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIANUS_2_LC_3_26_5  (
            .in0(N__29884),
            .in1(N__20529),
            .in2(_gnd_net_),
            .in3(N__22944),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_3_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_3_26_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_3_26_6  (
            .in0(N__22946),
            .in1(_gnd_net_),
            .in2(N__25490),
            .in3(N__29887),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_26_7  (
            .in0(N__29253),
            .in1(N__21824),
            .in2(_gnd_net_),
            .in3(N__19775),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_3_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_3_27_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_3_27_0  (
            .in0(N__20124),
            .in1(N__19757),
            .in2(N__23228),
            .in3(N__19751),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36033),
            .ce(),
            .sr(N__36763));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_3_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_3_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_3_27_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_3_27_1  (
            .in0(N__25184),
            .in1(N__22978),
            .in2(_gnd_net_),
            .in3(N__29912),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_3_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_3_27_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_3_27_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_3_27_2  (
            .in0(N__20125),
            .in1(N__19736),
            .in2(N__23229),
            .in3(N__19730),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36033),
            .ce(),
            .sr(N__36763));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_3_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_3_27_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_3_27_3  (
            .in0(N__19693),
            .in1(N__22982),
            .in2(_gnd_net_),
            .in3(N__29914),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_3_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_3_27_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_3_27_4  (
            .in0(N__29913),
            .in1(_gnd_net_),
            .in2(N__23044),
            .in3(N__19692),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_3_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_3_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_3_27_5 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_3_27_5  (
            .in0(N__19694),
            .in1(N__27941),
            .in2(N__30579),
            .in3(N__21446),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_3_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_3_27_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_3_27_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_3_27_7  (
            .in0(N__23201),
            .in1(N__19682),
            .in2(N__19673),
            .in3(N__20126),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36033),
            .ce(),
            .sr(N__36763));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_3_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_3_28_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_3_28_1  (
            .in0(N__19938),
            .in1(N__23293),
            .in2(N__24386),
            .in3(N__30028),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_3_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_3_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_3_28_2  (
            .in0(N__23294),
            .in1(N__20528),
            .in2(N__30087),
            .in3(N__19936),
            .lcout(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_3_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_3_28_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_3_28_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_3_28_3  (
            .in0(N__23193),
            .in1(N__20122),
            .in2(N__19964),
            .in3(N__19952),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36023),
            .ce(),
            .sr(N__36767));
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_3_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_3_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_3_28_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_3_28_4  (
            .in0(N__23295),
            .in1(N__24622),
            .in2(N__30088),
            .in3(N__19937),
            .lcout(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_6_LC_3_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_3_28_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_3_28_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_3_28_5  (
            .in0(N__23194),
            .in1(N__20123),
            .in2(N__19883),
            .in3(N__19868),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36023),
            .ce(),
            .sr(N__36767));
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_3_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_3_28_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIERUS_6_LC_3_28_6  (
            .in0(N__30027),
            .in1(N__24621),
            .in2(_gnd_net_),
            .in3(N__23030),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_3_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_3_28_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_3_28_7  (
            .in0(N__23029),
            .in1(N__24381),
            .in2(_gnd_net_),
            .in3(N__30026),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_3_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_3_29_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_3_29_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_3_29_0  (
            .in0(N__23167),
            .in1(N__20105),
            .in2(N__19811),
            .in3(N__19799),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36018),
            .ce(),
            .sr(N__36770));
    defparam \ppm_encoder_1.init_pulses_4_LC_3_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_3_29_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_3_29_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_3_29_3  (
            .in0(N__20106),
            .in1(N__19793),
            .in2(N__23191),
            .in3(N__19787),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36018),
            .ce(),
            .sr(N__36770));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_3_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_3_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_3_29_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_4_LC_3_29_4  (
            .in0(N__20136),
            .in1(N__23076),
            .in2(_gnd_net_),
            .in3(N__30035),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_3_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_3_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_3_29_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_3_29_5  (
            .in0(N__30036),
            .in1(_gnd_net_),
            .in2(N__23090),
            .in3(N__20137),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_3_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_3_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_3_29_6 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_3_29_6  (
            .in0(N__20138),
            .in1(N__27924),
            .in2(N__30584),
            .in3(N__26648),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_3_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_3_29_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_3_29_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_3_29_7  (
            .in0(N__20107),
            .in1(N__20027),
            .in2(N__23192),
            .in3(N__20021),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36018),
            .ce(),
            .sr(N__36770));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_3_30_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_3_30_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_3_30_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_3_30_0  (
            .in0(N__30042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36877),
            .lcout(\ppm_encoder_1.N_1014_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_3_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_3_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_3_30_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_3_30_1  (
            .in0(N__23087),
            .in1(N__24301),
            .in2(_gnd_net_),
            .in3(N__30041),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_3_30_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_3_30_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_3_30_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_3_30_3  (
            .in0(N__25296),
            .in1(N__22504),
            .in2(N__27923),
            .in3(N__25238),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_3_30_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_3_30_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_3_30_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_3_30_4  (
            .in0(N__27894),
            .in1(N__23338),
            .in2(_gnd_net_),
            .in3(N__21476),
            .lcout(),
            .ltout(\ppm_encoder_1.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_3_30_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_3_30_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_3_30_5 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_3_30_5  (
            .in0(N__30607),
            .in1(_gnd_net_),
            .in2(N__19982),
            .in3(N__30569),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_3_30_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_3_30_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_3_30_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_3_30_6  (
            .in0(N__30040),
            .in1(_gnd_net_),
            .in2(N__27839),
            .in3(N__23086),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_3_30_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_3_30_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_3_30_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_3_30_7  (
            .in0(N__30608),
            .in1(N__27895),
            .in2(N__20537),
            .in3(N__30570),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_4_5_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_4_5_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__30989),
            .in2(_gnd_net_),
            .in3(N__21634),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36160),
            .ce(N__25755),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_4_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_4_9_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_4_9_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_4_9_0  (
            .in0(N__20485),
            .in1(N__33644),
            .in2(N__28187),
            .in3(N__31690),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36146),
            .ce(),
            .sr(N__36690));
    defparam \pid_alt.error_i_reg_esr_6_LC_4_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_4_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20471),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36142),
            .ce(N__20300),
            .sr(N__21570));
    defparam \pid_alt.error_p_reg_esr_RNI69J71_6_LC_4_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI69J71_6_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI69J71_6_LC_4_10_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI69J71_6_LC_4_10_3  (
            .in0(N__20459),
            .in1(N__20421),
            .in2(_gnd_net_),
            .in3(N__20399),
            .lcout(\pid_alt.error_p_reg_esr_RNI69J71Z0Z_6 ),
            .ltout(\pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIFL6F2_7_LC_4_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIFL6F2_7_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIFL6F2_7_LC_4_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIFL6F2_7_LC_4_10_4  (
            .in0(N__20263),
            .in1(N__20238),
            .in2(N__20342),
            .in3(N__20224),
            .lcout(\pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_7_LC_4_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_4_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36142),
            .ce(N__20300),
            .sr(N__21570));
    defparam \pid_alt.error_p_reg_esr_RNI9CJ71_7_LC_4_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI9CJ71_7_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI9CJ71_7_LC_4_10_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI9CJ71_7_LC_4_10_6  (
            .in0(N__20264),
            .in1(N__20239),
            .in2(_gnd_net_),
            .in3(N__20225),
            .lcout(\pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_4_11_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26009),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36137),
            .ce(N__25636),
            .sr(N__36696));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_4_11_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26089),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36137),
            .ce(N__25636),
            .sr(N__36696));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_4_11_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_4_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26051),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36137),
            .ce(N__25636),
            .sr(N__36696));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_4_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26126),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36137),
            .ce(N__25636),
            .sr(N__36696));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_11_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26231),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36137),
            .ce(N__25636),
            .sr(N__36696));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_4_12_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_4_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26046),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36133),
            .ce(N__25704),
            .sr(N__36702));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_4_12_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26260),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36133),
            .ce(N__25704),
            .sr(N__36702));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_4_12_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_4_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26005),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36133),
            .ce(N__25704),
            .sr(N__36702));
    defparam \pid_alt.error_p_reg_esr_RNIF43K_18_LC_4_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIF43K_18_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIF43K_18_LC_4_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIF43K_18_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__20622),
            .in2(_gnd_net_),
            .in3(N__20572),
            .lcout(\pid_alt.error_p_reg_esr_RNIF43KZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI1O4K_20_LC_4_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI1O4K_20_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI1O4K_20_LC_4_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI1O4K_20_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__20861),
            .in2(_gnd_net_),
            .in3(N__20803),
            .lcout(\pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_4_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31475),
            .lcout(frame_decoder_CH2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_4_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_4_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_4_14_1  (
            .in0(N__31835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_4_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30867),
            .lcout(frame_decoder_CH2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_4_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31199),
            .lcout(frame_decoder_CH2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_4_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_4_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31691),
            .lcout(frame_decoder_CH2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_4_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_4_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30737),
            .lcout(frame_decoder_CH2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_4_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_4_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_4_14_6  (
            .in0(N__31361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_4_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_4_14_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_4_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30988),
            .lcout(frame_decoder_CH2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36123),
            .ce(N__23555),
            .sr(N__36708));
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_4_15_2 .C_ON=1'b0;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_4_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_4_15_2  (
            .in0(N__23804),
            .in1(N__21042),
            .in2(_gnd_net_),
            .in3(N__23762),
            .lcout(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.N_881_i_l_ofx_LC_4_15_4 .C_ON=1'b0;
    defparam \scaler_2.N_881_i_l_ofx_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.N_881_i_l_ofx_LC_4_15_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \scaler_2.N_881_i_l_ofx_LC_4_15_4  (
            .in0(N__21071),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23651),
            .lcout(\scaler_2.N_881_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_4_15_5 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_4_15_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_4_15_5  (
            .in0(N__23650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21070),
            .lcout(\scaler_2.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_4_15_7 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_4_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__29087),
            .in2(_gnd_net_),
            .in3(N__29066),
            .lcout(\scaler_3.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_4_16_0 .C_ON=1'b1;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_4_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__21050),
            .in2(N__21043),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_6_LC_4_16_1 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_6_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_6_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_6_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__20992),
            .in2(N__21044),
            .in3(N__20999),
            .lcout(scaler_2_data_6),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_1 ),
            .carryout(\scaler_2.un2_source_data_0_cry_2 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_7_LC_4_16_2 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_7_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_7_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_7_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__20950),
            .in2(N__20996),
            .in3(N__20957),
            .lcout(scaler_2_data_7),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_2 ),
            .carryout(\scaler_2.un2_source_data_0_cry_3 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_8_LC_4_16_3 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_8_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_8_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_8_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__20929),
            .in2(N__20954),
            .in3(N__20936),
            .lcout(scaler_2_data_8),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_3 ),
            .carryout(\scaler_2.un2_source_data_0_cry_4 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_9_LC_4_16_4 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_9_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_9_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_9_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__21295),
            .in2(N__20933),
            .in3(N__20885),
            .lcout(scaler_2_data_9),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_4 ),
            .carryout(\scaler_2.un2_source_data_0_cry_5 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_10_LC_4_16_5 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_10_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_10_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_10_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__21274),
            .in2(N__21299),
            .in3(N__21281),
            .lcout(scaler_2_data_10),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_5 ),
            .carryout(\scaler_2.un2_source_data_0_cry_6 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_11_LC_4_16_6 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_11_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_11_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_11_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__21226),
            .in2(N__21278),
            .in3(N__21233),
            .lcout(scaler_2_data_11),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_6 ),
            .carryout(\scaler_2.un2_source_data_0_cry_7 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_12_LC_4_16_7 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_12_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_12_LC_4_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_12_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(N__21208),
            .in2(N__21230),
            .in3(N__21212),
            .lcout(scaler_2_data_12),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_7 ),
            .carryout(\scaler_2.un2_source_data_0_cry_8 ),
            .clk(N__36112),
            .ce(N__29573),
            .sr(N__36714));
    defparam \scaler_2.source_data_1_esr_13_LC_4_17_0 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_13_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_13_LC_4_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_13_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__21209),
            .in2(N__21185),
            .in3(N__21170),
            .lcout(scaler_2_data_13),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_9 ),
            .clk(N__36106),
            .ce(N__29571),
            .sr(N__36719));
    defparam \scaler_2.source_data_1_esr_14_LC_4_17_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_14_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_14_LC_4_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_2.source_data_1_esr_14_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21167),
            .lcout(scaler_2_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36106),
            .ce(N__29571),
            .sr(N__36719));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_4_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_4_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_4_18_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__30987),
            .in2(_gnd_net_),
            .in3(N__21624),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36098),
            .ce(N__28041),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_1_LC_4_19_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_1_LC_4_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_1_LC_4_19_1 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_alt.pid_prereg_1_LC_4_19_1  (
            .in0(N__34132),
            .in1(N__21137),
            .in2(N__21119),
            .in3(N__21097),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36091),
            .ce(),
            .sr(N__36727));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_4_19_2 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_4_19_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__34131),
            .in2(_gnd_net_),
            .in3(N__36895),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_1_LC_4_19_4 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_4_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34133),
            .lcout(\pid_alt.N_60_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36091),
            .ce(),
            .sr(N__36727));
    defparam \pid_alt.state_RNICP2N1_0_LC_4_19_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_4_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__23825),
            .in2(_gnd_net_),
            .in3(N__21623),
            .lcout(\pid_alt.N_422_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_4_20_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_4_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23885),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36083),
            .ce(N__21482),
            .sr(N__36730));
    defparam \ppm_encoder_1.elevator_13_LC_4_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_4_21_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_4_21_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_4_21_0  (
            .in0(N__24419),
            .in1(N__29657),
            .in2(N__24936),
            .in3(N__24328),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.rudder_11_LC_4_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_4_21_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_4_21_1 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_4_21_1  (
            .in0(N__26908),
            .in1(N__24858),
            .in2(N__25529),
            .in3(N__21468),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.rudder_7_LC_4_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_4_21_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_4_21_2  (
            .in0(N__25595),
            .in1(N__26566),
            .in2(N__24937),
            .in3(N__21432),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.throttle_10_LC_4_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_4_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_4_21_3 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_4_21_3  (
            .in0(N__21416),
            .in1(N__24859),
            .in2(N__21386),
            .in3(N__22599),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.throttle_13_LC_4_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_4_21_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_4_21_4 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_4_21_4  (
            .in0(N__21371),
            .in1(N__21350),
            .in2(N__24938),
            .in3(N__23689),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.throttle_2_LC_4_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_4_21_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_4_21_5 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_4_21_5  (
            .in0(N__21338),
            .in1(N__24860),
            .in2(N__21326),
            .in3(N__22764),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.throttle_4_LC_4_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_4_21_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_4_21_6  (
            .in0(N__21815),
            .in1(N__21800),
            .in2(N__24939),
            .in3(N__21843),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36075),
            .ce(),
            .sr(N__36736));
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_4_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_4_22_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNII6JI2_12_LC_4_22_0  (
            .in0(N__21648),
            .in1(N__27789),
            .in2(N__22359),
            .in3(N__22251),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_4_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_4_22_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIFQRT5_12_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__21788),
            .in2(N__21770),
            .in3(N__21752),
            .lcout(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_4_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_4_22_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI25DH2_12_LC_4_22_2  (
            .in0(N__21696),
            .in1(N__21708),
            .in2(N__22124),
            .in3(N__22006),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_4_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_4_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_4_22_3  (
            .in0(N__29489),
            .in1(N__21649),
            .in2(_gnd_net_),
            .in3(N__21697),
            .lcout(),
            .ltout(\ppm_encoder_1.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_4_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_4_22_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_4_22_4  (
            .in0(N__29223),
            .in1(_gnd_net_),
            .in2(N__21746),
            .in3(N__21709),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_4_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_4_22_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_4_22_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_4_22_5  (
            .in0(N__21710),
            .in1(N__24929),
            .in2(N__21743),
            .in3(N__21719),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36064),
            .ce(),
            .sr(N__36740));
    defparam \ppm_encoder_1.elevator_12_LC_4_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_4_22_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_4_22_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_4_22_6  (
            .in0(N__21698),
            .in1(N__29705),
            .in2(N__24983),
            .in3(N__24428),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36064),
            .ce(),
            .sr(N__36740));
    defparam \ppm_encoder_1.throttle_12_LC_4_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_4_22_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_4_22_7  (
            .in0(N__21686),
            .in1(N__21662),
            .in2(N__24984),
            .in3(N__21650),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36064),
            .ce(),
            .sr(N__36740));
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_4_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_4_23_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIS5KK2_8_LC_4_23_0  (
            .in0(N__24225),
            .in1(N__21882),
            .in2(N__22343),
            .in3(N__22250),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_4_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_4_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIONI96_8_LC_4_23_1  (
            .in0(N__22163),
            .in1(_gnd_net_),
            .in2(N__22148),
            .in3(N__21944),
            .lcout(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_4_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_4_23_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNICKVN2_8_LC_4_23_2  (
            .in0(N__21936),
            .in1(N__22791),
            .in2(N__22110),
            .in3(N__22000),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_4_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_4_23_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_4_23_3  (
            .in0(N__21883),
            .in1(N__29480),
            .in2(_gnd_net_),
            .in3(N__21937),
            .lcout(\ppm_encoder_1.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_8_LC_4_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_4_23_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_4_23_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_4_23_4  (
            .in0(N__21938),
            .in1(N__24476),
            .in2(N__24982),
            .in3(N__28943),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36056),
            .ce(),
            .sr(N__36745));
    defparam \ppm_encoder_1.throttle_8_LC_4_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_4_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_4_23_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_4_23_5  (
            .in0(N__21884),
            .in1(N__24921),
            .in2(N__21926),
            .in3(N__21893),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36056),
            .ce(),
            .sr(N__36745));
    defparam \ppm_encoder_1.aileron_8_LC_4_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_4_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_4_23_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_4_23_6  (
            .in0(N__21872),
            .in1(N__21854),
            .in2(N__24981),
            .in3(N__22792),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36056),
            .ce(),
            .sr(N__36745));
    defparam \ppm_encoder_1.rudder_8_LC_4_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_4_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_4_23_7 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_4_23_7  (
            .in0(N__25577),
            .in1(N__24226),
            .in2(N__26525),
            .in3(N__24928),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36056),
            .ce(),
            .sr(N__36745));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_4_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_4_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_4_24_0  (
            .in0(N__26678),
            .in1(N__21845),
            .in2(_gnd_net_),
            .in3(N__22483),
            .lcout(\ppm_encoder_1.N_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_4_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_4_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_4_24_1 .LUT_INIT=16'b1111000111111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_4_24_1  (
            .in0(N__23046),
            .in1(N__22544),
            .in2(N__36914),
            .in3(N__29967),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_4_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_4_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_4_24_2 .LUT_INIT=16'b1101110011011110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_4_24_2  (
            .in0(N__29963),
            .in1(N__36901),
            .in2(N__29252),
            .in3(N__23047),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_4_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_4_24_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_4_24_3 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_4_24_3  (
            .in0(N__36900),
            .in1(N__29218),
            .in2(N__22528),
            .in3(N__29966),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_4_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_4_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_4_24_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_4_24_4  (
            .in0(N__29962),
            .in1(N__22640),
            .in2(N__22451),
            .in3(N__36909),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_24_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_24_5  (
            .in0(N__22484),
            .in1(N__29217),
            .in2(N__36913),
            .in3(N__29965),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_24_6 .LUT_INIT=16'b1111111101000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_24_6  (
            .in0(N__29964),
            .in1(N__25279),
            .in2(N__23083),
            .in3(N__36902),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_4_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_4_24_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_4_24_7  (
            .in0(_gnd_net_),
            .in1(N__22574),
            .in2(_gnd_net_),
            .in3(N__22446),
            .lcout(\ppm_encoder_1.N_227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_4_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_4_25_0 .LUT_INIT=16'b0101010110000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_4_25_0  (
            .in0(N__27955),
            .in1(N__29482),
            .in2(N__29222),
            .in3(N__25225),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_4_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_4_25_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_4_25_1  (
            .in0(N__22432),
            .in1(N__22942),
            .in2(_gnd_net_),
            .in3(N__22401),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_4_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_4_25_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22658),
            .in3(N__29908),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_4_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_4_25_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_4_25_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_4_25_3  (
            .in0(N__29910),
            .in1(N__22639),
            .in2(N__25236),
            .in3(N__36911),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36042),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_4_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_4_25_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_4_25_4  (
            .in0(N__22943),
            .in1(N__23339),
            .in2(_gnd_net_),
            .in3(N__29909),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_4_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_4_25_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_4_25_5  (
            .in0(N__29481),
            .in1(N__22607),
            .in2(_gnd_net_),
            .in3(N__24107),
            .lcout(),
            .ltout(\ppm_encoder_1.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_4_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_4_25_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_4_25_6  (
            .in0(N__29181),
            .in1(_gnd_net_),
            .in2(N__22580),
            .in3(N__24164),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_4_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_4_25_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_4_25_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_4_25_7  (
            .in0(N__29911),
            .in1(N__35063),
            .in2(N__23384),
            .in3(N__22577),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36042),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_4_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_4_26_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_4_26_0  (
            .in0(N__27422),
            .in1(N__27451),
            .in2(N__27398),
            .in3(N__27481),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_4_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_4_26_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_4_26_1  (
            .in0(_gnd_net_),
            .in1(N__30437),
            .in2(_gnd_net_),
            .in3(N__27605),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_4_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_4_26_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_4_26_2  (
            .in0(N__22553),
            .in1(N__27635),
            .in2(N__22547),
            .in3(N__27371),
            .lcout(\ppm_encoder_1.N_145_17 ),
            .ltout(\ppm_encoder_1.N_145_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_4_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_4_26_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_4_26_3  (
            .in0(N__30176),
            .in1(N__24680),
            .in2(N__22727),
            .in3(N__25142),
            .lcout(\ppm_encoder_1.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_4_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_4_26_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_4_26_5  (
            .in0(N__30175),
            .in1(N__24746),
            .in2(N__22724),
            .in3(N__25141),
            .lcout(\ppm_encoder_1.N_238 ),
            .ltout(\ppm_encoder_1.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_4_26_6 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_4_26_6  (
            .in0(N__25334),
            .in1(N__25396),
            .in2(N__22715),
            .in3(N__24740),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36034),
            .ce(),
            .sr(N__36758));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_4_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_4_26_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_4_26_7  (
            .in0(_gnd_net_),
            .in1(N__24737),
            .in2(_gnd_net_),
            .in3(N__25333),
            .lcout(\ppm_encoder_1.PPM_STATE_59_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_27_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_27_0  (
            .in0(N__22694),
            .in1(N__27452),
            .in2(N__22667),
            .in3(N__27482),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_4_27_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_4_27_1  (
            .in0(N__22712),
            .in1(N__22700),
            .in2(_gnd_net_),
            .in3(N__27110),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_27_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_4_27_2 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_4_27_2  (
            .in0(N__22688),
            .in1(N__22679),
            .in2(N__27122),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_4_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_4_27_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_4_27_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_4_27_3  (
            .in0(N__24491),
            .in1(N__27111),
            .in2(_gnd_net_),
            .in3(N__24344),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_4_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_4_27_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_4_27_4  (
            .in0(N__27109),
            .in1(N__25100),
            .in2(_gnd_net_),
            .in3(N__23348),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_27_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_4_27_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_4_27_5  (
            .in0(N__22862),
            .in1(N__27112),
            .in2(_gnd_net_),
            .in3(N__25424),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_4_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_4_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_4_27_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_4_27_6  (
            .in0(N__22853),
            .in1(N__27694),
            .in2(N__22817),
            .in3(N__27661),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_27_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_4_27_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_4_27_7  (
            .in0(N__22847),
            .in1(N__27113),
            .in2(_gnd_net_),
            .in3(N__22829),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36024),
            .ce(N__27014),
            .sr(N__36760));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_4_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_4_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_4_28_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_4_28_0  (
            .in0(N__29260),
            .in1(N__22808),
            .in2(_gnd_net_),
            .in3(N__22796),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_4_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_4_28_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_4_28_1  (
            .in0(_gnd_net_),
            .in1(N__27107),
            .in2(N__22778),
            .in3(N__24212),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36019),
            .ce(N__26997),
            .sr(N__36764));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_28_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_28_2  (
            .in0(N__29259),
            .in1(N__29461),
            .in2(_gnd_net_),
            .in3(N__22775),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_4_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_4_28_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_4_28_3  (
            .in0(_gnd_net_),
            .in1(N__27106),
            .in2(N__22748),
            .in3(N__22745),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36019),
            .ce(N__26997),
            .sr(N__36764));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_4_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_4_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_4_28_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_4_28_4  (
            .in0(N__27105),
            .in1(N__23096),
            .in2(_gnd_net_),
            .in3(N__25163),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36019),
            .ce(N__26997),
            .sr(N__36764));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_4_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_4_28_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_4_28_5  (
            .in0(N__22733),
            .in1(N__27730),
            .in2(N__23393),
            .in3(N__27367),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_28_6  (
            .in0(N__29261),
            .in1(N__23441),
            .in2(_gnd_net_),
            .in3(N__23429),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_4_28_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_4_28_7  (
            .in0(_gnd_net_),
            .in1(N__27108),
            .in2(N__23408),
            .in3(N__23405),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36019),
            .ce(N__26997),
            .sr(N__36764));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_4_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_4_29_1 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_4_29_1  (
            .in0(N__23081),
            .in1(N__29273),
            .in2(N__29484),
            .in3(N__27897),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_4_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_4_29_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_4_29_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_4_29_2  (
            .in0(N__27898),
            .in1(N__35078),
            .in2(N__23369),
            .in3(N__30039),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36014),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_29_3 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_29_3  (
            .in0(N__30531),
            .in1(N__27896),
            .in2(N__30618),
            .in3(N__23366),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_4_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_4_29_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_4_29_4  (
            .in0(N__23337),
            .in1(N__23080),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_4_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_4_29_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_4_29_5  (
            .in0(N__30038),
            .in1(N__30112),
            .in2(_gnd_net_),
            .in3(N__23297),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_4_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_4_29_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_4_29_6  (
            .in0(N__29272),
            .in1(N__29460),
            .in2(_gnd_net_),
            .in3(N__24773),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_4_30_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_4_30_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_4_30_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_4_30_5  (
            .in0(N__30390),
            .in1(N__23082),
            .in2(_gnd_net_),
            .in3(N__30043),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_4_30_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_4_30_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_4_30_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_4_30_6  (
            .in0(N__25297),
            .in1(N__29392),
            .in2(_gnd_net_),
            .in3(N__25237),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_0_LC_5_9_2 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_5_9_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_5_9_2  (
            .in0(N__34129),
            .in1(N__23996),
            .in2(_gnd_net_),
            .in3(N__23956),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36143),
            .ce(),
            .sr(N__36689));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_10_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26229),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36138),
            .ce(N__25705),
            .sr(N__36691));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_10_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25964),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36138),
            .ce(N__25705),
            .sr(N__36691));
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_5_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_5_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_1_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__30969),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23501),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_11_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23486),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_11_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23471),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31696),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36128),
            .ce(N__25877),
            .sr(N__36697));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30738),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36128),
            .ce(N__25877),
            .sr(N__36697));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31362),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36128),
            .ce(N__25877),
            .sr(N__36697));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30983),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36128),
            .ce(N__25877),
            .sr(N__36697));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_13_3 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_5_13_3  (
            .in0(N__36889),
            .in1(N__28148),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_5_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_5_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__36888),
            .in2(_gnd_net_),
            .in3(N__28268),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_5_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_5_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_0_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31474),
            .lcout(frame_decoder_OFF2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_5_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_1_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31822),
            .lcout(frame_decoder_OFF2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_5_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_2_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30857),
            .lcout(frame_decoder_OFF2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_5_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_5_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_3_LC_5_14_3  (
            .in0(N__31209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_5_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_4_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31695),
            .lcout(frame_decoder_OFF2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_5_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_5_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30736),
            .lcout(frame_decoder_OFF2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_5_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_5_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_6_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31343),
            .lcout(frame_decoder_OFF2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_5_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_5_14_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_ess_7_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30982),
            .lcout(frame_decoder_OFF2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36118),
            .ce(N__23642),
            .sr(N__36706));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_5_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_5_15_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_5_15_0  (
            .in0(N__25911),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24063),
            .lcout(\dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_5_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_5_15_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_5_15_6  (
            .in0(N__25912),
            .in1(N__24064),
            .in2(N__24029),
            .in3(N__32421),
            .lcout(\dron_frame_decoder_1.state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_LC_5_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_5_16_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_5_16_0  (
            .in0(N__36942),
            .in1(N__33628),
            .in2(N__32813),
            .in3(N__31892),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36107),
            .ce(),
            .sr(N__36712));
    defparam \dron_frame_decoder_1.state_0_LC_5_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_5_16_5 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_5_16_5 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_5_16_5  (
            .in0(N__24065),
            .in1(N__32186),
            .in2(N__23627),
            .in3(N__23597),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36107),
            .ce(),
            .sr(N__36712));
    defparam \dron_frame_decoder_1.source_data_valid_LC_5_16_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_5_16_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_5_16_6  (
            .in0(N__25916),
            .in1(N__32422),
            .in2(_gnd_net_),
            .in3(N__23981),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36107),
            .ce(),
            .sr(N__36712));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_5_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_5_17_2 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_5_17_2  (
            .in0(N__23618),
            .in1(N__24040),
            .in2(N__23609),
            .in3(N__23704),
            .lcout(\dron_frame_decoder_1.state_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_5_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_5_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__25958),
            .in2(_gnd_net_),
            .in3(N__26081),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_5_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_5_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_5_17_4  (
            .in0(N__26225),
            .in1(N__24062),
            .in2(N__24044),
            .in3(N__26004),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_5_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_5_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_5_17_5  (
            .in0(N__26118),
            .in1(N__32416),
            .in2(N__26050),
            .in3(N__24002),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_5_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_5_17_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_5_17_6  (
            .in0(N__24024),
            .in1(N__24041),
            .in2(N__24032),
            .in3(N__32174),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36099),
            .ce(),
            .sr(N__36715));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_5_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_5_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__26178),
            .in2(_gnd_net_),
            .in3(N__26259),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_18_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_18_4 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_5_18_4  (
            .in0(N__23985),
            .in1(N__23867),
            .in2(N__34130),
            .in3(N__36875),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_4_LC_5_19_0 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_4_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_4_LC_5_19_0 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_2.source_data_1_4_LC_5_19_0  (
            .in0(N__36958),
            .in1(N__23819),
            .in2(N__23737),
            .in3(N__23779),
            .lcout(scaler_2_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36084),
            .ce(),
            .sr(N__36724));
    defparam \dron_frame_decoder_1.state_3_LC_5_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_5_19_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_5_19_2  (
            .in0(N__32161),
            .in1(N__23720),
            .in2(N__32206),
            .in3(N__23708),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36084),
            .ce(),
            .sr(N__36724));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_5_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_5_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_5_20_0  (
            .in0(N__29485),
            .in1(N__23688),
            .in2(_gnd_net_),
            .in3(N__24327),
            .lcout(\ppm_encoder_1.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_5_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_5_21_0 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_5_21_0  (
            .in0(N__27958),
            .in1(N__30568),
            .in2(N__24308),
            .in3(N__25777),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_5_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_5_21_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_5_21_1  (
            .in0(N__30567),
            .in1(N__24266),
            .in2(N__24236),
            .in3(N__27959),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_12_LC_5_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_5_21_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_5_21_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_5_21_4  (
            .in0(N__26869),
            .in1(N__25508),
            .in2(N__27799),
            .in3(N__24879),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36065),
            .ce(),
            .sr(N__36731));
    defparam \ppm_encoder_1.aileron_10_LC_5_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_5_21_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_5_21_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_5_21_5  (
            .in0(N__24200),
            .in1(N__24176),
            .in2(N__24940),
            .in3(N__24153),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36065),
            .ce(),
            .sr(N__36731));
    defparam \ppm_encoder_1.aileron_13_LC_5_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_5_21_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_5_21_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_5_21_6  (
            .in0(N__24137),
            .in1(N__24116),
            .in2(N__24942),
            .in3(N__29523),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36065),
            .ce(),
            .sr(N__36731));
    defparam \ppm_encoder_1.elevator_10_LC_5_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_5_21_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_5_21_7  (
            .in0(N__28868),
            .in1(N__24449),
            .in2(N__24941),
            .in3(N__24096),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36065),
            .ce(),
            .sr(N__36731));
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_5_22_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_5_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_c_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__29023),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_5_22_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_5_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(N__28978),
            .in2(_gnd_net_),
            .in3(N__24068),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_5_22_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_5_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(N__28939),
            .in2(_gnd_net_),
            .in3(N__24470),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_5_22_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_5_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__28903),
            .in2(_gnd_net_),
            .in3(N__24452),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_5_22_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_5_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(N__28864),
            .in2(_gnd_net_),
            .in3(N__24443),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_5_22_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_5_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(N__29737),
            .in2(_gnd_net_),
            .in3(N__24431),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_5_22_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_5_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(N__29704),
            .in2(_gnd_net_),
            .in3(N__24422),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_5_22_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_5_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_5_22_7  (
            .in0(_gnd_net_),
            .in1(N__29656),
            .in2(N__28674),
            .in3(N__24413),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_5_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_5_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_5_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__29627),
            .in2(_gnd_net_),
            .in3(N__24410),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36050),
            .ce(N__27267),
            .sr(N__36741));
    defparam \ppm_encoder_1.rudder_10_LC_5_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_5_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_5_24_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_5_24_1  (
            .in0(N__26431),
            .in1(N__25541),
            .in2(N__25455),
            .in3(N__24947),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36043),
            .ce(),
            .sr(N__36746));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_5_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_5_24_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_5_24_2  (
            .in0(N__30558),
            .in1(N__27948),
            .in2(_gnd_net_),
            .in3(N__24385),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_5_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_5_24_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_5_24_3  (
            .in0(_gnd_net_),
            .in1(N__24943),
            .in2(_gnd_net_),
            .in3(N__36890),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_5_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_5_24_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_5_24_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_5_24_4  (
            .in0(N__24944),
            .in1(N__24656),
            .in2(_gnd_net_),
            .in3(N__29112),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36043),
            .ce(),
            .sr(N__36746));
    defparam \ppm_encoder_1.elevator_6_LC_5_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_5_24_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_5_24_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_5_24_5  (
            .in0(N__29301),
            .in1(N__29027),
            .in2(_gnd_net_),
            .in3(N__24946),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36043),
            .ce(),
            .sr(N__36746));
    defparam \ppm_encoder_1.rudder_6_LC_5_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_5_24_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_5_24_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_5_24_6  (
            .in0(N__24945),
            .in1(N__24606),
            .in2(_gnd_net_),
            .in3(N__26608),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36043),
            .ce(),
            .sr(N__36746));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_5_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_5_24_7 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_5_24_7  (
            .in0(N__27949),
            .in1(N__24632),
            .in2(N__24608),
            .in3(N__30557),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_5_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_5_25_0 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_5_25_0  (
            .in0(N__27947),
            .in1(N__24587),
            .in2(N__24559),
            .in3(N__30545),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_13_LC_5_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_5_25_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_5_25_1 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_5_25_1  (
            .in0(N__24985),
            .in1(N__24555),
            .in2(N__26816),
            .in3(N__25802),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36035),
            .ce(),
            .sr(N__36752));
    defparam \ppm_encoder_1.throttle_0_LC_5_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_5_25_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_5_25_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_5_25_2  (
            .in0(N__24508),
            .in1(N__24987),
            .in2(_gnd_net_),
            .in3(N__24536),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36035),
            .ce(),
            .sr(N__36752));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_25_3 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_25_3  (
            .in0(N__29195),
            .in1(N__29466),
            .in2(_gnd_net_),
            .in3(N__24507),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_5_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_5_25_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_5_25_4  (
            .in0(N__29467),
            .in1(N__29196),
            .in2(_gnd_net_),
            .in3(N__25053),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_1_LC_5_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_5_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_5_25_5 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_5_25_5  (
            .in0(N__24986),
            .in1(N__25054),
            .in2(N__25091),
            .in3(N__25076),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36035),
            .ce(),
            .sr(N__36752));
    defparam \ppm_encoder_1.throttle_3_LC_5_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_5_25_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_5_25_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_5_25_7  (
            .in0(N__25034),
            .in1(N__25022),
            .in2(N__25000),
            .in3(N__24768),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36035),
            .ce(),
            .sr(N__36752));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_26_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_26_0  (
            .in0(N__27505),
            .in1(N__24738),
            .in2(N__27563),
            .in3(N__27531),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_5_26_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_5_26_1  (
            .in0(_gnd_net_),
            .in1(N__25358),
            .in2(_gnd_net_),
            .in3(N__25411),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36025),
            .ce(),
            .sr(N__36755));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_5_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_5_26_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_5_26_2  (
            .in0(N__25357),
            .in1(N__25395),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ppm_encoder_1.N_140_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_5_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_5_26_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_5_26_3 .LUT_INIT=16'b1100110011110100;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_5_26_3  (
            .in0(N__24739),
            .in1(N__24691),
            .in2(N__24719),
            .in3(N__24716),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36025),
            .ce(),
            .sr(N__36755));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_26_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_26_4  (
            .in0(N__27506),
            .in1(N__27562),
            .in2(N__25363),
            .in3(N__27532),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_26_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_26_5  (
            .in0(N__24674),
            .in1(N__24665),
            .in2(N__27533),
            .in3(N__27504),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_26_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_26_6  (
            .in0(N__27558),
            .in1(N__25157),
            .in2(N__25151),
            .in3(N__26944),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_5_26_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_5_26_7  (
            .in0(N__26945),
            .in1(N__27698),
            .in2(N__27668),
            .in3(N__27731),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_5_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_5_27_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_5_27_0  (
            .in0(_gnd_net_),
            .in1(N__25133),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_5_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_5_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_5_27_1  (
            .in0(_gnd_net_),
            .in1(N__28686),
            .in2(N__25127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_5_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_5_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_5_27_2  (
            .in0(_gnd_net_),
            .in1(N__25118),
            .in2(N__28700),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_5_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_5_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_5_27_3  (
            .in0(_gnd_net_),
            .in1(N__28678),
            .in2(N__27239),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_5_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_5_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_5_27_4  (
            .in0(_gnd_net_),
            .in1(N__25112),
            .in2(N__28701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_5_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_5_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(N__25106),
            .in2(N__28658),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_5_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_5_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_5_27_6  (
            .in0(_gnd_net_),
            .in1(N__27152),
            .in2(N__28702),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_5_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_5_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_5_27_7  (
            .in0(_gnd_net_),
            .in1(N__28685),
            .in2(N__30413),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_5_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_5_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_5_28_0  (
            .in0(_gnd_net_),
            .in1(N__25601),
            .in2(N__28672),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_28_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_5_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_5_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_5_28_1  (
            .in0(_gnd_net_),
            .in1(N__30263),
            .in2(N__28703),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_5_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_5_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_5_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25493),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_5_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_5_28_3 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_5_28_3  (
            .in0(N__27925),
            .in1(N__25489),
            .in2(N__25460),
            .in3(N__30533),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_28_4 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_28_4  (
            .in0(N__25412),
            .in1(N__25382),
            .in2(N__25364),
            .in3(N__35059),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_28_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_28_5  (
            .in0(N__29427),
            .in1(N__25292),
            .in2(_gnd_net_),
            .in3(N__25229),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_28_6 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_28_6  (
            .in0(N__30532),
            .in1(N__27926),
            .in2(N__30626),
            .in3(N__25190),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_28_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_28_7  (
            .in0(N__30236),
            .in1(N__30214),
            .in2(N__30329),
            .in3(N__30371),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_5_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_5_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_5_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_5_29_0  (
            .in0(_gnd_net_),
            .in1(N__26609),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_29_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_5_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_5_29_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_5_29_1  (
            .in0(_gnd_net_),
            .in1(N__26567),
            .in2(_gnd_net_),
            .in3(N__25580),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_5_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_5_29_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_5_29_2  (
            .in0(_gnd_net_),
            .in1(N__26524),
            .in2(_gnd_net_),
            .in3(N__25562),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_5_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_5_29_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_5_29_3  (
            .in0(_gnd_net_),
            .in1(N__26473),
            .in2(_gnd_net_),
            .in3(N__25544),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_5_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_5_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_5_29_4  (
            .in0(_gnd_net_),
            .in1(N__26432),
            .in2(_gnd_net_),
            .in3(N__25532),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_5_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_5_29_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_5_29_5  (
            .in0(_gnd_net_),
            .in1(N__26912),
            .in2(_gnd_net_),
            .in3(N__25511),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_5_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_5_29_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_5_29_6  (
            .in0(_gnd_net_),
            .in1(N__26870),
            .in2(_gnd_net_),
            .in3(N__25496),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_5_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_5_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_5_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_5_29_7  (
            .in0(_gnd_net_),
            .in1(N__26815),
            .in2(N__28673),
            .in3(N__25790),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_5_30_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_5_30_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_5_30_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_5_30_0  (
            .in0(_gnd_net_),
            .in1(N__26786),
            .in2(_gnd_net_),
            .in3(N__25787),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36010),
            .ce(N__27293),
            .sr(N__36768));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_8_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_7_8_6  (
            .in0(N__28177),
            .in1(N__33643),
            .in2(_gnd_net_),
            .in3(N__36887),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31223),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36129),
            .ce(N__28111),
            .sr(N__36692));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_7_11_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_7_11_0 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_5_LC_7_11_0  (
            .in0(N__28079),
            .in1(N__28240),
            .in2(N__25910),
            .in3(N__36882),
            .lcout(\dron_frame_decoder_1.N_390_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_4_LC_7_11_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_7_11_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_7_11_2  (
            .in0(N__32413),
            .in1(N__28241),
            .in2(N__28099),
            .in3(N__32187),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36124),
            .ce(),
            .sr(N__36694));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_11_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_11_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_11_3  (
            .in0(N__28239),
            .in1(N__25897),
            .in2(N__25618),
            .in3(N__28078),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_11_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_11_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25655),
            .in3(N__35075),
            .lcout(\dron_frame_decoder_1.N_382_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_7_LC_7_11_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_7_11_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_7_11_6  (
            .in0(N__32415),
            .in1(N__25617),
            .in2(N__28100),
            .in3(N__32189),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36124),
            .ce(),
            .sr(N__36694));
    defparam \dron_frame_decoder_1.state_6_LC_7_11_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_7_11_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_7_11_7  (
            .in0(N__32188),
            .in1(N__25901),
            .in2(N__25619),
            .in3(N__32414),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36124),
            .ce(),
            .sr(N__36694));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__25828),
            .in2(_gnd_net_),
            .in3(N__36891),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_2_LC_7_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_7_12_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_7_12_1  (
            .in0(N__25862),
            .in1(N__31106),
            .in2(N__25856),
            .in3(N__32881),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36119),
            .ce(),
            .sr(N__36698));
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_12_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_2_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__31449),
            .in2(_gnd_net_),
            .in3(N__30945),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_2_LC_7_12_3  (
            .in0(N__30852),
            .in1(N__31088),
            .in2(N__25865),
            .in3(N__30711),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__25852),
            .in2(_gnd_net_),
            .in3(N__33631),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_3_LC_7_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_7_12_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_3_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__25814),
            .in2(N__25817),
            .in3(N__32882),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36119),
            .ce(),
            .sr(N__36698));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_2  (
            .in0(N__25813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33563),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__28216),
            .in2(_gnd_net_),
            .in3(N__36884),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_7_14_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_7_14_0  (
            .in0(N__33561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28204),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_7_14_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_7_14_1  (
            .in0(N__36874),
            .in1(_gnd_net_),
            .in2(N__26144),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_7_14_4.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_7_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36873),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__28132),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_7_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31652),
            .lcout(frame_decoder_CH3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36100),
            .ce(N__28464),
            .sr(N__36709));
    defparam \uart_drone.data_esr_0_LC_7_16_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28321),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_1_LC_7_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28307),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_2_LC_7_16_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28291),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_3_LC_7_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28415),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_4_LC_7_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34226),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_5_LC_7_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_7_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28403),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_6_LC_7_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_7_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28390),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \uart_drone.data_esr_7_LC_7_16_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_7_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34409),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(N__31520),
            .sr(N__31562));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31491),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31827),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30844),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31697),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30716),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_7_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31358),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_17_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30959),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36085),
            .ce(N__28121),
            .sr(N__36716));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31494),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31828),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30856),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_7_18_3  (
            .in0(N__31202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31670),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_7_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_7_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30717),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31359),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_7_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_7_18_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_7_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30981),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36076),
            .ce(N__26291),
            .sr(N__36720));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_7_19_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_7_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__26696),
            .in2(N__26738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_7_19_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__26279),
            .in2(N__26273),
            .in3(N__26408),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_7_19_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__26405),
            .in2(N__26396),
            .in3(N__26387),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_7_19_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__26384),
            .in2(N__26378),
            .in3(N__26366),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_7_19_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__26363),
            .in2(N__26354),
            .in3(N__26345),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_7_19_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__26342),
            .in2(N__26336),
            .in3(N__26324),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_7_19_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__26321),
            .in2(N__26315),
            .in3(N__26303),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_7_19_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_7_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__28334),
            .in2(_gnd_net_),
            .in3(N__26300),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_7_20_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__26624),
            .in2(N__28671),
            .in3(N__26297),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_7_20_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_7_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26294),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_20_2 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_20_2  (
            .in0(N__26762),
            .in1(N__26739),
            .in2(_gnd_net_),
            .in3(N__26706),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_905_i_l_ofx_LC_7_20_6 .C_ON=1'b0;
    defparam \scaler_4.N_905_i_l_ofx_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_905_i_l_ofx_LC_7_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_905_i_l_ofx_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__28373),
            .in2(_gnd_net_),
            .in3(N__28354),
            .lcout(\scaler_4.N_905_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_21_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_7_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__26763),
            .in2(N__26618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_7_21_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__26578),
            .in2(N__26770),
            .in3(N__26585),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_7_LC_7_21_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__26536),
            .in2(N__26582),
            .in3(N__26543),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_8_LC_7_21_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__26488),
            .in2(N__26540),
            .in3(N__26495),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_9_LC_7_21_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__26443),
            .in2(N__26492),
            .in3(N__26450),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_10_LC_7_21_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__26923),
            .in2(N__26447),
            .in3(N__26411),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_11_LC_7_21_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__26881),
            .in2(N__26927),
            .in3(N__26888),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_12_LC_7_21_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_7_21_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__26839),
            .in2(N__26885),
            .in3(N__26846),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__36051),
            .ce(N__29570),
            .sr(N__36732));
    defparam \scaler_4.source_data_1_esr_13_LC_7_22_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__26843),
            .in2(N__26828),
            .in3(N__26792),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__36044),
            .ce(N__29569),
            .sr(N__36737));
    defparam \scaler_4.source_data_1_esr_14_LC_7_22_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_7_22_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_7_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26789),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36044),
            .ce(N__29569),
            .sr(N__36737));
    defparam \scaler_4.source_data_1_esr_5_LC_7_22_5 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_7_22_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_7_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_7_22_5  (
            .in0(N__26771),
            .in1(N__26740),
            .in2(_gnd_net_),
            .in3(N__26708),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36044),
            .ce(N__29569),
            .sr(N__36737));
    defparam \scaler_4.source_data_1_4_LC_7_23_6 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_7_23_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_7_23_6  (
            .in0(N__36977),
            .in1(N__26741),
            .in2(N__26663),
            .in3(N__26707),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36036),
            .ce(),
            .sr(N__36742));
    defparam \ppm_encoder_1.elevator_esr_4_LC_7_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_4_LC_7_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_4_LC_7_24_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_4_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(N__32027),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36026),
            .ce(N__27283),
            .sr(N__36747));
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26662),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36026),
            .ce(N__27283),
            .sr(N__36747));
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_24_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_7_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27335),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36026),
            .ce(N__27283),
            .sr(N__36747));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_7_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_7_25_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_7_25_0  (
            .in0(N__27390),
            .in1(N__27212),
            .in2(N__27179),
            .in3(N__27417),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_7_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_7_25_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_7_25_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_7_25_1  (
            .in0(N__27224),
            .in1(N__27121),
            .in2(_gnd_net_),
            .in3(N__29093),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36020),
            .ce(N__27013),
            .sr(N__36753));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_7_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_7_25_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_7_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_7_25_2  (
            .in0(N__27206),
            .in1(N__27118),
            .in2(_gnd_net_),
            .in3(N__27191),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36020),
            .ce(N__27013),
            .sr(N__36753));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_7_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_7_25_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_7_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_7_25_3  (
            .in0(N__27170),
            .in1(N__27120),
            .in2(_gnd_net_),
            .in3(N__30452),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36020),
            .ce(N__27013),
            .sr(N__36753));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_7_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_7_25_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_7_25_4  (
            .in0(N__27601),
            .in1(N__27158),
            .in2(N__27131),
            .in3(N__27631),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_7_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_7_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_7_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_7_25_5  (
            .in0(N__27117),
            .in1(N__29504),
            .in2(_gnd_net_),
            .in3(N__27140),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36020),
            .ce(N__27013),
            .sr(N__36753));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_7_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_7_25_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_7_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_7_25_6  (
            .in0(N__27119),
            .in1(N__27044),
            .in2(_gnd_net_),
            .in3(N__27026),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36020),
            .ce(N__27013),
            .sr(N__36753));
    defparam \ppm_encoder_1.counter_0_LC_7_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_7_26_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_7_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(N__26943),
            .in2(N__26969),
            .in3(N__26968),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_1_LC_7_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_7_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_7_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_7_26_1  (
            .in0(_gnd_net_),
            .in1(N__27557),
            .in2(_gnd_net_),
            .in3(N__27536),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_2_LC_7_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_7_26_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_7_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(N__27527),
            .in2(_gnd_net_),
            .in3(N__27509),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_3_LC_7_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_7_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_7_26_3  (
            .in0(_gnd_net_),
            .in1(N__27503),
            .in2(_gnd_net_),
            .in3(N__27485),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_4_LC_7_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_7_26_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_7_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__27477),
            .in2(_gnd_net_),
            .in3(N__27455),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_5_LC_7_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_7_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_7_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_7_26_5  (
            .in0(_gnd_net_),
            .in1(N__27447),
            .in2(_gnd_net_),
            .in3(N__27425),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_6_LC_7_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_7_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_7_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__27421),
            .in2(_gnd_net_),
            .in3(N__27401),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_7_LC_7_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_7_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_7_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_7_26_7  (
            .in0(_gnd_net_),
            .in1(N__27394),
            .in2(_gnd_net_),
            .in3(N__27374),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__36015),
            .ce(),
            .sr(N__27974));
    defparam \ppm_encoder_1.counter_8_LC_7_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_7_27_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_7_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(N__27360),
            .in2(_gnd_net_),
            .in3(N__27338),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_9_LC_7_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_7_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(N__27723),
            .in2(_gnd_net_),
            .in3(N__27701),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_10_LC_7_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_7_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__27693),
            .in2(_gnd_net_),
            .in3(N__27671),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_11_LC_7_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_7_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(N__27660),
            .in2(_gnd_net_),
            .in3(N__27638),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_12_LC_7_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_7_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_7_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__27630),
            .in2(_gnd_net_),
            .in3(N__27608),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_13_LC_7_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_7_27_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_7_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(N__27600),
            .in2(_gnd_net_),
            .in3(N__27578),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_14_LC_7_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_7_27_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_7_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(N__30433),
            .in2(_gnd_net_),
            .in3(N__27575),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_15_LC_7_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_7_27_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_7_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__30251),
            .in2(_gnd_net_),
            .in3(N__27572),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__36013),
            .ce(),
            .sr(N__27973));
    defparam \ppm_encoder_1.counter_16_LC_7_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_7_28_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_7_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__30213),
            .in2(_gnd_net_),
            .in3(N__27569),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__36011),
            .ce(),
            .sr(N__27972));
    defparam \ppm_encoder_1.counter_17_LC_7_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_7_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_7_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__30235),
            .in2(_gnd_net_),
            .in3(N__27566),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__36011),
            .ce(),
            .sr(N__27972));
    defparam \ppm_encoder_1.counter_18_LC_7_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_7_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_7_28_2  (
            .in0(_gnd_net_),
            .in1(N__30191),
            .in2(_gnd_net_),
            .in3(N__27977),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36011),
            .ce(),
            .sr(N__27972));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_29_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_29_2  (
            .in0(N__27922),
            .in1(N__27837),
            .in2(_gnd_net_),
            .in3(N__27803),
            .lcout(\ppm_encoder_1.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_8_2_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27773),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36156),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_8_2_3 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_8_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31022),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36156),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_8_2_5 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_8_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27767),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36156),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_4 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_4_4  (
            .in0(N__27761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36150),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_8_7_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27752),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36139),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_8_8_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27743),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36134),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_8_9_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27737),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36130),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__31988),
            .in2(_gnd_net_),
            .in3(N__33632),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state51_i_LC_8_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state51_i_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state51_i_LC_8_11_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.un1_state51_i_LC_8_11_1  (
            .in0(N__33633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36880),
            .lcout(\Commands_frame_decoder.un1_state51_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_8_11_2  (
            .in0(N__36881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_11_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__32356),
            .in2(_gnd_net_),
            .in3(N__28092),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_11_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_8_11_7  (
            .in0(N__30821),
            .in1(N__31079),
            .in2(N__31477),
            .in3(N__28066),
            .lcout(\Commands_frame_decoder.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_11_LC_8_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_8_12_0 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_8_12_0  (
            .in0(N__33624),
            .in1(N__27988),
            .in2(N__32300),
            .in3(N__32909),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36113),
            .ce(),
            .sr(N__36703));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2  (
            .in0(N__33623),
            .in1(N__27987),
            .in2(_gnd_net_),
            .in3(N__36879),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_10_LC_8_12_3  (
            .in0(N__27989),
            .in1(N__28004),
            .in2(_gnd_net_),
            .in3(N__32873),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36113),
            .ce(),
            .sr(N__36703));
    defparam \Commands_frame_decoder.state_7_LC_8_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_8_12_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_8_12_4  (
            .in0(N__32874),
            .in1(N__28176),
            .in2(N__33642),
            .in3(N__28277),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36113),
            .ce(),
            .sr(N__36703));
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIJN1J_7_LC_8_12_6  (
            .in0(N__33622),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28276),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_8_LC_8_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_8_12_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__28253),
            .in2(N__28256),
            .in3(N__32875),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36113),
            .ce(),
            .sr(N__36703));
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIKO1J_8_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__28252),
            .in2(_gnd_net_),
            .in3(N__33562),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_13_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__33955),
            .in2(_gnd_net_),
            .in3(N__35076),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_5_LC_8_14_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_8_14_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_8_14_1  (
            .in0(N__32406),
            .in1(N__28238),
            .in2(N__32120),
            .in3(N__32178),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36101),
            .ce(),
            .sr(N__36710));
    defparam \Commands_frame_decoder.state_5_LC_8_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_8_14_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_5_LC_8_14_2  (
            .in0(N__32868),
            .in1(N__28205),
            .in2(_gnd_net_),
            .in3(N__28217),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36101),
            .ce(),
            .sr(N__36710));
    defparam \uart_pc.data_rdy_LC_8_14_5 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_8_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__36324),
            .in2(_gnd_net_),
            .in3(N__33956),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36101),
            .ce(),
            .sr(N__36710));
    defparam \Commands_frame_decoder.state_6_LC_8_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_8_14_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_6_LC_8_14_6  (
            .in0(N__32869),
            .in1(N__28169),
            .in2(_gnd_net_),
            .in3(N__28193),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36101),
            .ce(),
            .sr(N__36710));
    defparam \Commands_frame_decoder.state_4_LC_8_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_8_14_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_4_LC_8_14_7  (
            .in0(N__28133),
            .in1(N__28147),
            .in2(_gnd_net_),
            .in3(N__32867),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36101),
            .ce(),
            .sr(N__36710));
    defparam \uart_pc.data_6_LC_8_15_1 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_8_15_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_6_LC_8_15_1  (
            .in0(N__31877),
            .in1(N__31725),
            .in2(N__31946),
            .in3(N__30921),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36093),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_15_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_15_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_8_15_2  (
            .in0(N__36314),
            .in1(N__35077),
            .in2(_gnd_net_),
            .in3(N__33953),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_8_15_3 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_8_15_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \uart_pc.data_1_4_LC_8_15_3  (
            .in0(N__31875),
            .in1(N__32696),
            .in2(N__28376),
            .in3(N__30682),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36093),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_8_15_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_8_15_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_8_15_4  (
            .in0(N__37255),
            .in1(N__32471),
            .in2(_gnd_net_),
            .in3(N__36885),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_5 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__28372),
            .in2(_gnd_net_),
            .in3(N__28355),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_8_15_7 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_8_15_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \uart_pc.data_2_LC_8_15_7  (
            .in0(N__31876),
            .in1(N__30853),
            .in2(N__32732),
            .in3(N__31724),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36093),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_8_16_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_0_LC_8_16_0  (
            .in0(N__31919),
            .in1(N__34362),
            .in2(N__28322),
            .in3(N__34264),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_8_16_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_1_LC_8_16_1  (
            .in0(N__34265),
            .in1(N__28306),
            .in2(N__34379),
            .in3(N__32768),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_8_16_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_8_16_2  (
            .in0(N__31586),
            .in1(N__34363),
            .in2(N__28295),
            .in3(N__34266),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \uart_drone.data_Aux_3_LC_8_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_8_16_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_3_LC_8_16_3  (
            .in0(N__34267),
            .in1(N__28414),
            .in2(N__34380),
            .in3(N__31568),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \uart_drone.data_Aux_5_LC_8_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_8_16_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_5_LC_8_16_5  (
            .in0(N__34268),
            .in1(N__28402),
            .in2(N__34381),
            .in3(N__31574),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \uart_drone.data_Aux_6_LC_8_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_8_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_8_16_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_8_16_6  (
            .in0(N__31580),
            .in1(N__34364),
            .in2(N__28391),
            .in3(N__34269),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36086),
            .ce(),
            .sr(N__34182));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_8_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_8_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31492),
            .lcout(frame_decoder_CH3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36077),
            .ce(N__28472),
            .sr(N__36721));
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_8_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_8_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_0_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31490),
            .lcout(frame_decoder_OFF3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_8_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_8_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_1_LC_8_18_1  (
            .in0(N__31802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_8_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_8_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_2_LC_8_18_2  (
            .in0(N__30834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_8_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_8_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_3_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31200),
            .lcout(frame_decoder_OFF3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_8_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_8_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_4_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31651),
            .lcout(frame_decoder_OFF3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_8_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_8_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_5_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30715),
            .lcout(frame_decoder_OFF3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_8_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_8_18_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_8_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_6_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31356),
            .lcout(frame_decoder_OFF3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_8_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_8_18_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_8_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_ess_7_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30957),
            .lcout(frame_decoder_OFF3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36066),
            .ce(N__31928),
            .sr(N__36725));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_8_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_8_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_8_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31201),
            .lcout(frame_decoder_CH3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_8_19_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_8_19_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_8_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_8_19_1  (
            .in0(N__31823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_8_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_8_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30828),
            .lcout(frame_decoder_CH3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_8_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_8_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_8_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30724),
            .lcout(frame_decoder_CH3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_8_19_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_8_19_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_8_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31357),
            .lcout(frame_decoder_CH3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_8_19_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_8_19_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_8_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30958),
            .lcout(frame_decoder_CH3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36057),
            .ce(N__28468),
            .sr(N__36728));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_8_20_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_8_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__32045),
            .in2(N__32090),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_8_20_1 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__28436),
            .in2(N__28430),
            .in3(N__28418),
            .lcout(\scaler_3.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_0 ),
            .carryout(\scaler_3.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_8_20_2 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__28847),
            .in2(N__28841),
            .in3(N__28829),
            .lcout(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_1 ),
            .carryout(\scaler_3.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_8_20_3 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__28826),
            .in2(N__28817),
            .in3(N__28808),
            .lcout(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_2 ),
            .carryout(\scaler_3.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_8_20_4 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__28805),
            .in2(N__28793),
            .in3(N__28781),
            .lcout(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_3 ),
            .carryout(\scaler_3.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_8_20_5 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__28778),
            .in2(N__28772),
            .in3(N__28760),
            .lcout(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_4 ),
            .carryout(\scaler_3.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_8_20_6 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_8_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__28757),
            .in2(N__28751),
            .in3(N__28739),
            .lcout(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_5 ),
            .carryout(\scaler_3.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_8_20_7 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_8_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(N__28736),
            .in2(_gnd_net_),
            .in3(N__28721),
            .lcout(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_6 ),
            .carryout(\scaler_3.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_8_21_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_8_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(N__29042),
            .in2(N__28657),
            .in3(N__28478),
            .lcout(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_8_21_1 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_8_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28475),
            .lcout(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.N_893_i_l_ofx_LC_8_21_2 .C_ON=1'b0;
    defparam \scaler_3.N_893_i_l_ofx_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.N_893_i_l_ofx_LC_8_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_3.N_893_i_l_ofx_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(N__29086),
            .in2(_gnd_net_),
            .in3(N__29062),
            .lcout(\scaler_3.N_893_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_8_21_7 .C_ON=1'b0;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_8_21_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_8_21_7  (
            .in0(N__29609),
            .in1(N__32091),
            .in2(_gnd_net_),
            .in3(N__32055),
            .lcout(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_8_22_0 .C_ON=1'b1;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_8_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__29610),
            .in2(N__29036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.source_data_1_esr_6_LC_8_22_1 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_6_LC_8_22_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_6_LC_8_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_6_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__28999),
            .in2(N__29617),
            .in3(N__29006),
            .lcout(scaler_3_data_6),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_1 ),
            .carryout(\scaler_3.un2_source_data_0_cry_2 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_7_LC_8_22_2 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_7_LC_8_22_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_7_LC_8_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_7_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__28954),
            .in2(N__29003),
            .in3(N__28961),
            .lcout(scaler_3_data_7),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_2 ),
            .carryout(\scaler_3.un2_source_data_0_cry_3 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_8_LC_8_22_3 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_8_LC_8_22_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_8_LC_8_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_8_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__28918),
            .in2(N__28958),
            .in3(N__28925),
            .lcout(scaler_3_data_8),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_3 ),
            .carryout(\scaler_3.un2_source_data_0_cry_4 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_9_LC_8_22_4 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_9_LC_8_22_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_9_LC_8_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_9_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__28879),
            .in2(N__28922),
            .in3(N__28886),
            .lcout(scaler_3_data_9),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_4 ),
            .carryout(\scaler_3.un2_source_data_0_cry_5 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_10_LC_8_22_5 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_10_LC_8_22_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_10_LC_8_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_10_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(N__29749),
            .in2(N__28883),
            .in3(N__28850),
            .lcout(scaler_3_data_10),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_5 ),
            .carryout(\scaler_3.un2_source_data_0_cry_6 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_11_LC_8_22_6 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_11_LC_8_22_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_11_LC_8_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_11_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(N__29716),
            .in2(N__29753),
            .in3(N__29723),
            .lcout(scaler_3_data_11),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_6 ),
            .carryout(\scaler_3.un2_source_data_0_cry_7 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_12_LC_8_22_7 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_12_LC_8_22_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_12_LC_8_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_12_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(N__29680),
            .in2(N__29720),
            .in3(N__29687),
            .lcout(scaler_3_data_12),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_7 ),
            .carryout(\scaler_3.un2_source_data_0_cry_8 ),
            .clk(N__36037),
            .ce(N__29568),
            .sr(N__36743));
    defparam \scaler_3.source_data_1_esr_13_LC_8_23_0 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_13_LC_8_23_0 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_13_LC_8_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_13_LC_8_23_0  (
            .in0(_gnd_net_),
            .in1(N__29684),
            .in2(N__29669),
            .in3(N__29633),
            .lcout(scaler_3_data_13),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_9 ),
            .clk(N__36027),
            .ce(N__29567),
            .sr(N__36748));
    defparam \scaler_3.source_data_1_esr_14_LC_8_23_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_14_LC_8_23_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_14_LC_8_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_3.source_data_1_esr_14_LC_8_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29630),
            .lcout(scaler_3_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36027),
            .ce(N__29567),
            .sr(N__36748));
    defparam \scaler_3.source_data_1_esr_5_LC_8_23_6 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_5_LC_8_23_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_5_LC_8_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.source_data_1_esr_5_LC_8_23_6  (
            .in0(N__29618),
            .in1(N__32092),
            .in2(_gnd_net_),
            .in3(N__32059),
            .lcout(scaler_3_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36027),
            .ce(N__29567),
            .sr(N__36748));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_8_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_8_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_8_24_0  (
            .in0(N__29244),
            .in1(N__29546),
            .in2(_gnd_net_),
            .in3(N__29533),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_8_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_8_24_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_8_24_5  (
            .in0(N__29498),
            .in1(N__29333),
            .in2(_gnd_net_),
            .in3(N__29303),
            .lcout(),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_8_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_8_24_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_8_24_6  (
            .in0(N__29245),
            .in1(_gnd_net_),
            .in2(N__29126),
            .in3(N__29122),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_8_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_8_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_8_25_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_8_25_5  (
            .in0(N__30625),
            .in1(N__30571),
            .in2(_gnd_net_),
            .in3(N__30464),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_27_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_27_0  (
            .in0(N__30446),
            .in1(N__30249),
            .in2(N__29768),
            .in3(N__30429),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_16_LC_8_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_8_27_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_8_27_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_8_27_2  (
            .in0(N__30401),
            .in1(N__30367),
            .in2(N__30139),
            .in3(N__30085),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36012),
            .ce(),
            .sr(N__36761));
    defparam \ppm_encoder_1.pulses2count_17_LC_8_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_8_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_8_27_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_8_27_4  (
            .in0(N__30353),
            .in1(N__30322),
            .in2(N__30140),
            .in3(N__30086),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36012),
            .ce(),
            .sr(N__36761));
    defparam \ppm_encoder_1.pulses2count_18_LC_8_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_8_27_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_8_27_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_8_27_5  (
            .in0(N__30084),
            .in1(N__30308),
            .in2(N__30275),
            .in3(N__30137),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36012),
            .ce(),
            .sr(N__36761));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_8_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_8_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_8_27_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_8_27_6  (
            .in0(N__30189),
            .in1(N__30271),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_8_27_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_8_27_7  (
            .in0(N__30250),
            .in1(N__30234),
            .in2(N__30215),
            .in3(N__30190),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_15_LC_8_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_8_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_8_28_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_8_28_3  (
            .in0(N__30161),
            .in1(N__29767),
            .in2(N__30138),
            .in3(N__30083),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36009),
            .ce(),
            .sr(N__36765));
    defparam \uart_pc_sync.aux_1__0__0_LC_9_2_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31007),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36153),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_2_3 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31016),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36153),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_rdy_LC_9_10_6 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_9_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__34335),
            .in2(_gnd_net_),
            .in3(N__31544),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36120),
            .ce(),
            .sr(N__36699));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_9_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_9_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_9_11_2  (
            .in0(N__30854),
            .in1(N__30973),
            .in2(N__31476),
            .in3(N__30729),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_9_11_3 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_9_11_3  (
            .in0(N__31055),
            .in1(N__31101),
            .in2(N__31001),
            .in3(N__30998),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_9_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_9_11_4 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_9_11_4 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \Commands_frame_decoder.state_0_LC_9_11_4  (
            .in0(N__32872),
            .in1(N__31083),
            .in2(N__30992),
            .in3(N__31031),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36114),
            .ce(),
            .sr(N__36704));
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_9_11_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_1_LC_9_11_5  (
            .in0(N__30974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31445),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_9_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_9_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_9_11_6  (
            .in0(N__30855),
            .in1(N__31046),
            .in2(N__30752),
            .in3(N__30730),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_LC_9_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_9_11_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_9_11_7  (
            .in0(N__31084),
            .in1(N__31102),
            .in2(N__30629),
            .in3(N__32871),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36114),
            .ce(),
            .sr(N__36704));
    defparam \uart_pc.state_RNO_0_2_LC_9_12_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_9_12_0 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_9_12_0  (
            .in0(N__36339),
            .in1(N__33250),
            .in2(N__33420),
            .in3(N__36894),
            .lcout(\uart_pc.state_srsts_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_12_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_9_12_1  (
            .in0(N__32326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32590),
            .lcout(\uart_drone.N_126_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__31636),
            .in2(_gnd_net_),
            .in3(N__31818),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_12_3  (
            .in0(N__33621),
            .in1(N__31311),
            .in2(N__31109),
            .in3(N__31158),
            .lcout(\Commands_frame_decoder.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNI3NPK_1_LC_9_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI3NPK_1_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI3NPK_1_LC_9_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI3NPK_1_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__33467),
            .in2(_gnd_net_),
            .in3(N__31078),
            .lcout(\Commands_frame_decoder.N_308_2 ),
            .ltout(\Commands_frame_decoder.N_308_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_9_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_9_12_7 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_9_12_7  (
            .in0(N__31045),
            .in1(N__32290),
            .in2(N__31034),
            .in3(N__32908),
            .lcout(\Commands_frame_decoder.state_ns_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_9_13_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_9_13_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_9_13_2  (
            .in0(N__31510),
            .in1(N__34324),
            .in2(_gnd_net_),
            .in3(N__36896),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_9_13_3 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_9_13_3 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_9_13_3  (
            .in0(N__32278),
            .in1(N__32628),
            .in2(N__31025),
            .in3(N__32466),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36102),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_13_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_13_7 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_9_13_7  (
            .in0(N__32587),
            .in1(N__32325),
            .in2(N__32467),
            .in3(N__32627),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_9_14_1 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_9_14_1 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.state_1_LC_9_14_1  (
            .in0(N__31254),
            .in1(N__31511),
            .in2(N__34352),
            .in3(N__36899),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36094),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_9_14_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_9_14_2 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_9_14_2  (
            .in0(N__37236),
            .in1(N__32649),
            .in2(N__32543),
            .in3(N__32597),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_9_14_3 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_9_14_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \uart_pc.data_0_LC_9_14_3  (
            .in0(N__31415),
            .in1(N__31866),
            .in2(N__36194),
            .in3(N__31726),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36094),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_9_14_4 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_9_14_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \uart_pc.data_5_LC_9_14_4  (
            .in0(N__31727),
            .in1(N__31964),
            .in2(N__31878),
            .in3(N__31307),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36094),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_9_14_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_9_14_5 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_9_14_5  (
            .in0(N__32534),
            .in1(N__34323),
            .in2(N__31256),
            .in3(N__36898),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_9_14_6 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_9_14_6 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_9_14_6  (
            .in0(N__31255),
            .in1(N__32650),
            .in2(N__31238),
            .in3(N__32598),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36094),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_9_14_7 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_9_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_9_14_7  (
            .in0(N__31235),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36094),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_9_15_1 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_9_15_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \uart_pc.data_3_LC_9_15_1  (
            .in0(N__31723),
            .in1(N__31143),
            .in2(N__35372),
            .in3(N__31880),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36087),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_15_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_15_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_9_15_2  (
            .in0(N__34331),
            .in1(N__31539),
            .in2(_gnd_net_),
            .in3(N__35020),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__33166),
            .in2(_gnd_net_),
            .in3(N__33492),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_9_15_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_9_15_5 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_9_15_5  (
            .in0(N__32600),
            .in1(N__37227),
            .in2(N__32542),
            .in3(N__32651),
            .lcout(\uart_drone.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_9_15_6 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_9_15_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_LC_9_15_6  (
            .in0(N__31879),
            .in1(N__31722),
            .in2(N__32753),
            .in3(N__31786),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36087),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_9_15_7 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_9_15_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \uart_pc.data_4_LC_9_15_7  (
            .in0(N__31721),
            .in1(N__33954),
            .in2(N__31653),
            .in3(N__32710),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36087),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_16_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_16_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_9_16_2  (
            .in0(N__37189),
            .in1(N__37118),
            .in2(_gnd_net_),
            .in3(N__37061),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_16_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_9_16_3  (
            .in0(N__37064),
            .in1(_gnd_net_),
            .in2(N__37132),
            .in3(N__37192),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_9_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_9_16_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_9_16_5  (
            .in0(N__37063),
            .in1(_gnd_net_),
            .in2(N__37131),
            .in3(N__37191),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_16_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_9_16_6  (
            .in0(N__37190),
            .in1(N__37119),
            .in2(_gnd_net_),
            .in3(N__37062),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_16_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_16_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__31555),
            .in2(_gnd_net_),
            .in3(N__31540),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_6_LC_9_17_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_9_17_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_6_LC_9_17_3  (
            .in0(N__32792),
            .in1(N__36352),
            .in2(N__31963),
            .in3(N__36234),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36067),
            .ce(),
            .sr(N__35675));
    defparam \uart_pc.data_Aux_7_LC_9_17_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_9_17_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_7_LC_9_17_4  (
            .in0(N__36235),
            .in1(N__31939),
            .in2(N__36356),
            .in3(N__33859),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36067),
            .ce(),
            .sr(N__35675));
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIH58S_8_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__32008),
            .in2(_gnd_net_),
            .in3(N__36893),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_18_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_18_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_9_18_1  (
            .in0(N__37193),
            .in1(N__37133),
            .in2(_gnd_net_),
            .in3(N__37051),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_9_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_9_19_0 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_9_19_0  (
            .in0(N__33312),
            .in1(N__33291),
            .in2(_gnd_net_),
            .in3(N__31901),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_9_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_9_19_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_9_19_2  (
            .in0(N__33030),
            .in1(N__33051),
            .in2(_gnd_net_),
            .in3(N__33130),
            .lcout(\dron_frame_decoder_1.WDT10lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_19_3  (
            .in0(N__32935),
            .in1(N__33100),
            .in2(N__33086),
            .in3(N__32920),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_9_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_9_19_4 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_9_19_4  (
            .in0(N__33115),
            .in1(N__32219),
            .in2(N__31910),
            .in3(N__31907),
            .lcout(\dron_frame_decoder_1.WDT10lt14_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_19_5 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_19_5  (
            .in0(N__33292),
            .in1(N__33313),
            .in2(N__31895),
            .in3(N__32417),
            .lcout(\dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_9_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_9_20_7 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_9_20_7  (
            .in0(N__33067),
            .in1(N__33031),
            .in2(N__33011),
            .in3(N__33052),
            .lcout(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_2_LC_9_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_9_22_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_9_22_5  (
            .in0(N__32107),
            .in1(N__32423),
            .in2(N__32213),
            .in3(N__32160),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36028),
            .ce(),
            .sr(N__36749));
    defparam \scaler_3.source_data_1_4_LC_9_24_4 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_4_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_4_LC_9_24_4 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_3.source_data_1_4_LC_9_24_4  (
            .in0(N__36969),
            .in1(N__32096),
            .in2(N__32026),
            .in3(N__32060),
            .lcout(scaler_3_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36016),
            .ce(),
            .sr(N__36756));
    defparam \Commands_frame_decoder.state_9_LC_10_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_10_10_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_9_LC_10_10_0  (
            .in0(N__31987),
            .in1(N__32009),
            .in2(_gnd_net_),
            .in3(N__32870),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36108),
            .ce(),
            .sr(N__36700));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_11_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_10_11_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_10_11_0  (
            .in0(N__33224),
            .in1(N__33202),
            .in2(N__33227),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_11_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_10_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__32327),
            .in2(_gnd_net_),
            .in3(N__31973),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_11_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_10_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__32599),
            .in2(_gnd_net_),
            .in3(N__31970),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_11_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_10_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__32643),
            .in2(_gnd_net_),
            .in3(N__31967),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_10_12_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_10_12_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_1_LC_10_12_2  (
            .in0(N__33191),
            .in1(N__32492),
            .in2(N__32261),
            .in3(N__35057),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36095),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_10_12_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_10_12_4 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_drone.timer_Count_0_LC_10_12_4  (
            .in0(N__33226),
            .in1(N__32491),
            .in2(N__32260),
            .in3(N__35056),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36095),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_10_12_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_10_12_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.timer_Count_4_LC_10_12_5  (
            .in0(N__35055),
            .in1(N__32259),
            .in2(N__32501),
            .in3(N__32429),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36095),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_10_12_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_10_12_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__32389),
            .in2(_gnd_net_),
            .in3(N__36883),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_10_12_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_10_12_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.timer_Count_2_LC_10_12_7  (
            .in0(N__35054),
            .in1(N__32258),
            .in2(N__32500),
            .in3(N__32333),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36095),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_13_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_13_1 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_10_13_1  (
            .in0(N__32464),
            .in1(N__32309),
            .in2(N__32279),
            .in3(N__37247),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIG8P51_2_LC_10_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIG8P51_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIG8P51_2_LC_10_13_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \Commands_frame_decoder.count_RNIG8P51_2_LC_10_13_2  (
            .in0(N__33629),
            .in1(N__33149),
            .in2(_gnd_net_),
            .in3(N__33490),
            .lcout(\Commands_frame_decoder.state_ns_i_a3_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIDLVE1_2_LC_10_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIDLVE1_2_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIDLVE1_2_LC_10_13_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \Commands_frame_decoder.count_RNIDLVE1_2_LC_10_13_3  (
            .in0(N__33491),
            .in1(N__33630),
            .in2(N__33159),
            .in3(N__36892),
            .lcout(\Commands_frame_decoder.count_RNIDLVE1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_10_13_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_10_13_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_10_13_4  (
            .in0(N__32642),
            .in1(N__32465),
            .in2(N__35065),
            .in3(N__32274),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_10_13_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_10_13_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_10_13_5  (
            .in0(N__35032),
            .in1(N__32242),
            .in2(N__32231),
            .in3(N__32228),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36088),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_10_13_6 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_10_13_6 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \uart_pc.state_2_LC_10_13_6  (
            .in0(N__35270),
            .in1(N__35348),
            .in2(N__33251),
            .in3(N__32660),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36088),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_10_14_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_10_14_0 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_10_14_0  (
            .in0(N__32588),
            .in1(N__32644),
            .in2(N__37240),
            .in3(N__32460),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_14_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_14_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_10_14_2  (
            .in0(N__33830),
            .in1(N__34472),
            .in2(_gnd_net_),
            .in3(N__34571),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_10_14_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_10_14_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_10_14_3  (
            .in0(N__35344),
            .in1(N__35269),
            .in2(N__33425),
            .in3(N__33903),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_10_14_4 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_10_14_4 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \uart_pc.state_3_LC_10_14_4  (
            .in0(N__35035),
            .in1(N__33971),
            .in2(N__32654),
            .in3(N__33424),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36079),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_14_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_10_14_5  (
            .in0(N__32645),
            .in1(N__37327),
            .in2(_gnd_net_),
            .in3(N__32589),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(\uart_drone.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_10_14_6 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_10_14_6 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \uart_drone.state_3_LC_10_14_6  (
            .in0(N__32552),
            .in1(N__32535),
            .in2(N__32510),
            .in3(N__35034),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36079),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_10_14_7 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_10_14_7 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \uart_drone.state_4_LC_10_14_7  (
            .in0(N__35033),
            .in1(N__32507),
            .in2(N__32499),
            .in3(N__37226),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36079),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_10_15_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_10_15_2 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_10_15_2  (
            .in0(N__35297),
            .in1(N__34757),
            .in2(N__34697),
            .in3(N__33901),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(\uart_pc.un1_state_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_1_LC_10_15_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_10_15_3 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \uart_pc.data_Aux_1_LC_10_15_3  (
            .in0(N__32749),
            .in1(N__32786),
            .in2(N__32756),
            .in3(N__36325),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36069),
            .ce(),
            .sr(N__35679));
    defparam \uart_pc.data_Aux_2_LC_10_15_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_10_15_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_pc.data_Aux_2_LC_10_15_4  (
            .in0(N__36326),
            .in1(N__32738),
            .in2(N__32728),
            .in3(N__36216),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36069),
            .ce(),
            .sr(N__35679));
    defparam \uart_pc.data_Aux_4_LC_10_15_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_10_15_6 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_pc.data_Aux_4_LC_10_15_6  (
            .in0(N__36327),
            .in1(N__32777),
            .in2(N__32711),
            .in3(N__36217),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36069),
            .ce(),
            .sr(N__35679));
    defparam \uart_pc.data_Aux_5_LC_10_15_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_10_15_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_pc.data_Aux_5_LC_10_15_7  (
            .in0(N__36218),
            .in1(N__32993),
            .in2(N__32695),
            .in3(N__36328),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36069),
            .ce(),
            .sr(N__35679));
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_10_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_10_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_4_LC_10_16_0  (
            .in0(N__33745),
            .in1(N__33328),
            .in2(N__33731),
            .in3(N__33343),
            .lcout(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_10_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_10_16_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Commands_frame_decoder.WDT_RNID7P31_6_LC_10_16_1  (
            .in0(N__33697),
            .in1(N__33775),
            .in2(_gnd_net_),
            .in3(N__33679),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_10_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_10_16_2 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_10_16_2  (
            .in0(N__33760),
            .in1(N__32666),
            .in2(N__32678),
            .in3(N__32675),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(\Commands_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_10_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_10_16_3 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \Commands_frame_decoder.preinit_RNIF92K5_LC_10_16_3  (
            .in0(N__32805),
            .in1(N__34040),
            .in2(N__32669),
            .in3(N__34010),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_10_16_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_10_16_4 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_10_16_4  (
            .in0(N__33678),
            .in1(N__33696),
            .in2(N__33662),
            .in3(N__33712),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_10_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_10_16_5 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_10_16_5  (
            .in0(N__34041),
            .in1(N__34011),
            .in2(N__33640),
            .in3(N__32890),
            .lcout(\Commands_frame_decoder.N_303_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_10_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_10_16_6 .LUT_INIT=16'b0000001100010011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_10_16_6  (
            .in0(N__32891),
            .in1(N__33617),
            .in2(N__34016),
            .in3(N__34042),
            .lcout(\Commands_frame_decoder.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_10_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_10_16_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_10_16_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_10_16_7  (
            .in0(N__32806),
            .in1(_gnd_net_),
            .in2(N__33641),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36059),
            .ce(),
            .sr(N__36722));
    defparam \uart_pc.state_RNIEAGS_4_LC_10_17_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_10_17_0 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_10_17_0  (
            .in0(N__33905),
            .in1(_gnd_net_),
            .in2(N__34756),
            .in3(N__36886),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_17_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_17_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_10_17_1  (
            .in0(N__34560),
            .in1(N__33814),
            .in2(_gnd_net_),
            .in3(N__34452),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_10_17_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_10_17_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_10_17_2  (
            .in0(N__33812),
            .in1(N__34450),
            .in2(_gnd_net_),
            .in3(N__34558),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_17_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_17_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_10_17_3  (
            .in0(N__34559),
            .in1(N__33813),
            .in2(_gnd_net_),
            .in3(N__34451),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_10_17_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_10_17_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_10_17_5  (
            .in0(N__35326),
            .in1(_gnd_net_),
            .in2(N__35264),
            .in3(N__33858),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_10_17_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_10_17_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_10_17_6  (
            .in0(N__37185),
            .in1(N__37127),
            .in2(_gnd_net_),
            .in3(N__37043),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_10_17_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_10_17_7 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_10_17_7  (
            .in0(N__35325),
            .in1(N__34747),
            .in2(N__35263),
            .in3(N__33904),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_18_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_18_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_10_18_3  (
            .in0(N__33811),
            .in1(N__34449),
            .in2(_gnd_net_),
            .in3(N__34547),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_10_18_5 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_10_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__34500),
            .in2(_gnd_net_),
            .in3(N__34548),
            .lcout(\uart_pc.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_10_18_7 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_10_18_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_10_18_7  (
            .in0(N__33810),
            .in1(N__34448),
            .in2(_gnd_net_),
            .in3(N__34546),
            .lcout(\uart_pc.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_10_19_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_10_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__32969),
            .in2(N__32984),
            .in3(N__32983),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_1_LC_10_19_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_10_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__32963),
            .in2(_gnd_net_),
            .in3(N__32957),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_2_LC_10_19_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_10_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__32954),
            .in2(_gnd_net_),
            .in3(N__32948),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_3_LC_10_19_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_10_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__32945),
            .in2(_gnd_net_),
            .in3(N__32939),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_4_LC_10_19_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_10_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__32936),
            .in2(_gnd_net_),
            .in3(N__32924),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_5_LC_10_19_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_10_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__32921),
            .in2(_gnd_net_),
            .in3(N__33134),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_6_LC_10_19_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_10_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__33131),
            .in2(_gnd_net_),
            .in3(N__33119),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_7_LC_10_19_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_10_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__33116),
            .in2(_gnd_net_),
            .in3(N__33104),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__36039),
            .ce(),
            .sr(N__33277));
    defparam \dron_frame_decoder_1.WDT_8_LC_10_20_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_10_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__33101),
            .in2(_gnd_net_),
            .in3(N__33089),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_9_LC_10_20_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_10_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__33085),
            .in2(_gnd_net_),
            .in3(N__33071),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_10_LC_10_20_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_10_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__33068),
            .in2(_gnd_net_),
            .in3(N__33056),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_11_LC_10_20_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_10_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__33053),
            .in2(_gnd_net_),
            .in3(N__33035),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_12_LC_10_20_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_10_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__33032),
            .in2(_gnd_net_),
            .in3(N__33014),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_13_LC_10_20_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_10_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(_gnd_net_),
            .in3(N__32996),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_14_LC_10_20_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_10_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__33314),
            .in2(_gnd_net_),
            .in3(N__33299),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \dron_frame_decoder_1.WDT_15_LC_10_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_10_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__33293),
            .in2(_gnd_net_),
            .in3(N__33296),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36030),
            .ce(),
            .sr(N__33278));
    defparam \uart_pc.state_1_LC_11_12_1 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_11_12_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_11_12_1  (
            .in0(N__33249),
            .in1(N__36343),
            .in2(N__34718),
            .in3(N__36910),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36089),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_11_12_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_11_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__33225),
            .in2(_gnd_net_),
            .in3(N__33203),
            .lcout(\uart_drone.timer_Count_RNO_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_13_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_13_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_11_13_1  (
            .in0(N__33826),
            .in1(N__34467),
            .in2(_gnd_net_),
            .in3(N__34566),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIE6P51_0_LC_11_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIE6P51_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIE6P51_0_LC_11_14_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Commands_frame_decoder.count_RNIE6P51_0_LC_11_14_0  (
            .in0(N__33433),
            .in1(N__33612),
            .in2(_gnd_net_),
            .in3(N__33493),
            .lcout(\Commands_frame_decoder.CO0 ),
            .ltout(\Commands_frame_decoder.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_1_LC_11_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_1_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_1_LC_11_14_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \Commands_frame_decoder.count_1_LC_11_14_1  (
            .in0(N__33448),
            .in1(_gnd_net_),
            .in2(N__33185),
            .in3(N__33175),
            .lcout(\Commands_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36070),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_11_14_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_11_14_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_11_14_2  (
            .in0(N__33825),
            .in1(N__34466),
            .in2(_gnd_net_),
            .in3(N__34565),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_2_LC_11_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_2_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_2_LC_11_14_3 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \Commands_frame_decoder.count_2_LC_11_14_3  (
            .in0(N__33449),
            .in1(N__33182),
            .in2(N__33167),
            .in3(N__33176),
            .lcout(\Commands_frame_decoder.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_11_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_11_14_4 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_11_14_4  (
            .in0(N__33613),
            .in1(N__33494),
            .in2(N__33437),
            .in3(N__33447),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36070),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_14_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_14_6 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_11_14_6  (
            .in0(N__35268),
            .in1(N__35337),
            .in2(N__33419),
            .in3(N__33902),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_11_15_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33377),
            .in2(N__33392),
            .in3(N__33391),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_1_LC_11_15_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__33371),
            .in2(_gnd_net_),
            .in3(N__33365),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_2_LC_11_15_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__33362),
            .in2(_gnd_net_),
            .in3(N__33356),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_3_LC_11_15_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__33353),
            .in2(_gnd_net_),
            .in3(N__33347),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_4_LC_11_15_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_11_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33344),
            .in2(_gnd_net_),
            .in3(N__33332),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_5_LC_11_15_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_11_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__33329),
            .in2(_gnd_net_),
            .in3(N__33317),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_6_LC_11_15_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__33776),
            .in2(_gnd_net_),
            .in3(N__33764),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_7_LC_11_15_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__33761),
            .in2(_gnd_net_),
            .in3(N__33749),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__36060),
            .ce(),
            .sr(N__33991));
    defparam \Commands_frame_decoder.WDT_8_LC_11_16_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_11_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__33746),
            .in2(_gnd_net_),
            .in3(N__33734),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_9_LC_11_16_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_11_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__33730),
            .in2(_gnd_net_),
            .in3(N__33716),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_10_LC_11_16_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_11_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__33713),
            .in2(_gnd_net_),
            .in3(N__33701),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_11_LC_11_16_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__33698),
            .in2(_gnd_net_),
            .in3(N__33683),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_12_LC_11_16_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_11_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__33680),
            .in2(_gnd_net_),
            .in3(N__33665),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_13_LC_11_16_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_11_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__33661),
            .in2(_gnd_net_),
            .in3(N__33647),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_14_LC_11_16_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_11_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__34043),
            .in2(_gnd_net_),
            .in3(N__34022),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \Commands_frame_decoder.WDT_15_LC_11_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_11_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__34015),
            .in2(_gnd_net_),
            .in3(N__34019),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36053),
            .ce(),
            .sr(N__33995));
    defparam \uart_pc.state_4_LC_11_17_0 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_11_17_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \uart_pc.state_4_LC_11_17_0  (
            .in0(N__33907),
            .in1(N__33970),
            .in2(N__35064),
            .in3(N__35152),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36046),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_17_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_17_1 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_11_17_1  (
            .in0(N__35184),
            .in1(N__35324),
            .in2(N__35246),
            .in3(N__34746),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_11_17_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_11_17_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_11_17_2  (
            .in0(N__37175),
            .in1(N__37126),
            .in2(_gnd_net_),
            .in3(N__37042),
            .lcout(\uart_drone.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_11_17_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_11_17_5 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_11_17_5  (
            .in0(N__34499),
            .in1(N__33906),
            .in2(_gnd_net_),
            .in3(N__33857),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_11_17_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_11_17_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_3_LC_11_17_7  (
            .in0(N__35058),
            .in1(N__35114),
            .in2(N__35156),
            .in3(N__34679),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36046),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_0_LC_11_18_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_11_18_0 .LUT_INIT=16'b0011000000111000;
    LogicCell40 \uart_pc.bit_Count_0_LC_11_18_0  (
            .in0(N__33911),
            .in1(N__34504),
            .in2(N__34570),
            .in3(N__33860),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36040),
            .ce(),
            .sr(N__36733));
    defparam \uart_pc.bit_Count_2_LC_11_18_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_11_18_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_11_18_2  (
            .in0(N__34481),
            .in1(N__33824),
            .in2(N__34471),
            .in3(N__33836),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36040),
            .ce(),
            .sr(N__36733));
    defparam \uart_pc.bit_Count_1_LC_11_18_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_11_18_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uart_pc.bit_Count_1_LC_11_18_3  (
            .in0(N__34561),
            .in1(N__34462),
            .in2(N__34505),
            .in3(N__34480),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36040),
            .ce(),
            .sr(N__36733));
    defparam \uart_drone.data_Aux_7_LC_11_19_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_11_19_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_11_19_1  (
            .in0(N__34378),
            .in1(N__34270),
            .in2(N__34405),
            .in3(N__37325),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36031),
            .ce(),
            .sr(N__34201));
    defparam \uart_drone.data_Aux_4_LC_11_20_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_11_20_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_4_LC_11_20_6  (
            .in0(N__36989),
            .in1(N__34377),
            .in2(N__34219),
            .in3(N__34274),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36021),
            .ce(),
            .sr(N__34202));
    defparam \pid_alt.state_RNIH1EN_0_LC_12_2_2 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_2_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__34166),
            .in2(_gnd_net_),
            .in3(N__36878),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_12_12_0 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_12_12_0 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \reset_module_System.count_2_LC_12_12_0  (
            .in0(N__35548),
            .in1(N__34052),
            .in2(N__35468),
            .in3(N__35565),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36078),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_12_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_12_12_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_12_12_2  (
            .in0(N__34601),
            .in1(N__34622),
            .in2(N__34643),
            .in3(N__34064),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(\reset_module_System.reset6_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_12_12_3 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_12_12_3 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \reset_module_System.reset_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__35464),
            .in2(N__34067),
            .in3(N__35547),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36078),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_12_13_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__35534),
            .in2(N__35588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_12_13_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_12_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__34063),
            .in2(_gnd_net_),
            .in3(N__34046),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_12_13_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_12_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__34621),
            .in2(_gnd_net_),
            .in3(N__34610),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_12_13_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_12_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__34772),
            .in2(_gnd_net_),
            .in3(N__34607),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_12_13_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_12_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__34798),
            .in2(_gnd_net_),
            .in3(N__34604),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_12_13_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_12_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__34600),
            .in2(_gnd_net_),
            .in3(N__34589),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_12_13_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_12_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__34814),
            .in2(_gnd_net_),
            .in3(N__34586),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_12_13_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_12_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__34826),
            .in2(_gnd_net_),
            .in3(N__34583),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__36068),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_12_14_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_12_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__34784),
            .in2(_gnd_net_),
            .in3(N__34580),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_12_14_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_12_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__35479),
            .in2(_gnd_net_),
            .in3(N__34577),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_12_14_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_12_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__35506),
            .in2(_gnd_net_),
            .in3(N__34574),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_12_14_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_12_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__35605),
            .in2(_gnd_net_),
            .in3(N__34667),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_12_14_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_12_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__35402),
            .in2(_gnd_net_),
            .in3(N__34664),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_12_14_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_12_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__35518),
            .in2(_gnd_net_),
            .in3(N__34661),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_12_14_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_12_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__35429),
            .in2(_gnd_net_),
            .in3(N__34658),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_12_14_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_12_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__35630),
            .in2(_gnd_net_),
            .in3(N__34655),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__36058),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_12_15_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_12_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__35491),
            .in2(_gnd_net_),
            .in3(N__34652),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__36052),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_12_15_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_12_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__35644),
            .in2(_gnd_net_),
            .in3(N__34649),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__36052),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_12_15_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_12_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__35441),
            .in2(_gnd_net_),
            .in3(N__34646),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__36052),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_12_15_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_12_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__34639),
            .in2(_gnd_net_),
            .in3(N__34625),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__36052),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_12_15_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_12_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__35416),
            .in2(_gnd_net_),
            .in3(N__34760),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36052),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_12_16_1 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_12_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__37028),
            .in2(_gnd_net_),
            .in3(N__37286),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_12_16_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_12_16_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_12_16_4  (
            .in0(N__35292),
            .in1(N__34751),
            .in2(N__35256),
            .in3(N__35021),
            .lcout(\uart_pc.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_12_16_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_12_16_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_12_16_6  (
            .in0(N__34708),
            .in1(N__36351),
            .in2(_gnd_net_),
            .in3(N__36897),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_12_16_7 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_12_16_7 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart_pc.state_0_LC_12_16_7  (
            .in0(N__34752),
            .in1(N__35240),
            .in2(N__34721),
            .in3(N__35293),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36045),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_12_17_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_12_17_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_12_17_0  (
            .in0(N__34847),
            .in1(N__35167),
            .in2(N__34850),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_12_17_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_12_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35189),
            .in3(N__34682),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_12_17_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_12_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__35328),
            .in2(_gnd_net_),
            .in3(N__34673),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_12_17_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_12_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__35236),
            .in2(_gnd_net_),
            .in3(N__34670),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_17_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__35327),
            .in2(_gnd_net_),
            .in3(N__35185),
            .lcout(\uart_pc.N_126_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_12_17_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_12_17_6 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_4_LC_12_17_6  (
            .in0(N__35022),
            .in1(N__35108),
            .in2(N__35155),
            .in3(N__35276),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36038),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_12_17_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_12_17_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_2_LC_12_17_7  (
            .in0(N__35195),
            .in1(N__35145),
            .in2(N__35115),
            .in3(N__35023),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36038),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_12_18_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__34848),
            .in2(_gnd_net_),
            .in3(N__35168),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_12_18_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_12_18_5 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \uart_pc.timer_Count_1_LC_12_18_5  (
            .in0(N__35154),
            .in1(N__35024),
            .in2(N__35171),
            .in3(N__35119),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36029),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_12_18_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_12_18_6 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_12_18_6  (
            .in0(N__34849),
            .in1(N__35153),
            .in2(N__35120),
            .in3(N__35025),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36029),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_13_13_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_13_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_13_13_0  (
            .in0(N__34825),
            .in1(N__34813),
            .in2(N__34802),
            .in3(N__34783),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_13_13_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_13_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__34771),
            .in2(_gnd_net_),
            .in3(N__35532),
            .lcout(),
            .ltout(\reset_module_System.reset6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_13_13_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_13_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_13_13_3  (
            .in0(N__35645),
            .in1(N__35629),
            .in2(N__35618),
            .in3(N__35615),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_13_13_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_13_13_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_13_13_4  (
            .in0(N__35390),
            .in1(N__35609),
            .in2(N__35594),
            .in3(N__35585),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_13_13_5 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_13_13_5 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_13_13_5  (
            .in0(N__35587),
            .in1(N__35566),
            .in2(N__35591),
            .in3(N__35463),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36080),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_13_13_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_13_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__35586),
            .in2(_gnd_net_),
            .in3(N__35533),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_13_13_7 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_13_13_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_13_13_7  (
            .in0(N__35462),
            .in1(N__35567),
            .in2(N__35552),
            .in3(N__35549),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36080),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_13_14_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_13_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_13_14_5  (
            .in0(N__35519),
            .in1(N__35507),
            .in2(N__35495),
            .in3(N__35480),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_14_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_13_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_13_14_6  (
            .in0(N__35440),
            .in1(N__35428),
            .in2(N__35417),
            .in3(N__35401),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_3_LC_13_15_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_13_15_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_3_LC_13_15_2  (
            .in0(N__35384),
            .in1(N__36344),
            .in2(N__35365),
            .in3(N__36230),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36061),
            .ce(),
            .sr(N__35683));
    defparam \uart_drone.state_RNI63LK2_3_LC_13_16_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_13_16_0 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_13_16_0  (
            .in0(N__37287),
            .in1(N__37328),
            .in2(_gnd_net_),
            .in3(N__37251),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(\uart_drone.un1_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_13_16_1 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_13_16_1 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \uart_drone.bit_Count_1_LC_13_16_1  (
            .in0(N__37106),
            .in1(N__37041),
            .in2(N__37346),
            .in3(N__37288),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36054),
            .ce(),
            .sr(N__36734));
    defparam \uart_drone.bit_Count_2_LC_13_16_3 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_13_16_3 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \uart_drone.bit_Count_2_LC_13_16_3  (
            .in0(N__37107),
            .in1(N__37161),
            .in2(N__37343),
            .in3(N__37334),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36054),
            .ce(),
            .sr(N__36734));
    defparam \uart_drone.bit_Count_0_LC_13_17_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_13_17_6 .LUT_INIT=16'b0011010000110000;
    LogicCell40 \uart_drone.bit_Count_0_LC_13_17_6  (
            .in0(N__37326),
            .in1(N__37289),
            .in2(N__37050),
            .in3(N__37256),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36047),
            .ce(),
            .sr(N__36738));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_13_18_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_13_18_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_13_18_6  (
            .in0(N__37174),
            .in1(N__37117),
            .in2(_gnd_net_),
            .in3(N__37029),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_23_0 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_23_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_2.source_data_1_esr_ctle_14_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__36965),
            .in2(_gnd_net_),
            .in3(N__36876),
            .lcout(debug_CH3_20A_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_14_15_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_14_15_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_14_15_2  (
            .in0(N__36368),
            .in1(N__36345),
            .in2(N__36184),
            .in3(N__36236),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36071),
            .ce(),
            .sr(N__35684));
endmodule // Pc2drone
