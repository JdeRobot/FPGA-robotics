// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 16 2019 21:18:00

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2Drone" view "INTERFACE"

module Pc2Drone (
    ppm_output,
    uart_input_debug,
    uart_input,
    frame_decoder_dv,
    clk_system);

    output ppm_output;
    output uart_input_debug;
    input uart_input;
    output frame_decoder_dv;
    input clk_system;

    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24838;
    wire N__24837;
    wire N__24836;
    wire N__24829;
    wire N__24828;
    wire N__24827;
    wire N__24820;
    wire N__24819;
    wire N__24818;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24770;
    wire N__24769;
    wire N__24768;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24747;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24742;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24716;
    wire N__24713;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24690;
    wire N__24687;
    wire N__24682;
    wire N__24679;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24660;
    wire N__24651;
    wire N__24644;
    wire N__24641;
    wire N__24634;
    wire N__24629;
    wire N__24624;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24587;
    wire N__24582;
    wire N__24579;
    wire N__24578;
    wire N__24577;
    wire N__24570;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24558;
    wire N__24555;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24534;
    wire N__24533;
    wire N__24530;
    wire N__24529;
    wire N__24528;
    wire N__24525;
    wire N__24524;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24487;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24467;
    wire N__24464;
    wire N__24463;
    wire N__24462;
    wire N__24457;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24411;
    wire N__24408;
    wire N__24407;
    wire N__24406;
    wire N__24405;
    wire N__24402;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24394;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24379;
    wire N__24374;
    wire N__24371;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24347;
    wire N__24346;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24240;
    wire N__24237;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24208;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24178;
    wire N__24165;
    wire N__24162;
    wire N__24161;
    wire N__24158;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24147;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24131;
    wire N__24126;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24118;
    wire N__24117;
    wire N__24116;
    wire N__24113;
    wire N__24108;
    wire N__24103;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24089;
    wire N__24088;
    wire N__24087;
    wire N__24086;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24078;
    wire N__24077;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24069;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24041;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24025;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24006;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23982;
    wire N__23981;
    wire N__23980;
    wire N__23977;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23960;
    wire N__23959;
    wire N__23956;
    wire N__23947;
    wire N__23944;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23920;
    wire N__23911;
    wire N__23908;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23882;
    wire N__23881;
    wire N__23880;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23876;
    wire N__23875;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23860;
    wire N__23859;
    wire N__23858;
    wire N__23857;
    wire N__23856;
    wire N__23855;
    wire N__23854;
    wire N__23853;
    wire N__23852;
    wire N__23851;
    wire N__23850;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23846;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23841;
    wire N__23840;
    wire N__23839;
    wire N__23838;
    wire N__23837;
    wire N__23836;
    wire N__23835;
    wire N__23834;
    wire N__23833;
    wire N__23832;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23823;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23815;
    wire N__23814;
    wire N__23813;
    wire N__23812;
    wire N__23811;
    wire N__23810;
    wire N__23809;
    wire N__23808;
    wire N__23807;
    wire N__23806;
    wire N__23805;
    wire N__23804;
    wire N__23803;
    wire N__23802;
    wire N__23801;
    wire N__23800;
    wire N__23799;
    wire N__23798;
    wire N__23797;
    wire N__23796;
    wire N__23795;
    wire N__23794;
    wire N__23793;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23789;
    wire N__23788;
    wire N__23787;
    wire N__23786;
    wire N__23785;
    wire N__23784;
    wire N__23783;
    wire N__23782;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23570;
    wire N__23569;
    wire N__23568;
    wire N__23567;
    wire N__23566;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23562;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23534;
    wire N__23533;
    wire N__23532;
    wire N__23531;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23523;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23490;
    wire N__23487;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23450;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23405;
    wire N__23404;
    wire N__23403;
    wire N__23402;
    wire N__23401;
    wire N__23400;
    wire N__23399;
    wire N__23398;
    wire N__23397;
    wire N__23396;
    wire N__23395;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23387;
    wire N__23386;
    wire N__23385;
    wire N__23384;
    wire N__23383;
    wire N__23382;
    wire N__23381;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23364;
    wire N__23363;
    wire N__23362;
    wire N__23361;
    wire N__23360;
    wire N__23359;
    wire N__23358;
    wire N__23357;
    wire N__23356;
    wire N__23355;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23351;
    wire N__23350;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23018;
    wire N__23017;
    wire N__23014;
    wire N__23009;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22967;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22937;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22863;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22841;
    wire N__22840;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22836;
    wire N__22835;
    wire N__22832;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22814;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22763;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22733;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22689;
    wire N__22684;
    wire N__22681;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22577;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22549;
    wire N__22544;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22526;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22495;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22469;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22427;
    wire N__22424;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22368;
    wire N__22367;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22350;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22329;
    wire N__22328;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22311;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22287;
    wire N__22284;
    wire N__22283;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22258;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22235;
    wire N__22232;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22154;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22134;
    wire N__22133;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22122;
    wire N__22121;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22117;
    wire N__22116;
    wire N__22111;
    wire N__22110;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22098;
    wire N__22097;
    wire N__22096;
    wire N__22091;
    wire N__22084;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22068;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22058;
    wire N__22053;
    wire N__22050;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22020;
    wire N__22015;
    wire N__22008;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21982;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21973;
    wire N__21968;
    wire N__21967;
    wire N__21966;
    wire N__21965;
    wire N__21964;
    wire N__21961;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21925;
    wire N__21920;
    wire N__21915;
    wire N__21908;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21896;
    wire N__21893;
    wire N__21888;
    wire N__21883;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21864;
    wire N__21861;
    wire N__21856;
    wire N__21849;
    wire N__21844;
    wire N__21831;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21786;
    wire N__21785;
    wire N__21782;
    wire N__21781;
    wire N__21780;
    wire N__21779;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21762;
    wire N__21761;
    wire N__21760;
    wire N__21753;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21734;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21703;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21691;
    wire N__21688;
    wire N__21687;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21679;
    wire N__21676;
    wire N__21669;
    wire N__21666;
    wire N__21659;
    wire N__21654;
    wire N__21651;
    wire N__21644;
    wire N__21637;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21615;
    wire N__21614;
    wire N__21611;
    wire N__21610;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21594;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21571;
    wire N__21566;
    wire N__21563;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21545;
    wire N__21540;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21513;
    wire N__21512;
    wire N__21511;
    wire N__21508;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21484;
    wire N__21481;
    wire N__21476;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21450;
    wire N__21449;
    wire N__21446;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21276;
    wire N__21273;
    wire N__21272;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21234;
    wire N__21233;
    wire N__21232;
    wire N__21231;
    wire N__21230;
    wire N__21229;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21223;
    wire N__21222;
    wire N__21221;
    wire N__21220;
    wire N__21219;
    wire N__21218;
    wire N__21217;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21207;
    wire N__21206;
    wire N__21205;
    wire N__21204;
    wire N__21203;
    wire N__21202;
    wire N__21201;
    wire N__21192;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21155;
    wire N__21146;
    wire N__21145;
    wire N__21140;
    wire N__21131;
    wire N__21130;
    wire N__21123;
    wire N__21120;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21090;
    wire N__21089;
    wire N__21088;
    wire N__21087;
    wire N__21086;
    wire N__21085;
    wire N__21084;
    wire N__21083;
    wire N__21080;
    wire N__21073;
    wire N__21070;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21053;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21021;
    wire N__21010;
    wire N__21005;
    wire N__21002;
    wire N__20993;
    wire N__20984;
    wire N__20979;
    wire N__20970;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20930;
    wire N__20927;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20894;
    wire N__20889;
    wire N__20886;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20817;
    wire N__20816;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20777;
    wire N__20772;
    wire N__20771;
    wire N__20770;
    wire N__20767;
    wire N__20762;
    wire N__20757;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20736;
    wire N__20733;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20663;
    wire N__20660;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20592;
    wire N__20591;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20540;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20515;
    wire N__20512;
    wire N__20507;
    wire N__20502;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20450;
    wire N__20449;
    wire N__20444;
    wire N__20441;
    wire N__20440;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20421;
    wire N__20420;
    wire N__20419;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20392;
    wire N__20391;
    wire N__20388;
    wire N__20381;
    wire N__20376;
    wire N__20371;
    wire N__20368;
    wire N__20363;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20351;
    wire N__20350;
    wire N__20349;
    wire N__20348;
    wire N__20347;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20342;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20321;
    wire N__20316;
    wire N__20311;
    wire N__20302;
    wire N__20299;
    wire N__20294;
    wire N__20287;
    wire N__20274;
    wire N__20273;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20258;
    wire N__20257;
    wire N__20256;
    wire N__20255;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20243;
    wire N__20242;
    wire N__20241;
    wire N__20240;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20222;
    wire N__20219;
    wire N__20218;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20203;
    wire N__20200;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20182;
    wire N__20177;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20152;
    wire N__20151;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20116;
    wire N__20115;
    wire N__20110;
    wire N__20105;
    wire N__20104;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20072;
    wire N__20067;
    wire N__20060;
    wire N__20043;
    wire N__20040;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20018;
    wire N__20015;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19988;
    wire N__19985;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19973;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19937;
    wire N__19932;
    wire N__19931;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19862;
    wire N__19861;
    wire N__19860;
    wire N__19859;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19844;
    wire N__19841;
    wire N__19830;
    wire N__19827;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19790;
    wire N__19785;
    wire N__19770;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19766;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19746;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19706;
    wire N__19705;
    wire N__19702;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19690;
    wire N__19689;
    wire N__19688;
    wire N__19687;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19655;
    wire N__19650;
    wire N__19643;
    wire N__19632;
    wire N__19631;
    wire N__19630;
    wire N__19627;
    wire N__19626;
    wire N__19625;
    wire N__19624;
    wire N__19623;
    wire N__19622;
    wire N__19621;
    wire N__19620;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19598;
    wire N__19597;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19591;
    wire N__19588;
    wire N__19587;
    wire N__19582;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19558;
    wire N__19555;
    wire N__19554;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19548;
    wire N__19541;
    wire N__19540;
    wire N__19539;
    wire N__19538;
    wire N__19533;
    wire N__19526;
    wire N__19521;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19502;
    wire N__19497;
    wire N__19492;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19468;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19444;
    wire N__19441;
    wire N__19436;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19410;
    wire N__19407;
    wire N__19406;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19374;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19338;
    wire N__19337;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19296;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19266;
    wire N__19263;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19239;
    wire N__19236;
    wire N__19235;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19014;
    wire N__19011;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18921;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18903;
    wire N__18902;
    wire N__18901;
    wire N__18900;
    wire N__18899;
    wire N__18898;
    wire N__18897;
    wire N__18894;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18886;
    wire N__18885;
    wire N__18882;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18876;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18860;
    wire N__18855;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18827;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18805;
    wire N__18802;
    wire N__18789;
    wire N__18788;
    wire N__18787;
    wire N__18784;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18776;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18764;
    wire N__18763;
    wire N__18760;
    wire N__18759;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18735;
    wire N__18732;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18687;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18590;
    wire N__18589;
    wire N__18586;
    wire N__18581;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18571;
    wire N__18568;
    wire N__18563;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18551;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18534;
    wire N__18533;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18516;
    wire N__18513;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18494;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18449;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18419;
    wire N__18414;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18392;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18290;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18253;
    wire N__18250;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18145;
    wire N__18140;
    wire N__18137;
    wire N__18132;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18040;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17872;
    wire N__17871;
    wire N__17866;
    wire N__17865;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17850;
    wire N__17847;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17817;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17808;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17782;
    wire N__17777;
    wire N__17772;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17737;
    wire N__17736;
    wire N__17735;
    wire N__17730;
    wire N__17723;
    wire N__17718;
    wire N__17717;
    wire N__17716;
    wire N__17715;
    wire N__17714;
    wire N__17713;
    wire N__17712;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17705;
    wire N__17704;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17669;
    wire N__17668;
    wire N__17667;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17637;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17618;
    wire N__17613;
    wire N__17604;
    wire N__17601;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17568;
    wire N__17565;
    wire N__17564;
    wire N__17563;
    wire N__17562;
    wire N__17561;
    wire N__17560;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17541;
    wire N__17540;
    wire N__17539;
    wire N__17536;
    wire N__17535;
    wire N__17534;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17524;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17496;
    wire N__17493;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17476;
    wire N__17473;
    wire N__17468;
    wire N__17463;
    wire N__17462;
    wire N__17461;
    wire N__17460;
    wire N__17459;
    wire N__17458;
    wire N__17455;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17435;
    wire N__17434;
    wire N__17433;
    wire N__17432;
    wire N__17429;
    wire N__17414;
    wire N__17411;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17390;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17367;
    wire N__17364;
    wire N__17359;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17325;
    wire N__17310;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17301;
    wire N__17296;
    wire N__17293;
    wire N__17288;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17192;
    wire N__17189;
    wire N__17188;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17182;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17162;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17088;
    wire N__17087;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17037;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17007;
    wire N__17002;
    wire N__16997;
    wire N__16994;
    wire N__16989;
    wire N__16984;
    wire N__16981;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16922;
    wire N__16921;
    wire N__16920;
    wire N__16919;
    wire N__16918;
    wire N__16915;
    wire N__16914;
    wire N__16911;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16896;
    wire N__16889;
    wire N__16882;
    wire N__16881;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16877;
    wire N__16876;
    wire N__16875;
    wire N__16872;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16843;
    wire N__16838;
    wire N__16833;
    wire N__16826;
    wire N__16823;
    wire N__16816;
    wire N__16813;
    wire N__16800;
    wire N__16799;
    wire N__16798;
    wire N__16797;
    wire N__16796;
    wire N__16795;
    wire N__16794;
    wire N__16793;
    wire N__16792;
    wire N__16791;
    wire N__16790;
    wire N__16789;
    wire N__16788;
    wire N__16787;
    wire N__16786;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16767;
    wire N__16762;
    wire N__16759;
    wire N__16748;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16262;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16250;
    wire N__16245;
    wire N__16244;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16193;
    wire N__16188;
    wire N__16185;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15867;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15806;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15740;
    wire N__15737;
    wire N__15732;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15674;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15651;
    wire N__15650;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15629;
    wire N__15626;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15371;
    wire N__15368;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15311;
    wire N__15310;
    wire N__15307;
    wire N__15302;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15267;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15230;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15222;
    wire N__15219;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15195;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15153;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15135;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15095;
    wire N__15094;
    wire N__15093;
    wire N__15090;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15073;
    wire N__15070;
    wire N__15061;
    wire N__15058;
    wire N__15057;
    wire N__15056;
    wire N__15053;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14939;
    wire N__14934;
    wire N__14933;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14906;
    wire N__14901;
    wire N__14896;
    wire N__14893;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14793;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14781;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14769;
    wire N__14766;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14747;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14696;
    wire N__14691;
    wire N__14688;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14676;
    wire N__14675;
    wire N__14672;
    wire N__14667;
    wire N__14664;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14652;
    wire N__14649;
    wire N__14648;
    wire N__14647;
    wire N__14646;
    wire N__14641;
    wire N__14636;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14607;
    wire N__14606;
    wire N__14603;
    wire N__14602;
    wire N__14599;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14587;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14472;
    wire N__14469;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14457;
    wire N__14454;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14442;
    wire N__14439;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14427;
    wire N__14424;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14412;
    wire N__14409;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14397;
    wire N__14394;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14379;
    wire N__14376;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14364;
    wire N__14361;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14349;
    wire N__14346;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14327;
    wire N__14326;
    wire N__14325;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14311;
    wire N__14308;
    wire N__14301;
    wire N__14298;
    wire N__14297;
    wire N__14292;
    wire N__14291;
    wire N__14290;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14268;
    wire N__14265;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14249;
    wire N__14248;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14233;
    wire N__14228;
    wire N__14227;
    wire N__14224;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14197;
    wire N__14184;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14148;
    wire N__14145;
    wire N__14144;
    wire N__14143;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14125;
    wire N__14118;
    wire N__14117;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14100;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14081;
    wire N__14080;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14058;
    wire N__14057;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14034;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13973;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13950;
    wire N__13949;
    wire N__13948;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13936;
    wire N__13929;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13921;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13909;
    wire N__13902;
    wire N__13899;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13797;
    wire N__13794;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13782;
    wire N__13779;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13593;
    wire N__13590;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13560;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13509;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13473;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13461;
    wire N__13460;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13368;
    wire N__13361;
    wire N__13360;
    wire N__13355;
    wire N__13352;
    wire N__13347;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13329;
    wire N__13326;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13290;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13254;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13246;
    wire N__13241;
    wire N__13238;
    wire N__13237;
    wire N__13236;
    wire N__13235;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13218;
    wire N__13209;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13169;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13161;
    wire N__13158;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13149;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13110;
    wire N__13107;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13099;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13062;
    wire N__13061;
    wire N__13054;
    wire N__13051;
    wire N__13044;
    wire N__13039;
    wire N__13032;
    wire N__13027;
    wire N__13020;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12993;
    wire N__12992;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12982;
    wire N__12981;
    wire N__12978;
    wire N__12977;
    wire N__12976;
    wire N__12975;
    wire N__12974;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12950;
    wire N__12939;
    wire N__12936;
    wire N__12935;
    wire N__12930;
    wire N__12929;
    wire N__12926;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12921;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12907;
    wire N__12904;
    wire N__12899;
    wire N__12892;
    wire N__12879;
    wire N__12878;
    wire N__12877;
    wire N__12876;
    wire N__12871;
    wire N__12866;
    wire N__12863;
    wire N__12862;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12858;
    wire N__12857;
    wire N__12856;
    wire N__12855;
    wire N__12850;
    wire N__12847;
    wire N__12842;
    wire N__12831;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12779;
    wire N__12778;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12752;
    wire N__12745;
    wire N__12742;
    wire N__12741;
    wire N__12740;
    wire N__12739;
    wire N__12736;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12704;
    wire N__12699;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12681;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12659;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12644;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12634;
    wire N__12633;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12603;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12595;
    wire N__12592;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12571;
    wire N__12564;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12528;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12509;
    wire N__12500;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12490;
    wire N__12487;
    wire N__12484;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12402;
    wire N__12399;
    wire N__12398;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12369;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12361;
    wire N__12356;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12334;
    wire N__12329;
    wire N__12326;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12292;
    wire N__12285;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12277;
    wire N__12276;
    wire N__12275;
    wire N__12274;
    wire N__12273;
    wire N__12272;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12250;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12215;
    wire N__12214;
    wire N__12213;
    wire N__12210;
    wire N__12209;
    wire N__12208;
    wire N__12207;
    wire N__12206;
    wire N__12203;
    wire N__12202;
    wire N__12197;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12086;
    wire N__12085;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12053;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12033;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12021;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12009;
    wire N__12006;
    wire N__12005;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11966;
    wire N__11965;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11961;
    wire N__11960;
    wire N__11959;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11839;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11825;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11810;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11795;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11780;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11765;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11739;
    wire N__11736;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11683;
    wire N__11682;
    wire N__11679;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11658;
    wire N__11655;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11612;
    wire N__11607;
    wire N__11604;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11554;
    wire N__11553;
    wire N__11548;
    wire N__11545;
    wire N__11544;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11519;
    wire N__11514;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11463;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11403;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11375;
    wire N__11370;
    wire N__11367;
    wire N__11366;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11351;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11336;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11306;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11291;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11213;
    wire N__11212;
    wire N__11211;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11184;
    wire N__11177;
    wire N__11166;
    wire N__11165;
    wire N__11162;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11137;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11112;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11094;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11082;
    wire N__11081;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11051;
    wire N__11048;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11023;
    wire N__11018;
    wire N__11007;
    wire N__11004;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10986;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10975;
    wire N__10974;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10953;
    wire N__10946;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10922;
    wire N__10917;
    wire N__10908;
    wire N__10905;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10893;
    wire N__10890;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10793;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10693;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10661;
    wire N__10656;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10646;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10631;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10616;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10601;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10586;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10491;
    wire N__10482;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10474;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10439;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10420;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10266;
    wire N__10265;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10253;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10020;
    wire N__10017;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10002;
    wire N__10001;
    wire N__9998;
    wire N__9997;
    wire N__9994;
    wire N__9989;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9978;
    wire N__9971;
    wire N__9966;
    wire N__9965;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9949;
    wire N__9942;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9934;
    wire N__9929;
    wire N__9924;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9912;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9887;
    wire N__9882;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9843;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9819;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9804;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9768;
    wire N__9767;
    wire N__9764;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9747;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9737;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9533;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9515;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9446;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9428;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9410;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9284;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9272;
    wire N__9269;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire VCCG0;
    wire GNDG0;
    wire \uart_frame_decoder.WDTZ0Z_0 ;
    wire bfn_1_17_0_;
    wire \uart_frame_decoder.WDTZ0Z_1 ;
    wire \uart_frame_decoder.un1_WDT_cry_0 ;
    wire \uart_frame_decoder.WDTZ0Z_2 ;
    wire \uart_frame_decoder.un1_WDT_cry_1 ;
    wire \uart_frame_decoder.WDTZ0Z_3 ;
    wire \uart_frame_decoder.un1_WDT_cry_2 ;
    wire \uart_frame_decoder.un1_WDT_cry_3 ;
    wire \uart_frame_decoder.un1_WDT_cry_4 ;
    wire \uart_frame_decoder.un1_WDT_cry_5 ;
    wire \uart_frame_decoder.un1_WDT_cry_6 ;
    wire \uart_frame_decoder.un1_WDT_cry_7 ;
    wire bfn_1_18_0_;
    wire \uart_frame_decoder.un1_WDT_cry_8 ;
    wire \uart_frame_decoder.un1_WDT_cry_9 ;
    wire \uart_frame_decoder.un1_WDT_cry_10 ;
    wire \uart_frame_decoder.un1_WDT_cry_11 ;
    wire \uart_frame_decoder.un1_WDT_cry_12 ;
    wire \uart_frame_decoder.un1_WDT_cry_13 ;
    wire \uart_frame_decoder.un1_WDT_cry_14 ;
    wire bfn_1_19_0_;
    wire \uart_frame_decoder.count8_axb_1 ;
    wire \uart_frame_decoder.count8_cry_0 ;
    wire \uart_frame_decoder.count_i_2 ;
    wire \uart_frame_decoder.count8_cry_1 ;
    wire \uart_frame_decoder.count8 ;
    wire \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21 ;
    wire \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_ ;
    wire \uart_frame_decoder.count_RNIV5MSZ0Z_0 ;
    wire \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ;
    wire \uart_frame_decoder.count8_0_i ;
    wire bfn_1_23_0_;
    wire \scaler_3.un3_source_data_0_cry_0 ;
    wire frame_decoder_OFF3data_2;
    wire \scaler_3.un3_source_data_0_cry_1 ;
    wire frame_decoder_OFF3data_3;
    wire \scaler_3.un3_source_data_0_cry_2 ;
    wire frame_decoder_OFF3data_4;
    wire \scaler_3.un3_source_data_0_cry_3 ;
    wire frame_decoder_OFF3data_5;
    wire \scaler_3.un3_source_data_0_cry_4 ;
    wire frame_decoder_OFF3data_6;
    wire \scaler_3.un3_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_7 ;
    wire bfn_1_24_0_;
    wire \scaler_3.un3_source_data_0_cry_8 ;
    wire \scaler_3.N_795_i_l_ofxZ0 ;
    wire \scaler_3.un2_source_data_0_cry_1_c_RNO_1 ;
    wire bfn_1_25_0_;
    wire \scaler_3.un2_source_data_0_cry_1 ;
    wire \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ;
    wire \scaler_3.un2_source_data_0_cry_2 ;
    wire \scaler_3.un3_source_data_0_cry_2_c_RNIR08I ;
    wire \scaler_3.un2_source_data_0_cry_3 ;
    wire \scaler_3.un3_source_data_0_cry_3_c_RNIU49I ;
    wire \scaler_3.un2_source_data_0_cry_4 ;
    wire \scaler_3.un3_source_data_0_cry_4_c_RNI19AI ;
    wire \scaler_3.un2_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ;
    wire \scaler_3.un2_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ;
    wire \scaler_3.un2_source_data_0_cry_7 ;
    wire \scaler_3.un2_source_data_0_cry_8 ;
    wire \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ;
    wire \scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ;
    wire bfn_1_26_0_;
    wire \scaler_3.un2_source_data_0_cry_9 ;
    wire \uart_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire bfn_1_29_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_OFF4data_5;
    wire frame_decoder_CH4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire bfn_1_30_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire frame_decoder_OFF4data_7;
    wire \scaler_4.N_807_i_l_ofxZ0 ;
    wire \uart_frame_decoder.WDTZ0Z_8 ;
    wire \uart_frame_decoder.WDTZ0Z_11 ;
    wire \uart_frame_decoder.WDTZ0Z_10 ;
    wire \uart_frame_decoder.WDTZ0Z_13 ;
    wire \uart_frame_decoder.WDTZ0Z_12 ;
    wire \uart_frame_decoder.WDTZ0Z_9 ;
    wire \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ;
    wire \uart_frame_decoder.WDT8lto13_1 ;
    wire \uart_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \uart_frame_decoder.WDT8_0_i ;
    wire \uart_frame_decoder.WDTZ0Z_6 ;
    wire \uart_frame_decoder.WDTZ0Z_5 ;
    wire \uart_frame_decoder.WDTZ0Z_7 ;
    wire \uart_frame_decoder.WDTZ0Z_4 ;
    wire \uart_frame_decoder.WDT_RNIM6B11Z0Z_4 ;
    wire \uart_frame_decoder.WDTZ0Z_15 ;
    wire \uart_frame_decoder.WDTZ0Z_14 ;
    wire \uart_frame_decoder.WDT8lt14_0 ;
    wire \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_ ;
    wire \uart_frame_decoder.state_1Z0Z_3 ;
    wire \uart_frame_decoder.state_1Z0Z_2 ;
    wire \uart_frame_decoder.state_1Z0Z_4 ;
    wire \uart_frame_decoder.countZ0Z_2 ;
    wire \uart_frame_decoder.countZ0Z_1 ;
    wire \uart_frame_decoder.count8_0 ;
    wire \uart_frame_decoder.state_1_ns_i_i_0_0_cascade_ ;
    wire bfn_2_21_0_;
    wire frame_decoder_CH2data_1;
    wire frame_decoder_OFF2data_1;
    wire \scaler_2.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH2data_2;
    wire frame_decoder_OFF2data_2;
    wire \scaler_2.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH2data_3;
    wire frame_decoder_OFF2data_3;
    wire \scaler_2.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH2data_4;
    wire frame_decoder_OFF2data_4;
    wire \scaler_2.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH2data_5;
    wire frame_decoder_OFF2data_5;
    wire \scaler_2.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH2data_6;
    wire frame_decoder_OFF2data_6;
    wire \scaler_2.un3_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_7 ;
    wire bfn_2_22_0_;
    wire \scaler_2.un3_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_axb_7 ;
    wire \uart_frame_decoder.source_CH1data_1_sqmuxa ;
    wire \uart_frame_decoder.source_offset2data_1_sqmuxa_0 ;
    wire frame_decoder_CH2data_7;
    wire frame_decoder_OFF2data_7;
    wire \scaler_2.N_783_i_l_ofxZ0 ;
    wire \uart_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \uart_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire \uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire frame_decoder_OFF3data_7;
    wire \scaler_3.un3_source_data_0_axb_7 ;
    wire \uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ;
    wire frame_decoder_CH3data_1;
    wire frame_decoder_CH3data_2;
    wire frame_decoder_CH3data_3;
    wire frame_decoder_CH3data_4;
    wire frame_decoder_CH3data_5;
    wire frame_decoder_CH3data_6;
    wire frame_decoder_CH3data_7;
    wire bfn_2_27_0_;
    wire frame_decoder_CH1data_1;
    wire frame_decoder_OFF1data_1;
    wire \scaler_1.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH1data_2;
    wire frame_decoder_OFF1data_2;
    wire \scaler_1.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH1data_3;
    wire frame_decoder_OFF1data_3;
    wire \scaler_1.un3_source_data_0_cry_2 ;
    wire frame_decoder_OFF1data_4;
    wire \scaler_1.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH1data_5;
    wire frame_decoder_OFF1data_5;
    wire \scaler_1.un3_source_data_0_cry_4 ;
    wire frame_decoder_OFF1data_6;
    wire frame_decoder_CH1data_6;
    wire \scaler_1.un3_source_data_0_cry_5 ;
    wire \scaler_1.un3_source_data_0_cry_6 ;
    wire \scaler_1.un3_source_data_0_cry_7 ;
    wire bfn_2_28_0_;
    wire \scaler_1.un3_source_data_0_cry_8 ;
    wire \scaler_1.N_771_i_l_ofxZ0 ;
    wire frame_decoder_CH4data_0;
    wire frame_decoder_OFF4data_0;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNO_2 ;
    wire bfn_2_29_0_;
    wire \scaler_4.un2_source_data_0 ;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNI15MI ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNI49NI ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire bfn_2_30_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire \uart.CO1 ;
    wire \uart.N_133_0 ;
    wire \uart.N_177_cascade_ ;
    wire \uart.state_srsts_i_0_3 ;
    wire \uart.N_168_1_cascade_ ;
    wire \uart.N_154_0 ;
    wire \uart.data_Auxce_0_0_0 ;
    wire \uart.data_Auxce_0_1 ;
    wire \uart.data_Auxce_0_3 ;
    wire \uart.data_Auxce_0_5 ;
    wire \uart.data_Auxce_0_6 ;
    wire \uart.N_177 ;
    wire \uart.state_srsts_0_0_0_cascade_ ;
    wire \uart_frame_decoder.state_1_RNI592GZ0Z_10 ;
    wire \uart_frame_decoder.state_1_RNO_3Z0Z_0 ;
    wire \uart_frame_decoder.N_168_i_1 ;
    wire \uart_frame_decoder.state_1_RNO_2Z0Z_0 ;
    wire \uart_frame_decoder.state_1Z0Z_7 ;
    wire \uart_frame_decoder.state_1Z0Z_0 ;
    wire \uart_frame_decoder.N_79_4 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ;
    wire \uart.data_AuxZ1Z_0 ;
    wire uart_data_0;
    wire \uart_frame_decoder.state_1Z0Z_1 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_2 ;
    wire \uart.data_AuxZ0Z_5 ;
    wire uart_data_5;
    wire \uart.data_AuxZ1Z_2 ;
    wire uart_data_2;
    wire \uart.data_AuxZ0Z_7 ;
    wire \uart.data_AuxZ1Z_1 ;
    wire bfn_3_21_0_;
    wire \scaler_2.un2_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_1_c_RNILSPH ;
    wire \scaler_2.un2_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ;
    wire \scaler_2.un2_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ;
    wire \scaler_2.un2_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ;
    wire \scaler_2.un2_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ;
    wire \scaler_2.un2_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ;
    wire \scaler_2.un2_source_data_0_cry_7 ;
    wire \scaler_2.un2_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ;
    wire \scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ;
    wire bfn_3_22_0_;
    wire \scaler_2.un2_source_data_0_cry_9 ;
    wire \scaler_3.un2_source_data_0 ;
    wire \uart_frame_decoder.source_offset2data_1_sqmuxa ;
    wire \uart_frame_decoder.state_1Z0Z_8 ;
    wire \uart_frame_decoder.source_offset3data_1_sqmuxa ;
    wire \uart_frame_decoder.state_1Z0Z_9 ;
    wire \uart_frame_decoder.state_1Z0Z_5 ;
    wire \uart_frame_decoder.source_CH4data_1_sqmuxa ;
    wire uart_data_7;
    wire frame_decoder_CH4data_7;
    wire \uart_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire \uart_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \uart_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire frame_decoder_OFF1data_0;
    wire frame_decoder_CH1data_0;
    wire frame_decoder_OFF1data_7;
    wire frame_decoder_CH1data_7;
    wire \scaler_1.un3_source_data_0_axb_7 ;
    wire bfn_3_26_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire scaler_4_data_14;
    wire bfn_3_27_0_;
    wire \scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_3_28_0_;
    wire \scaler_1.un2_source_data_0 ;
    wire \scaler_1.un2_source_data_0_cry_1 ;
    wire \scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ;
    wire \scaler_1.un2_source_data_0_cry_2 ;
    wire \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ;
    wire \scaler_1.un2_source_data_0_cry_3 ;
    wire \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ;
    wire \scaler_1.un2_source_data_0_cry_4 ;
    wire \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ;
    wire \scaler_1.un2_source_data_0_cry_5 ;
    wire \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ;
    wire \scaler_1.un2_source_data_0_cry_6 ;
    wire \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ;
    wire \scaler_1.un2_source_data_0_cry_7 ;
    wire \scaler_1.un2_source_data_0_cry_8 ;
    wire \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ;
    wire \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ;
    wire bfn_3_29_0_;
    wire \scaler_1.un2_source_data_0_cry_9 ;
    wire frame_decoder_dv_c_0_g;
    wire frame_decoder_OFF3data_1;
    wire \uart_frame_decoder.source_offset3data_1_sqmuxa_0 ;
    wire \uart_sync.aux_2__0_Z0Z_0 ;
    wire \uart_sync.aux_3__0_Z0Z_0 ;
    wire \uart.N_151 ;
    wire \uart.stateZ0Z_2 ;
    wire \uart.N_159 ;
    wire \uart.timer_Count_0_sqmuxa_1_cascade_ ;
    wire \uart.N_180 ;
    wire \uart.N_180_cascade_ ;
    wire \uart.un1_state_5_0 ;
    wire \uart.N_143_0 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \uart.N_153_0_cascade_ ;
    wire \uart.state_srsts_i_a3_0_0_3_cascade_ ;
    wire \uart.N_170 ;
    wire \uart.un1_state_2_0_a3_2 ;
    wire \uart.N_146_0 ;
    wire \uart.un1_state_2_0 ;
    wire \reset_module_System.reset6_11_cascade_ ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \uart.data_Auxce_0_0_4 ;
    wire \reset_module_System.reset6_14 ;
    wire \uart.state_RNIAFHLZ0Z_3 ;
    wire \uart.N_153_0 ;
    wire \uart.stateZ0Z_3 ;
    wire \uart.N_168_1 ;
    wire \uart.N_167 ;
    wire \uart.stateZ0Z_4 ;
    wire \uart.bit_CountZ0Z_2 ;
    wire \uart.bit_CountZ0Z_1 ;
    wire \uart.bit_CountZ0Z_0 ;
    wire \uart.data_Auxce_0_0_2 ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.reset6_3 ;
    wire \reset_module_System.reset6_17 ;
    wire uart_data_1;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ;
    wire \uart.stateZ0Z_0 ;
    wire \uart.stateZ0Z_1 ;
    wire uart_input_sync;
    wire \uart.data_AuxZ0Z_3 ;
    wire uart_data_3;
    wire \uart.data_AuxZ0Z_6 ;
    wire uart_data_6;
    wire \uart_frame_decoder.state_1Z0Z_6 ;
    wire \uart_frame_decoder.source_offset1data_1_sqmuxa ;
    wire \uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_ ;
    wire \uart_frame_decoder.source_offset1data_1_sqmuxa_0 ;
    wire \uart.data_rdyc_1 ;
    wire \uart.data_AuxZ0Z_4 ;
    wire \uart.state_RNIQABT2Z0Z_4 ;
    wire \uart_frame_decoder.state_1_ns_0_i_o2_0_10 ;
    wire \uart_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \uart_frame_decoder.state_1Z0Z_10 ;
    wire uart_data_rdy;
    wire \uart_frame_decoder.count8_THRU_CO ;
    wire scaler_4_data_6;
    wire frame_decoder_OFF3data_0;
    wire frame_decoder_CH3data_0;
    wire bfn_4_24_0_;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire scaler_2_data_11;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire scaler_2_data_14;
    wire bfn_4_25_0_;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire scaler_4_data_10;
    wire scaler_2_data_10;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire scaler_3_data_6;
    wire bfn_4_27_0_;
    wire scaler_3_data_7;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire scaler_3_data_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire scaler_3_data_12;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire scaler_3_data_14;
    wire bfn_4_28_0_;
    wire scaler_1_data_6;
    wire bfn_4_29_0_;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire scaler_1_data_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire scaler_1_data_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire scaler_1_data_14;
    wire bfn_4_30_0_;
    wire \uart_sync.aux_1__0_Z0Z_0 ;
    wire \uart.timer_CountZ0Z_1 ;
    wire bfn_5_15_0_;
    wire \uart.timer_CountZ0Z_2 ;
    wire \uart.un4_timer_Count_1_cry_1 ;
    wire \uart.timer_CountZ0Z_3 ;
    wire \uart.un4_timer_Count_1_cry_2 ;
    wire \uart.un4_timer_Count_1_cry_3 ;
    wire \uart.timer_CountZ0Z_5 ;
    wire \uart.un4_timer_Count_1_cry_4 ;
    wire \uart.timer_CountZ0Z_6 ;
    wire \uart.un4_timer_Count_1_cry_5 ;
    wire \uart.un4_timer_Count_1_cry_6 ;
    wire \uart.timer_CountZ0Z_7 ;
    wire \uart.timer_Count_1_sqmuxa_i ;
    wire \uart.timer_CountZ0Z_0 ;
    wire \uart.timer_CountZ0Z_4 ;
    wire \uart.un1_state_2_0_a3_0 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire bfn_5_17_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_5_18_0_;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_5_19_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_15 ;
    wire scaler_3_data_4;
    wire \scaler_2.un2_source_data_0 ;
    wire \scaler_2.un2_source_data_0_cry_1_c_RNO_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire scaler_2_data_6;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_rn_0_6 ;
    wire \ppm_encoder_1.un2_throttle_0_6_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_sn_6 ;
    wire \ppm_encoder_1.N_415 ;
    wire \ppm_encoder_1.N_414_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.N_412 ;
    wire \ppm_encoder_1.N_411_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire scaler_2_data_9;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire scaler_4_data_9;
    wire scaler_3_data_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire frame_decoder_OFF2data_0;
    wire frame_decoder_CH2data_0;
    wire scaler_2_data_4;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire uart_data_4;
    wire frame_decoder_CH1data_4;
    wire \uart_frame_decoder.source_CH1data_1_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire scaler_1_data_12;
    wire scaler_1_data_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire frame_decoder_dv_c;
    wire frame_decoder_dv_c_0;
    wire uart_input_c;
    wire \uart_sync.aux_0__0_Z0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_o2_0_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_ ;
    wire \ppm_encoder_1.N_462 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_i_i_1_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ;
    wire bfn_7_23_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.init_pulses_RNI398E4Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire bfn_7_24_0_;
    wire \ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_7_25_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14 ;
    wire \ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15 ;
    wire \ppm_encoder_1.N_403 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.N_114_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.N_348_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.init_pulses_18_i_0_14_cascade_ ;
    wire \ppm_encoder_1.init_pulses_18_i_a2_0_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.N_241_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_ ;
    wire scaler_2_data_13;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13 ;
    wire scaler_3_data_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_11 ;
    wire scaler_3_data_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire scaler_1_data_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire scaler_2_data_12;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.N_418 ;
    wire \ppm_encoder_1.N_417_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_ ;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire scaler_2_data_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire scaler_1_data_8;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire scaler_3_data_8;
    wire scaler_3_data_5;
    wire scaler_4_data_4;
    wire scaler_1_data_4;
    wire scaler_1_data_5;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0 ;
    wire scaler_2_data_5;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire scaler_4_data_5;
    wire \ppm_encoder_1.scaler_1_dv_0 ;
    wire \ppm_encoder_1.N_252_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_8 ;
    wire \ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8 ;
    wire \ppm_encoder_1.N_235_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7 ;
    wire \ppm_encoder_1.N_114 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_12 ;
    wire \ppm_encoder_1.N_407_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_14 ;
    wire \ppm_encoder_1.N_251_i_i ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_i_o2_0_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.N_245_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.N_241 ;
    wire \ppm_encoder_1.N_348 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire scaler_1_data_7;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire scaler_4_data_7;
    wire \ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_0_0_7_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_rn_0_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire scaler_2_data_7;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1 ;
    wire \ppm_encoder_1.N_426 ;
    wire \ppm_encoder_1.N_246 ;
    wire \ppm_encoder_1.N_426_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3 ;
    wire scaler_1_dv;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.N_248_i_i ;
    wire \ppm_encoder_1.N_250_i_i ;
    wire \ppm_encoder_1.N_254_i_i ;
    wire \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.N_246_i_i ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.N_256_i_i ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.N_305 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_ ;
    wire \ppm_encoder_1.N_260_i_i ;
    wire \ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI83R42Z0Z_0 ;
    wire bfn_9_26_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2 ;
    wire \ppm_encoder_1.N_249_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6 ;
    wire \ppm_encoder_1.N_253_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire bfn_9_27_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.N_259_i_i ;
    wire \ppm_encoder_1.init_pulses_RNIKON03Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire bfn_9_28_0_;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.N_204_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.N_379_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_i_o2_0_7 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_8 ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.N_391 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.N_396 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.N_325 ;
    wire \ppm_encoder_1.N_327_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_i_o2_0_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.N_204 ;
    wire \ppm_encoder_1.N_255_i_i ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.N_258_i_i ;
    wire \ppm_encoder_1.N_257_i_i ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_6 ;
    wire \ppm_encoder_1.N_301 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.N_302 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_12 ;
    wire \ppm_encoder_1.N_393 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.PPM_STATE_fastZ0Z_0 ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.init_pulses_RNILB4MZ0Z_0 ;
    wire \ppm_encoder_1.N_247_i_i ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.N_441_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_18 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.N_383 ;
    wire \ppm_encoder_1.N_385_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.N_369 ;
    wire \ppm_encoder_1.N_371_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.N_360 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.N_365 ;
    wire \ppm_encoder_1.N_443 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_1 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire bfn_11_24_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_11_25_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_11_26_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_512_g ;
    wire \ppm_encoder_1.N_247 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_11 ;
    wire \ppm_encoder_1.N_388 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_13 ;
    wire \ppm_encoder_1.N_303 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ;
    wire \ppm_encoder_1.N_238_i_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.N_235 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ;
    wire \ppm_encoder_1.N_304 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.N_300 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_ ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ;
    wire \ppm_encoder_1.N_431_cascade_ ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_1_9 ;
    wire \ppm_encoder_1.N_441 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.N_244 ;
    wire \ppm_encoder_1.pulses2count_9_0_1_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire clk_system_c_g;
    wire \ppm_encoder_1.N_238_i_0_g ;
    wire reset_system_g;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_13_24_0_;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire bfn_13_25_0_;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire CONSTANT_ONE_NET;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.N_330 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire reset_system;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire _gnd_net_;

    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__24856),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__24858),
            .DIN(N__24857),
            .DOUT(N__24856),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__24858),
            .PADOUT(N__24857),
            .PADIN(N__24856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__24847),
            .DIN(N__24846),
            .DOUT(N__24845),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__24847),
            .PADOUT(N__24846),
            .PADIN(N__24845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam frame_decoder_dv_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD frame_decoder_dv_obuf_iopad (
            .OE(N__24838),
            .DIN(N__24837),
            .DOUT(N__24836),
            .PACKAGEPIN(frame_decoder_dv));
    defparam frame_decoder_dv_obuf_preio.NEG_TRIGGER=1'b0;
    defparam frame_decoder_dv_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO frame_decoder_dv_obuf_preio (
            .PADOEN(N__24838),
            .PADOUT(N__24837),
            .PADIN(N__24836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14955),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_ibuf_iopad (
            .OE(N__24829),
            .DIN(N__24828),
            .DOUT(N__24827),
            .PACKAGEPIN(uart_input));
    defparam uart_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_ibuf_preio (
            .PADOEN(N__24829),
            .PADOUT(N__24828),
            .PADIN(N__24827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_debug_obuf_iopad (
            .OE(N__24820),
            .DIN(N__24819),
            .DOUT(N__24818),
            .PACKAGEPIN(uart_input_debug));
    defparam uart_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_input_debug_obuf_preio (
            .PADOEN(N__24820),
            .PADOUT(N__24819),
            .PADIN(N__24818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15410),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5994 (
            .O(N__24801),
            .I(N__24798));
    LocalMux I__5993 (
            .O(N__24798),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__5992 (
            .O(N__24795),
            .I(N__24792));
    LocalMux I__5991 (
            .O(N__24792),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    CascadeMux I__5990 (
            .O(N__24789),
            .I(N__24786));
    InMux I__5989 (
            .O(N__24786),
            .I(N__24783));
    LocalMux I__5988 (
            .O(N__24783),
            .I(N__24780));
    Odrv4 I__5987 (
            .O(N__24780),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__5986 (
            .O(N__24777),
            .I(N__24774));
    LocalMux I__5985 (
            .O(N__24774),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    CascadeMux I__5984 (
            .O(N__24771),
            .I(N__24764));
    CascadeMux I__5983 (
            .O(N__24770),
            .I(N__24761));
    CascadeMux I__5982 (
            .O(N__24769),
            .I(N__24758));
    CascadeMux I__5981 (
            .O(N__24768),
            .I(N__24754));
    CascadeMux I__5980 (
            .O(N__24767),
            .I(N__24751));
    InMux I__5979 (
            .O(N__24764),
            .I(N__24738));
    InMux I__5978 (
            .O(N__24761),
            .I(N__24735));
    InMux I__5977 (
            .O(N__24758),
            .I(N__24732));
    CascadeMux I__5976 (
            .O(N__24757),
            .I(N__24729));
    InMux I__5975 (
            .O(N__24754),
            .I(N__24726));
    InMux I__5974 (
            .O(N__24751),
            .I(N__24723));
    CascadeMux I__5973 (
            .O(N__24750),
            .I(N__24720));
    CascadeMux I__5972 (
            .O(N__24749),
            .I(N__24717));
    CascadeMux I__5971 (
            .O(N__24748),
            .I(N__24713));
    CascadeMux I__5970 (
            .O(N__24747),
            .I(N__24709));
    CascadeMux I__5969 (
            .O(N__24746),
            .I(N__24706));
    CascadeMux I__5968 (
            .O(N__24745),
            .I(N__24703));
    CascadeMux I__5967 (
            .O(N__24744),
            .I(N__24700));
    CascadeMux I__5966 (
            .O(N__24743),
            .I(N__24697));
    CascadeMux I__5965 (
            .O(N__24742),
            .I(N__24694));
    CascadeMux I__5964 (
            .O(N__24741),
            .I(N__24691));
    LocalMux I__5963 (
            .O(N__24738),
            .I(N__24687));
    LocalMux I__5962 (
            .O(N__24735),
            .I(N__24682));
    LocalMux I__5961 (
            .O(N__24732),
            .I(N__24682));
    InMux I__5960 (
            .O(N__24729),
            .I(N__24679));
    LocalMux I__5959 (
            .O(N__24726),
            .I(N__24674));
    LocalMux I__5958 (
            .O(N__24723),
            .I(N__24674));
    InMux I__5957 (
            .O(N__24720),
            .I(N__24671));
    InMux I__5956 (
            .O(N__24717),
            .I(N__24668));
    InMux I__5955 (
            .O(N__24716),
            .I(N__24665));
    InMux I__5954 (
            .O(N__24713),
            .I(N__24660));
    InMux I__5953 (
            .O(N__24712),
            .I(N__24660));
    InMux I__5952 (
            .O(N__24709),
            .I(N__24651));
    InMux I__5951 (
            .O(N__24706),
            .I(N__24651));
    InMux I__5950 (
            .O(N__24703),
            .I(N__24651));
    InMux I__5949 (
            .O(N__24700),
            .I(N__24651));
    InMux I__5948 (
            .O(N__24697),
            .I(N__24644));
    InMux I__5947 (
            .O(N__24694),
            .I(N__24644));
    InMux I__5946 (
            .O(N__24691),
            .I(N__24644));
    CascadeMux I__5945 (
            .O(N__24690),
            .I(N__24641));
    Span4Mux_h I__5944 (
            .O(N__24687),
            .I(N__24634));
    Span4Mux_v I__5943 (
            .O(N__24682),
            .I(N__24634));
    LocalMux I__5942 (
            .O(N__24679),
            .I(N__24634));
    Span4Mux_v I__5941 (
            .O(N__24674),
            .I(N__24629));
    LocalMux I__5940 (
            .O(N__24671),
            .I(N__24629));
    LocalMux I__5939 (
            .O(N__24668),
            .I(N__24624));
    LocalMux I__5938 (
            .O(N__24665),
            .I(N__24624));
    LocalMux I__5937 (
            .O(N__24660),
            .I(N__24617));
    LocalMux I__5936 (
            .O(N__24651),
            .I(N__24617));
    LocalMux I__5935 (
            .O(N__24644),
            .I(N__24617));
    InMux I__5934 (
            .O(N__24641),
            .I(N__24614));
    Span4Mux_v I__5933 (
            .O(N__24634),
            .I(N__24611));
    Sp12to4 I__5932 (
            .O(N__24629),
            .I(N__24608));
    Span4Mux_v I__5931 (
            .O(N__24624),
            .I(N__24605));
    Sp12to4 I__5930 (
            .O(N__24617),
            .I(N__24602));
    LocalMux I__5929 (
            .O(N__24614),
            .I(N__24599));
    Span4Mux_h I__5928 (
            .O(N__24611),
            .I(N__24596));
    Span12Mux_s11_v I__5927 (
            .O(N__24608),
            .I(N__24587));
    Sp12to4 I__5926 (
            .O(N__24605),
            .I(N__24587));
    Span12Mux_s11_v I__5925 (
            .O(N__24602),
            .I(N__24587));
    Span12Mux_s2_h I__5924 (
            .O(N__24599),
            .I(N__24587));
    Odrv4 I__5923 (
            .O(N__24596),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5922 (
            .O(N__24587),
            .I(CONSTANT_ONE_NET));
    InMux I__5921 (
            .O(N__24582),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__5920 (
            .O(N__24579),
            .I(N__24570));
    InMux I__5919 (
            .O(N__24578),
            .I(N__24570));
    InMux I__5918 (
            .O(N__24577),
            .I(N__24570));
    LocalMux I__5917 (
            .O(N__24570),
            .I(N__24566));
    InMux I__5916 (
            .O(N__24569),
            .I(N__24563));
    Odrv4 I__5915 (
            .O(N__24566),
            .I(\ppm_encoder_1.N_330 ));
    LocalMux I__5914 (
            .O(N__24563),
            .I(\ppm_encoder_1.N_330 ));
    InMux I__5913 (
            .O(N__24558),
            .I(N__24555));
    LocalMux I__5912 (
            .O(N__24555),
            .I(N__24551));
    InMux I__5911 (
            .O(N__24554),
            .I(N__24547));
    Span12Mux_s5_v I__5910 (
            .O(N__24551),
            .I(N__24544));
    InMux I__5909 (
            .O(N__24550),
            .I(N__24541));
    LocalMux I__5908 (
            .O(N__24547),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv12 I__5907 (
            .O(N__24544),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__5906 (
            .O(N__24541),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    CascadeMux I__5905 (
            .O(N__24534),
            .I(N__24530));
    CascadeMux I__5904 (
            .O(N__24533),
            .I(N__24525));
    InMux I__5903 (
            .O(N__24530),
            .I(N__24517));
    InMux I__5902 (
            .O(N__24529),
            .I(N__24517));
    InMux I__5901 (
            .O(N__24528),
            .I(N__24517));
    InMux I__5900 (
            .O(N__24525),
            .I(N__24514));
    IoInMux I__5899 (
            .O(N__24524),
            .I(N__24511));
    LocalMux I__5898 (
            .O(N__24517),
            .I(N__24508));
    LocalMux I__5897 (
            .O(N__24514),
            .I(N__24504));
    LocalMux I__5896 (
            .O(N__24511),
            .I(N__24501));
    Span4Mux_h I__5895 (
            .O(N__24508),
            .I(N__24497));
    InMux I__5894 (
            .O(N__24507),
            .I(N__24494));
    Span4Mux_v I__5893 (
            .O(N__24504),
            .I(N__24491));
    IoSpan4Mux I__5892 (
            .O(N__24501),
            .I(N__24488));
    InMux I__5891 (
            .O(N__24500),
            .I(N__24483));
    Span4Mux_h I__5890 (
            .O(N__24497),
            .I(N__24480));
    LocalMux I__5889 (
            .O(N__24494),
            .I(N__24477));
    Span4Mux_h I__5888 (
            .O(N__24491),
            .I(N__24474));
    Span4Mux_s3_v I__5887 (
            .O(N__24488),
            .I(N__24471));
    InMux I__5886 (
            .O(N__24487),
            .I(N__24468));
    InMux I__5885 (
            .O(N__24486),
            .I(N__24464));
    LocalMux I__5884 (
            .O(N__24483),
            .I(N__24457));
    Span4Mux_v I__5883 (
            .O(N__24480),
            .I(N__24457));
    Span4Mux_h I__5882 (
            .O(N__24477),
            .I(N__24452));
    Span4Mux_h I__5881 (
            .O(N__24474),
            .I(N__24452));
    Span4Mux_v I__5880 (
            .O(N__24471),
            .I(N__24449));
    LocalMux I__5879 (
            .O(N__24468),
            .I(N__24446));
    InMux I__5878 (
            .O(N__24467),
            .I(N__24443));
    LocalMux I__5877 (
            .O(N__24464),
            .I(N__24440));
    InMux I__5876 (
            .O(N__24463),
            .I(N__24435));
    InMux I__5875 (
            .O(N__24462),
            .I(N__24435));
    Span4Mux_v I__5874 (
            .O(N__24457),
            .I(N__24432));
    Span4Mux_v I__5873 (
            .O(N__24452),
            .I(N__24429));
    Span4Mux_v I__5872 (
            .O(N__24449),
            .I(N__24426));
    Odrv12 I__5871 (
            .O(N__24446),
            .I(reset_system));
    LocalMux I__5870 (
            .O(N__24443),
            .I(reset_system));
    Odrv4 I__5869 (
            .O(N__24440),
            .I(reset_system));
    LocalMux I__5868 (
            .O(N__24435),
            .I(reset_system));
    Odrv4 I__5867 (
            .O(N__24432),
            .I(reset_system));
    Odrv4 I__5866 (
            .O(N__24429),
            .I(reset_system));
    Odrv4 I__5865 (
            .O(N__24426),
            .I(reset_system));
    InMux I__5864 (
            .O(N__24411),
            .I(N__24408));
    LocalMux I__5863 (
            .O(N__24408),
            .I(N__24402));
    InMux I__5862 (
            .O(N__24407),
            .I(N__24398));
    InMux I__5861 (
            .O(N__24406),
            .I(N__24395));
    CascadeMux I__5860 (
            .O(N__24405),
            .I(N__24390));
    Span4Mux_h I__5859 (
            .O(N__24402),
            .I(N__24387));
    InMux I__5858 (
            .O(N__24401),
            .I(N__24384));
    LocalMux I__5857 (
            .O(N__24398),
            .I(N__24379));
    LocalMux I__5856 (
            .O(N__24395),
            .I(N__24379));
    InMux I__5855 (
            .O(N__24394),
            .I(N__24374));
    InMux I__5854 (
            .O(N__24393),
            .I(N__24374));
    InMux I__5853 (
            .O(N__24390),
            .I(N__24371));
    Odrv4 I__5852 (
            .O(N__24387),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__5851 (
            .O(N__24384),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__5850 (
            .O(N__24379),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__5849 (
            .O(N__24374),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__5848 (
            .O(N__24371),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    IoInMux I__5847 (
            .O(N__24360),
            .I(N__24357));
    LocalMux I__5846 (
            .O(N__24357),
            .I(N__24354));
    Span12Mux_s5_v I__5845 (
            .O(N__24354),
            .I(N__24351));
    Odrv12 I__5844 (
            .O(N__24351),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__5843 (
            .O(N__24348),
            .I(N__24342));
    InMux I__5842 (
            .O(N__24347),
            .I(N__24339));
    InMux I__5841 (
            .O(N__24346),
            .I(N__24336));
    InMux I__5840 (
            .O(N__24345),
            .I(N__24333));
    LocalMux I__5839 (
            .O(N__24342),
            .I(N__24330));
    LocalMux I__5838 (
            .O(N__24339),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__5837 (
            .O(N__24336),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__5836 (
            .O(N__24333),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv12 I__5835 (
            .O(N__24330),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__5834 (
            .O(N__24321),
            .I(N__24318));
    LocalMux I__5833 (
            .O(N__24318),
            .I(N__24315));
    Odrv12 I__5832 (
            .O(N__24315),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__5831 (
            .O(N__24312),
            .I(N__24309));
    InMux I__5830 (
            .O(N__24309),
            .I(N__24306));
    LocalMux I__5829 (
            .O(N__24306),
            .I(N__24303));
    Odrv4 I__5828 (
            .O(N__24303),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__5827 (
            .O(N__24300),
            .I(N__24295));
    InMux I__5826 (
            .O(N__24299),
            .I(N__24292));
    InMux I__5825 (
            .O(N__24298),
            .I(N__24289));
    LocalMux I__5824 (
            .O(N__24295),
            .I(N__24286));
    LocalMux I__5823 (
            .O(N__24292),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__5822 (
            .O(N__24289),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__5821 (
            .O(N__24286),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__5820 (
            .O(N__24279),
            .I(N__24276));
    LocalMux I__5819 (
            .O(N__24276),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__5818 (
            .O(N__24273),
            .I(N__24270));
    LocalMux I__5817 (
            .O(N__24270),
            .I(N__24267));
    Span4Mux_v I__5816 (
            .O(N__24267),
            .I(N__24264));
    Odrv4 I__5815 (
            .O(N__24264),
            .I(\ppm_encoder_1.pulses2count_9_i_0_1_9 ));
    InMux I__5814 (
            .O(N__24261),
            .I(N__24250));
    InMux I__5813 (
            .O(N__24260),
            .I(N__24247));
    InMux I__5812 (
            .O(N__24259),
            .I(N__24240));
    InMux I__5811 (
            .O(N__24258),
            .I(N__24240));
    InMux I__5810 (
            .O(N__24257),
            .I(N__24240));
    InMux I__5809 (
            .O(N__24256),
            .I(N__24237));
    InMux I__5808 (
            .O(N__24255),
            .I(N__24232));
    InMux I__5807 (
            .O(N__24254),
            .I(N__24229));
    CascadeMux I__5806 (
            .O(N__24253),
            .I(N__24226));
    LocalMux I__5805 (
            .O(N__24250),
            .I(N__24222));
    LocalMux I__5804 (
            .O(N__24247),
            .I(N__24219));
    LocalMux I__5803 (
            .O(N__24240),
            .I(N__24216));
    LocalMux I__5802 (
            .O(N__24237),
            .I(N__24213));
    InMux I__5801 (
            .O(N__24236),
            .I(N__24208));
    InMux I__5800 (
            .O(N__24235),
            .I(N__24208));
    LocalMux I__5799 (
            .O(N__24232),
            .I(N__24203));
    LocalMux I__5798 (
            .O(N__24229),
            .I(N__24203));
    InMux I__5797 (
            .O(N__24226),
            .I(N__24200));
    InMux I__5796 (
            .O(N__24225),
            .I(N__24197));
    Span4Mux_v I__5795 (
            .O(N__24222),
            .I(N__24194));
    Span4Mux_v I__5794 (
            .O(N__24219),
            .I(N__24191));
    Span4Mux_h I__5793 (
            .O(N__24216),
            .I(N__24188));
    Span12Mux_v I__5792 (
            .O(N__24213),
            .I(N__24185));
    LocalMux I__5791 (
            .O(N__24208),
            .I(N__24178));
    Span4Mux_h I__5790 (
            .O(N__24203),
            .I(N__24178));
    LocalMux I__5789 (
            .O(N__24200),
            .I(N__24178));
    LocalMux I__5788 (
            .O(N__24197),
            .I(\ppm_encoder_1.N_441 ));
    Odrv4 I__5787 (
            .O(N__24194),
            .I(\ppm_encoder_1.N_441 ));
    Odrv4 I__5786 (
            .O(N__24191),
            .I(\ppm_encoder_1.N_441 ));
    Odrv4 I__5785 (
            .O(N__24188),
            .I(\ppm_encoder_1.N_441 ));
    Odrv12 I__5784 (
            .O(N__24185),
            .I(\ppm_encoder_1.N_441 ));
    Odrv4 I__5783 (
            .O(N__24178),
            .I(\ppm_encoder_1.N_441 ));
    CascadeMux I__5782 (
            .O(N__24165),
            .I(N__24162));
    InMux I__5781 (
            .O(N__24162),
            .I(N__24158));
    InMux I__5780 (
            .O(N__24161),
            .I(N__24154));
    LocalMux I__5779 (
            .O(N__24158),
            .I(N__24151));
    InMux I__5778 (
            .O(N__24157),
            .I(N__24148));
    LocalMux I__5777 (
            .O(N__24154),
            .I(N__24144));
    Span4Mux_h I__5776 (
            .O(N__24151),
            .I(N__24139));
    LocalMux I__5775 (
            .O(N__24148),
            .I(N__24139));
    InMux I__5774 (
            .O(N__24147),
            .I(N__24136));
    Span4Mux_v I__5773 (
            .O(N__24144),
            .I(N__24131));
    Span4Mux_v I__5772 (
            .O(N__24139),
            .I(N__24131));
    LocalMux I__5771 (
            .O(N__24136),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    Odrv4 I__5770 (
            .O(N__24131),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    CascadeMux I__5769 (
            .O(N__24126),
            .I(N__24122));
    CascadeMux I__5768 (
            .O(N__24125),
            .I(N__24119));
    InMux I__5767 (
            .O(N__24122),
            .I(N__24113));
    InMux I__5766 (
            .O(N__24119),
            .I(N__24108));
    InMux I__5765 (
            .O(N__24118),
            .I(N__24108));
    InMux I__5764 (
            .O(N__24117),
            .I(N__24103));
    InMux I__5763 (
            .O(N__24116),
            .I(N__24103));
    LocalMux I__5762 (
            .O(N__24113),
            .I(\ppm_encoder_1.N_244 ));
    LocalMux I__5761 (
            .O(N__24108),
            .I(\ppm_encoder_1.N_244 ));
    LocalMux I__5760 (
            .O(N__24103),
            .I(\ppm_encoder_1.N_244 ));
    InMux I__5759 (
            .O(N__24096),
            .I(N__24093));
    LocalMux I__5758 (
            .O(N__24093),
            .I(\ppm_encoder_1.pulses2count_9_0_1_0 ));
    CascadeMux I__5757 (
            .O(N__24090),
            .I(N__24082));
    CascadeMux I__5756 (
            .O(N__24089),
            .I(N__24079));
    CascadeMux I__5755 (
            .O(N__24088),
            .I(N__24074));
    CascadeMux I__5754 (
            .O(N__24087),
            .I(N__24070));
    CascadeMux I__5753 (
            .O(N__24086),
            .I(N__24063));
    CascadeMux I__5752 (
            .O(N__24085),
            .I(N__24060));
    InMux I__5751 (
            .O(N__24082),
            .I(N__24057));
    InMux I__5750 (
            .O(N__24079),
            .I(N__24053));
    InMux I__5749 (
            .O(N__24078),
            .I(N__24050));
    InMux I__5748 (
            .O(N__24077),
            .I(N__24041));
    InMux I__5747 (
            .O(N__24074),
            .I(N__24041));
    InMux I__5746 (
            .O(N__24073),
            .I(N__24041));
    InMux I__5745 (
            .O(N__24070),
            .I(N__24041));
    InMux I__5744 (
            .O(N__24069),
            .I(N__24032));
    InMux I__5743 (
            .O(N__24068),
            .I(N__24032));
    InMux I__5742 (
            .O(N__24067),
            .I(N__24032));
    InMux I__5741 (
            .O(N__24066),
            .I(N__24032));
    InMux I__5740 (
            .O(N__24063),
            .I(N__24029));
    InMux I__5739 (
            .O(N__24060),
            .I(N__24026));
    LocalMux I__5738 (
            .O(N__24057),
            .I(N__24021));
    InMux I__5737 (
            .O(N__24056),
            .I(N__24018));
    LocalMux I__5736 (
            .O(N__24053),
            .I(N__24014));
    LocalMux I__5735 (
            .O(N__24050),
            .I(N__24011));
    LocalMux I__5734 (
            .O(N__24041),
            .I(N__24006));
    LocalMux I__5733 (
            .O(N__24032),
            .I(N__24006));
    LocalMux I__5732 (
            .O(N__24029),
            .I(N__23999));
    LocalMux I__5731 (
            .O(N__24026),
            .I(N__23996));
    InMux I__5730 (
            .O(N__24025),
            .I(N__23991));
    InMux I__5729 (
            .O(N__24024),
            .I(N__23991));
    Span4Mux_v I__5728 (
            .O(N__24021),
            .I(N__23986));
    LocalMux I__5727 (
            .O(N__24018),
            .I(N__23986));
    InMux I__5726 (
            .O(N__24017),
            .I(N__23983));
    Span4Mux_h I__5725 (
            .O(N__24014),
            .I(N__23977));
    Span4Mux_v I__5724 (
            .O(N__24011),
            .I(N__23972));
    Span4Mux_v I__5723 (
            .O(N__24006),
            .I(N__23972));
    CascadeMux I__5722 (
            .O(N__24005),
            .I(N__23969));
    InMux I__5721 (
            .O(N__24004),
            .I(N__23966));
    CascadeMux I__5720 (
            .O(N__24003),
            .I(N__23963));
    CascadeMux I__5719 (
            .O(N__24002),
            .I(N__23956));
    Span4Mux_v I__5718 (
            .O(N__23999),
            .I(N__23947));
    Span4Mux_h I__5717 (
            .O(N__23996),
            .I(N__23947));
    LocalMux I__5716 (
            .O(N__23991),
            .I(N__23947));
    Span4Mux_h I__5715 (
            .O(N__23986),
            .I(N__23947));
    LocalMux I__5714 (
            .O(N__23983),
            .I(N__23944));
    InMux I__5713 (
            .O(N__23982),
            .I(N__23937));
    InMux I__5712 (
            .O(N__23981),
            .I(N__23937));
    InMux I__5711 (
            .O(N__23980),
            .I(N__23937));
    Span4Mux_v I__5710 (
            .O(N__23977),
            .I(N__23934));
    Span4Mux_h I__5709 (
            .O(N__23972),
            .I(N__23931));
    InMux I__5708 (
            .O(N__23969),
            .I(N__23928));
    LocalMux I__5707 (
            .O(N__23966),
            .I(N__23925));
    InMux I__5706 (
            .O(N__23963),
            .I(N__23920));
    InMux I__5705 (
            .O(N__23962),
            .I(N__23920));
    InMux I__5704 (
            .O(N__23961),
            .I(N__23911));
    InMux I__5703 (
            .O(N__23960),
            .I(N__23911));
    InMux I__5702 (
            .O(N__23959),
            .I(N__23911));
    InMux I__5701 (
            .O(N__23956),
            .I(N__23911));
    Span4Mux_v I__5700 (
            .O(N__23947),
            .I(N__23908));
    Odrv4 I__5699 (
            .O(N__23944),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5698 (
            .O(N__23937),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5697 (
            .O(N__23934),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5696 (
            .O(N__23931),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5695 (
            .O(N__23928),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__5694 (
            .O(N__23925),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5693 (
            .O(N__23920),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5692 (
            .O(N__23911),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5691 (
            .O(N__23908),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__5690 (
            .O(N__23889),
            .I(N__23886));
    LocalMux I__5689 (
            .O(N__23886),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    ClkMux I__5688 (
            .O(N__23883),
            .I(N__23577));
    ClkMux I__5687 (
            .O(N__23882),
            .I(N__23577));
    ClkMux I__5686 (
            .O(N__23881),
            .I(N__23577));
    ClkMux I__5685 (
            .O(N__23880),
            .I(N__23577));
    ClkMux I__5684 (
            .O(N__23879),
            .I(N__23577));
    ClkMux I__5683 (
            .O(N__23878),
            .I(N__23577));
    ClkMux I__5682 (
            .O(N__23877),
            .I(N__23577));
    ClkMux I__5681 (
            .O(N__23876),
            .I(N__23577));
    ClkMux I__5680 (
            .O(N__23875),
            .I(N__23577));
    ClkMux I__5679 (
            .O(N__23874),
            .I(N__23577));
    ClkMux I__5678 (
            .O(N__23873),
            .I(N__23577));
    ClkMux I__5677 (
            .O(N__23872),
            .I(N__23577));
    ClkMux I__5676 (
            .O(N__23871),
            .I(N__23577));
    ClkMux I__5675 (
            .O(N__23870),
            .I(N__23577));
    ClkMux I__5674 (
            .O(N__23869),
            .I(N__23577));
    ClkMux I__5673 (
            .O(N__23868),
            .I(N__23577));
    ClkMux I__5672 (
            .O(N__23867),
            .I(N__23577));
    ClkMux I__5671 (
            .O(N__23866),
            .I(N__23577));
    ClkMux I__5670 (
            .O(N__23865),
            .I(N__23577));
    ClkMux I__5669 (
            .O(N__23864),
            .I(N__23577));
    ClkMux I__5668 (
            .O(N__23863),
            .I(N__23577));
    ClkMux I__5667 (
            .O(N__23862),
            .I(N__23577));
    ClkMux I__5666 (
            .O(N__23861),
            .I(N__23577));
    ClkMux I__5665 (
            .O(N__23860),
            .I(N__23577));
    ClkMux I__5664 (
            .O(N__23859),
            .I(N__23577));
    ClkMux I__5663 (
            .O(N__23858),
            .I(N__23577));
    ClkMux I__5662 (
            .O(N__23857),
            .I(N__23577));
    ClkMux I__5661 (
            .O(N__23856),
            .I(N__23577));
    ClkMux I__5660 (
            .O(N__23855),
            .I(N__23577));
    ClkMux I__5659 (
            .O(N__23854),
            .I(N__23577));
    ClkMux I__5658 (
            .O(N__23853),
            .I(N__23577));
    ClkMux I__5657 (
            .O(N__23852),
            .I(N__23577));
    ClkMux I__5656 (
            .O(N__23851),
            .I(N__23577));
    ClkMux I__5655 (
            .O(N__23850),
            .I(N__23577));
    ClkMux I__5654 (
            .O(N__23849),
            .I(N__23577));
    ClkMux I__5653 (
            .O(N__23848),
            .I(N__23577));
    ClkMux I__5652 (
            .O(N__23847),
            .I(N__23577));
    ClkMux I__5651 (
            .O(N__23846),
            .I(N__23577));
    ClkMux I__5650 (
            .O(N__23845),
            .I(N__23577));
    ClkMux I__5649 (
            .O(N__23844),
            .I(N__23577));
    ClkMux I__5648 (
            .O(N__23843),
            .I(N__23577));
    ClkMux I__5647 (
            .O(N__23842),
            .I(N__23577));
    ClkMux I__5646 (
            .O(N__23841),
            .I(N__23577));
    ClkMux I__5645 (
            .O(N__23840),
            .I(N__23577));
    ClkMux I__5644 (
            .O(N__23839),
            .I(N__23577));
    ClkMux I__5643 (
            .O(N__23838),
            .I(N__23577));
    ClkMux I__5642 (
            .O(N__23837),
            .I(N__23577));
    ClkMux I__5641 (
            .O(N__23836),
            .I(N__23577));
    ClkMux I__5640 (
            .O(N__23835),
            .I(N__23577));
    ClkMux I__5639 (
            .O(N__23834),
            .I(N__23577));
    ClkMux I__5638 (
            .O(N__23833),
            .I(N__23577));
    ClkMux I__5637 (
            .O(N__23832),
            .I(N__23577));
    ClkMux I__5636 (
            .O(N__23831),
            .I(N__23577));
    ClkMux I__5635 (
            .O(N__23830),
            .I(N__23577));
    ClkMux I__5634 (
            .O(N__23829),
            .I(N__23577));
    ClkMux I__5633 (
            .O(N__23828),
            .I(N__23577));
    ClkMux I__5632 (
            .O(N__23827),
            .I(N__23577));
    ClkMux I__5631 (
            .O(N__23826),
            .I(N__23577));
    ClkMux I__5630 (
            .O(N__23825),
            .I(N__23577));
    ClkMux I__5629 (
            .O(N__23824),
            .I(N__23577));
    ClkMux I__5628 (
            .O(N__23823),
            .I(N__23577));
    ClkMux I__5627 (
            .O(N__23822),
            .I(N__23577));
    ClkMux I__5626 (
            .O(N__23821),
            .I(N__23577));
    ClkMux I__5625 (
            .O(N__23820),
            .I(N__23577));
    ClkMux I__5624 (
            .O(N__23819),
            .I(N__23577));
    ClkMux I__5623 (
            .O(N__23818),
            .I(N__23577));
    ClkMux I__5622 (
            .O(N__23817),
            .I(N__23577));
    ClkMux I__5621 (
            .O(N__23816),
            .I(N__23577));
    ClkMux I__5620 (
            .O(N__23815),
            .I(N__23577));
    ClkMux I__5619 (
            .O(N__23814),
            .I(N__23577));
    ClkMux I__5618 (
            .O(N__23813),
            .I(N__23577));
    ClkMux I__5617 (
            .O(N__23812),
            .I(N__23577));
    ClkMux I__5616 (
            .O(N__23811),
            .I(N__23577));
    ClkMux I__5615 (
            .O(N__23810),
            .I(N__23577));
    ClkMux I__5614 (
            .O(N__23809),
            .I(N__23577));
    ClkMux I__5613 (
            .O(N__23808),
            .I(N__23577));
    ClkMux I__5612 (
            .O(N__23807),
            .I(N__23577));
    ClkMux I__5611 (
            .O(N__23806),
            .I(N__23577));
    ClkMux I__5610 (
            .O(N__23805),
            .I(N__23577));
    ClkMux I__5609 (
            .O(N__23804),
            .I(N__23577));
    ClkMux I__5608 (
            .O(N__23803),
            .I(N__23577));
    ClkMux I__5607 (
            .O(N__23802),
            .I(N__23577));
    ClkMux I__5606 (
            .O(N__23801),
            .I(N__23577));
    ClkMux I__5605 (
            .O(N__23800),
            .I(N__23577));
    ClkMux I__5604 (
            .O(N__23799),
            .I(N__23577));
    ClkMux I__5603 (
            .O(N__23798),
            .I(N__23577));
    ClkMux I__5602 (
            .O(N__23797),
            .I(N__23577));
    ClkMux I__5601 (
            .O(N__23796),
            .I(N__23577));
    ClkMux I__5600 (
            .O(N__23795),
            .I(N__23577));
    ClkMux I__5599 (
            .O(N__23794),
            .I(N__23577));
    ClkMux I__5598 (
            .O(N__23793),
            .I(N__23577));
    ClkMux I__5597 (
            .O(N__23792),
            .I(N__23577));
    ClkMux I__5596 (
            .O(N__23791),
            .I(N__23577));
    ClkMux I__5595 (
            .O(N__23790),
            .I(N__23577));
    ClkMux I__5594 (
            .O(N__23789),
            .I(N__23577));
    ClkMux I__5593 (
            .O(N__23788),
            .I(N__23577));
    ClkMux I__5592 (
            .O(N__23787),
            .I(N__23577));
    ClkMux I__5591 (
            .O(N__23786),
            .I(N__23577));
    ClkMux I__5590 (
            .O(N__23785),
            .I(N__23577));
    ClkMux I__5589 (
            .O(N__23784),
            .I(N__23577));
    ClkMux I__5588 (
            .O(N__23783),
            .I(N__23577));
    ClkMux I__5587 (
            .O(N__23782),
            .I(N__23577));
    GlobalMux I__5586 (
            .O(N__23577),
            .I(N__23574));
    gio2CtrlBuf I__5585 (
            .O(N__23574),
            .I(clk_system_c_g));
    CEMux I__5584 (
            .O(N__23571),
            .I(N__23541));
    CEMux I__5583 (
            .O(N__23570),
            .I(N__23541));
    CEMux I__5582 (
            .O(N__23569),
            .I(N__23541));
    CEMux I__5581 (
            .O(N__23568),
            .I(N__23541));
    CEMux I__5580 (
            .O(N__23567),
            .I(N__23541));
    CEMux I__5579 (
            .O(N__23566),
            .I(N__23541));
    CEMux I__5578 (
            .O(N__23565),
            .I(N__23541));
    CEMux I__5577 (
            .O(N__23564),
            .I(N__23541));
    CEMux I__5576 (
            .O(N__23563),
            .I(N__23541));
    CEMux I__5575 (
            .O(N__23562),
            .I(N__23541));
    GlobalMux I__5574 (
            .O(N__23541),
            .I(N__23538));
    gio2CtrlBuf I__5573 (
            .O(N__23538),
            .I(\ppm_encoder_1.N_238_i_0_g ));
    CascadeMux I__5572 (
            .O(N__23535),
            .I(N__23527));
    CascadeMux I__5571 (
            .O(N__23534),
            .I(N__23524));
    CascadeMux I__5570 (
            .O(N__23533),
            .I(N__23517));
    CascadeMux I__5569 (
            .O(N__23532),
            .I(N__23514));
    CascadeMux I__5568 (
            .O(N__23531),
            .I(N__23508));
    InMux I__5567 (
            .O(N__23530),
            .I(N__23487));
    InMux I__5566 (
            .O(N__23527),
            .I(N__23482));
    InMux I__5565 (
            .O(N__23524),
            .I(N__23482));
    InMux I__5564 (
            .O(N__23523),
            .I(N__23479));
    InMux I__5563 (
            .O(N__23522),
            .I(N__23476));
    InMux I__5562 (
            .O(N__23521),
            .I(N__23473));
    InMux I__5561 (
            .O(N__23520),
            .I(N__23470));
    InMux I__5560 (
            .O(N__23517),
            .I(N__23463));
    InMux I__5559 (
            .O(N__23514),
            .I(N__23463));
    InMux I__5558 (
            .O(N__23513),
            .I(N__23463));
    InMux I__5557 (
            .O(N__23512),
            .I(N__23460));
    InMux I__5556 (
            .O(N__23511),
            .I(N__23457));
    InMux I__5555 (
            .O(N__23508),
            .I(N__23450));
    InMux I__5554 (
            .O(N__23507),
            .I(N__23450));
    InMux I__5553 (
            .O(N__23506),
            .I(N__23450));
    InMux I__5552 (
            .O(N__23505),
            .I(N__23445));
    InMux I__5551 (
            .O(N__23504),
            .I(N__23445));
    InMux I__5550 (
            .O(N__23503),
            .I(N__23442));
    InMux I__5549 (
            .O(N__23502),
            .I(N__23439));
    InMux I__5548 (
            .O(N__23501),
            .I(N__23436));
    InMux I__5547 (
            .O(N__23500),
            .I(N__23433));
    InMux I__5546 (
            .O(N__23499),
            .I(N__23428));
    InMux I__5545 (
            .O(N__23498),
            .I(N__23428));
    InMux I__5544 (
            .O(N__23497),
            .I(N__23425));
    InMux I__5543 (
            .O(N__23496),
            .I(N__23422));
    InMux I__5542 (
            .O(N__23495),
            .I(N__23415));
    InMux I__5541 (
            .O(N__23494),
            .I(N__23415));
    InMux I__5540 (
            .O(N__23493),
            .I(N__23415));
    InMux I__5539 (
            .O(N__23492),
            .I(N__23412));
    InMux I__5538 (
            .O(N__23491),
            .I(N__23409));
    InMux I__5537 (
            .O(N__23490),
            .I(N__23406));
    LocalMux I__5536 (
            .O(N__23487),
            .I(N__23338));
    LocalMux I__5535 (
            .O(N__23482),
            .I(N__23335));
    LocalMux I__5534 (
            .O(N__23479),
            .I(N__23332));
    LocalMux I__5533 (
            .O(N__23476),
            .I(N__23329));
    LocalMux I__5532 (
            .O(N__23473),
            .I(N__23326));
    LocalMux I__5531 (
            .O(N__23470),
            .I(N__23323));
    LocalMux I__5530 (
            .O(N__23463),
            .I(N__23320));
    LocalMux I__5529 (
            .O(N__23460),
            .I(N__23317));
    LocalMux I__5528 (
            .O(N__23457),
            .I(N__23314));
    LocalMux I__5527 (
            .O(N__23450),
            .I(N__23311));
    LocalMux I__5526 (
            .O(N__23445),
            .I(N__23308));
    LocalMux I__5525 (
            .O(N__23442),
            .I(N__23305));
    LocalMux I__5524 (
            .O(N__23439),
            .I(N__23302));
    LocalMux I__5523 (
            .O(N__23436),
            .I(N__23299));
    LocalMux I__5522 (
            .O(N__23433),
            .I(N__23296));
    LocalMux I__5521 (
            .O(N__23428),
            .I(N__23293));
    LocalMux I__5520 (
            .O(N__23425),
            .I(N__23290));
    LocalMux I__5519 (
            .O(N__23422),
            .I(N__23287));
    LocalMux I__5518 (
            .O(N__23415),
            .I(N__23284));
    LocalMux I__5517 (
            .O(N__23412),
            .I(N__23281));
    LocalMux I__5516 (
            .O(N__23409),
            .I(N__23278));
    LocalMux I__5515 (
            .O(N__23406),
            .I(N__23275));
    SRMux I__5514 (
            .O(N__23405),
            .I(N__23100));
    SRMux I__5513 (
            .O(N__23404),
            .I(N__23100));
    SRMux I__5512 (
            .O(N__23403),
            .I(N__23100));
    SRMux I__5511 (
            .O(N__23402),
            .I(N__23100));
    SRMux I__5510 (
            .O(N__23401),
            .I(N__23100));
    SRMux I__5509 (
            .O(N__23400),
            .I(N__23100));
    SRMux I__5508 (
            .O(N__23399),
            .I(N__23100));
    SRMux I__5507 (
            .O(N__23398),
            .I(N__23100));
    SRMux I__5506 (
            .O(N__23397),
            .I(N__23100));
    SRMux I__5505 (
            .O(N__23396),
            .I(N__23100));
    SRMux I__5504 (
            .O(N__23395),
            .I(N__23100));
    SRMux I__5503 (
            .O(N__23394),
            .I(N__23100));
    SRMux I__5502 (
            .O(N__23393),
            .I(N__23100));
    SRMux I__5501 (
            .O(N__23392),
            .I(N__23100));
    SRMux I__5500 (
            .O(N__23391),
            .I(N__23100));
    SRMux I__5499 (
            .O(N__23390),
            .I(N__23100));
    SRMux I__5498 (
            .O(N__23389),
            .I(N__23100));
    SRMux I__5497 (
            .O(N__23388),
            .I(N__23100));
    SRMux I__5496 (
            .O(N__23387),
            .I(N__23100));
    SRMux I__5495 (
            .O(N__23386),
            .I(N__23100));
    SRMux I__5494 (
            .O(N__23385),
            .I(N__23100));
    SRMux I__5493 (
            .O(N__23384),
            .I(N__23100));
    SRMux I__5492 (
            .O(N__23383),
            .I(N__23100));
    SRMux I__5491 (
            .O(N__23382),
            .I(N__23100));
    SRMux I__5490 (
            .O(N__23381),
            .I(N__23100));
    SRMux I__5489 (
            .O(N__23380),
            .I(N__23100));
    SRMux I__5488 (
            .O(N__23379),
            .I(N__23100));
    SRMux I__5487 (
            .O(N__23378),
            .I(N__23100));
    SRMux I__5486 (
            .O(N__23377),
            .I(N__23100));
    SRMux I__5485 (
            .O(N__23376),
            .I(N__23100));
    SRMux I__5484 (
            .O(N__23375),
            .I(N__23100));
    SRMux I__5483 (
            .O(N__23374),
            .I(N__23100));
    SRMux I__5482 (
            .O(N__23373),
            .I(N__23100));
    SRMux I__5481 (
            .O(N__23372),
            .I(N__23100));
    SRMux I__5480 (
            .O(N__23371),
            .I(N__23100));
    SRMux I__5479 (
            .O(N__23370),
            .I(N__23100));
    SRMux I__5478 (
            .O(N__23369),
            .I(N__23100));
    SRMux I__5477 (
            .O(N__23368),
            .I(N__23100));
    SRMux I__5476 (
            .O(N__23367),
            .I(N__23100));
    SRMux I__5475 (
            .O(N__23366),
            .I(N__23100));
    SRMux I__5474 (
            .O(N__23365),
            .I(N__23100));
    SRMux I__5473 (
            .O(N__23364),
            .I(N__23100));
    SRMux I__5472 (
            .O(N__23363),
            .I(N__23100));
    SRMux I__5471 (
            .O(N__23362),
            .I(N__23100));
    SRMux I__5470 (
            .O(N__23361),
            .I(N__23100));
    SRMux I__5469 (
            .O(N__23360),
            .I(N__23100));
    SRMux I__5468 (
            .O(N__23359),
            .I(N__23100));
    SRMux I__5467 (
            .O(N__23358),
            .I(N__23100));
    SRMux I__5466 (
            .O(N__23357),
            .I(N__23100));
    SRMux I__5465 (
            .O(N__23356),
            .I(N__23100));
    SRMux I__5464 (
            .O(N__23355),
            .I(N__23100));
    SRMux I__5463 (
            .O(N__23354),
            .I(N__23100));
    SRMux I__5462 (
            .O(N__23353),
            .I(N__23100));
    SRMux I__5461 (
            .O(N__23352),
            .I(N__23100));
    SRMux I__5460 (
            .O(N__23351),
            .I(N__23100));
    SRMux I__5459 (
            .O(N__23350),
            .I(N__23100));
    SRMux I__5458 (
            .O(N__23349),
            .I(N__23100));
    SRMux I__5457 (
            .O(N__23348),
            .I(N__23100));
    SRMux I__5456 (
            .O(N__23347),
            .I(N__23100));
    SRMux I__5455 (
            .O(N__23346),
            .I(N__23100));
    SRMux I__5454 (
            .O(N__23345),
            .I(N__23100));
    SRMux I__5453 (
            .O(N__23344),
            .I(N__23100));
    SRMux I__5452 (
            .O(N__23343),
            .I(N__23100));
    SRMux I__5451 (
            .O(N__23342),
            .I(N__23100));
    SRMux I__5450 (
            .O(N__23341),
            .I(N__23100));
    Glb2LocalMux I__5449 (
            .O(N__23338),
            .I(N__23100));
    Glb2LocalMux I__5448 (
            .O(N__23335),
            .I(N__23100));
    Glb2LocalMux I__5447 (
            .O(N__23332),
            .I(N__23100));
    Glb2LocalMux I__5446 (
            .O(N__23329),
            .I(N__23100));
    Glb2LocalMux I__5445 (
            .O(N__23326),
            .I(N__23100));
    Glb2LocalMux I__5444 (
            .O(N__23323),
            .I(N__23100));
    Glb2LocalMux I__5443 (
            .O(N__23320),
            .I(N__23100));
    Glb2LocalMux I__5442 (
            .O(N__23317),
            .I(N__23100));
    Glb2LocalMux I__5441 (
            .O(N__23314),
            .I(N__23100));
    Glb2LocalMux I__5440 (
            .O(N__23311),
            .I(N__23100));
    Glb2LocalMux I__5439 (
            .O(N__23308),
            .I(N__23100));
    Glb2LocalMux I__5438 (
            .O(N__23305),
            .I(N__23100));
    Glb2LocalMux I__5437 (
            .O(N__23302),
            .I(N__23100));
    Glb2LocalMux I__5436 (
            .O(N__23299),
            .I(N__23100));
    Glb2LocalMux I__5435 (
            .O(N__23296),
            .I(N__23100));
    Glb2LocalMux I__5434 (
            .O(N__23293),
            .I(N__23100));
    Glb2LocalMux I__5433 (
            .O(N__23290),
            .I(N__23100));
    Glb2LocalMux I__5432 (
            .O(N__23287),
            .I(N__23100));
    Glb2LocalMux I__5431 (
            .O(N__23284),
            .I(N__23100));
    Glb2LocalMux I__5430 (
            .O(N__23281),
            .I(N__23100));
    Glb2LocalMux I__5429 (
            .O(N__23278),
            .I(N__23100));
    Glb2LocalMux I__5428 (
            .O(N__23275),
            .I(N__23100));
    GlobalMux I__5427 (
            .O(N__23100),
            .I(N__23097));
    gio2CtrlBuf I__5426 (
            .O(N__23097),
            .I(reset_system_g));
    InMux I__5425 (
            .O(N__23094),
            .I(N__23091));
    LocalMux I__5424 (
            .O(N__23091),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__5423 (
            .O(N__23088),
            .I(N__23085));
    LocalMux I__5422 (
            .O(N__23085),
            .I(N__23082));
    Span4Mux_h I__5421 (
            .O(N__23082),
            .I(N__23079));
    Odrv4 I__5420 (
            .O(N__23079),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__5419 (
            .O(N__23076),
            .I(N__23073));
    LocalMux I__5418 (
            .O(N__23073),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__5417 (
            .O(N__23070),
            .I(N__23067));
    LocalMux I__5416 (
            .O(N__23067),
            .I(N__23064));
    Odrv4 I__5415 (
            .O(N__23064),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__5414 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__5413 (
            .O(N__23058),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__5412 (
            .O(N__23055),
            .I(N__23052));
    LocalMux I__5411 (
            .O(N__23052),
            .I(N__23049));
    Odrv4 I__5410 (
            .O(N__23049),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1 ));
    CascadeMux I__5409 (
            .O(N__23046),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_ ));
    InMux I__5408 (
            .O(N__23043),
            .I(N__23040));
    LocalMux I__5407 (
            .O(N__23040),
            .I(N__23037));
    Span4Mux_v I__5406 (
            .O(N__23037),
            .I(N__23034));
    Odrv4 I__5405 (
            .O(N__23034),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    CascadeMux I__5404 (
            .O(N__23031),
            .I(N__23028));
    InMux I__5403 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__5402 (
            .O(N__23025),
            .I(N__23022));
    Odrv4 I__5401 (
            .O(N__23022),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__5400 (
            .O(N__23019),
            .I(N__23014));
    InMux I__5399 (
            .O(N__23018),
            .I(N__23009));
    InMux I__5398 (
            .O(N__23017),
            .I(N__23009));
    LocalMux I__5397 (
            .O(N__23014),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__5396 (
            .O(N__23009),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__5395 (
            .O(N__23004),
            .I(N__23001));
    LocalMux I__5394 (
            .O(N__23001),
            .I(N__22998));
    Odrv4 I__5393 (
            .O(N__22998),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__5392 (
            .O(N__22995),
            .I(N__22991));
    InMux I__5391 (
            .O(N__22994),
            .I(N__22987));
    LocalMux I__5390 (
            .O(N__22991),
            .I(N__22984));
    InMux I__5389 (
            .O(N__22990),
            .I(N__22981));
    LocalMux I__5388 (
            .O(N__22987),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv4 I__5387 (
            .O(N__22984),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__5386 (
            .O(N__22981),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__5385 (
            .O(N__22974),
            .I(N__22971));
    LocalMux I__5384 (
            .O(N__22971),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3 ));
    InMux I__5383 (
            .O(N__22968),
            .I(N__22963));
    InMux I__5382 (
            .O(N__22967),
            .I(N__22960));
    InMux I__5381 (
            .O(N__22966),
            .I(N__22957));
    LocalMux I__5380 (
            .O(N__22963),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__5379 (
            .O(N__22960),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__5378 (
            .O(N__22957),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    CascadeMux I__5377 (
            .O(N__22950),
            .I(N__22947));
    InMux I__5376 (
            .O(N__22947),
            .I(N__22944));
    LocalMux I__5375 (
            .O(N__22944),
            .I(N__22941));
    Odrv4 I__5374 (
            .O(N__22941),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4 ));
    InMux I__5373 (
            .O(N__22938),
            .I(N__22933));
    InMux I__5372 (
            .O(N__22937),
            .I(N__22930));
    InMux I__5371 (
            .O(N__22936),
            .I(N__22927));
    LocalMux I__5370 (
            .O(N__22933),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__5369 (
            .O(N__22930),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__5368 (
            .O(N__22927),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__5367 (
            .O(N__22920),
            .I(N__22917));
    LocalMux I__5366 (
            .O(N__22917),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2 ));
    InMux I__5365 (
            .O(N__22914),
            .I(N__22911));
    LocalMux I__5364 (
            .O(N__22911),
            .I(N__22908));
    Odrv4 I__5363 (
            .O(N__22908),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1 ));
    InMux I__5362 (
            .O(N__22905),
            .I(N__22902));
    LocalMux I__5361 (
            .O(N__22902),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4 ));
    CascadeMux I__5360 (
            .O(N__22899),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_ ));
    InMux I__5359 (
            .O(N__22896),
            .I(N__22892));
    InMux I__5358 (
            .O(N__22895),
            .I(N__22889));
    LocalMux I__5357 (
            .O(N__22892),
            .I(N__22886));
    LocalMux I__5356 (
            .O(N__22889),
            .I(N__22883));
    Span4Mux_v I__5355 (
            .O(N__22886),
            .I(N__22880));
    Span4Mux_h I__5354 (
            .O(N__22883),
            .I(N__22877));
    Odrv4 I__5353 (
            .O(N__22880),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5 ));
    Odrv4 I__5352 (
            .O(N__22877),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5 ));
    CascadeMux I__5351 (
            .O(N__22872),
            .I(N__22869));
    InMux I__5350 (
            .O(N__22869),
            .I(N__22863));
    InMux I__5349 (
            .O(N__22868),
            .I(N__22863));
    LocalMux I__5348 (
            .O(N__22863),
            .I(N__22859));
    InMux I__5347 (
            .O(N__22862),
            .I(N__22856));
    Odrv12 I__5346 (
            .O(N__22859),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ));
    LocalMux I__5345 (
            .O(N__22856),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ));
    CascadeMux I__5344 (
            .O(N__22851),
            .I(\ppm_encoder_1.N_431_cascade_ ));
    InMux I__5343 (
            .O(N__22848),
            .I(N__22845));
    LocalMux I__5342 (
            .O(N__22845),
            .I(N__22842));
    Span4Mux_h I__5341 (
            .O(N__22842),
            .I(N__22832));
    InMux I__5340 (
            .O(N__22841),
            .I(N__22825));
    InMux I__5339 (
            .O(N__22840),
            .I(N__22825));
    InMux I__5338 (
            .O(N__22839),
            .I(N__22825));
    InMux I__5337 (
            .O(N__22838),
            .I(N__22822));
    InMux I__5336 (
            .O(N__22837),
            .I(N__22819));
    InMux I__5335 (
            .O(N__22836),
            .I(N__22814));
    InMux I__5334 (
            .O(N__22835),
            .I(N__22814));
    Odrv4 I__5333 (
            .O(N__22832),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__5332 (
            .O(N__22825),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__5331 (
            .O(N__22822),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__5330 (
            .O(N__22819),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__5329 (
            .O(N__22814),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    IoInMux I__5328 (
            .O(N__22803),
            .I(N__22800));
    LocalMux I__5327 (
            .O(N__22800),
            .I(N__22797));
    IoSpan4Mux I__5326 (
            .O(N__22797),
            .I(N__22794));
    Span4Mux_s3_v I__5325 (
            .O(N__22794),
            .I(N__22791));
    Sp12to4 I__5324 (
            .O(N__22791),
            .I(N__22788));
    Span12Mux_v I__5323 (
            .O(N__22788),
            .I(N__22784));
    InMux I__5322 (
            .O(N__22787),
            .I(N__22781));
    Odrv12 I__5321 (
            .O(N__22784),
            .I(ppm_output_c));
    LocalMux I__5320 (
            .O(N__22781),
            .I(ppm_output_c));
    InMux I__5319 (
            .O(N__22776),
            .I(N__22773));
    LocalMux I__5318 (
            .O(N__22773),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    CascadeMux I__5317 (
            .O(N__22770),
            .I(N__22767));
    InMux I__5316 (
            .O(N__22767),
            .I(N__22763));
    InMux I__5315 (
            .O(N__22766),
            .I(N__22759));
    LocalMux I__5314 (
            .O(N__22763),
            .I(N__22756));
    InMux I__5313 (
            .O(N__22762),
            .I(N__22753));
    LocalMux I__5312 (
            .O(N__22759),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__5311 (
            .O(N__22756),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__5310 (
            .O(N__22753),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    CascadeMux I__5309 (
            .O(N__22746),
            .I(N__22743));
    InMux I__5308 (
            .O(N__22743),
            .I(N__22740));
    LocalMux I__5307 (
            .O(N__22740),
            .I(N__22737));
    Odrv12 I__5306 (
            .O(N__22737),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__5305 (
            .O(N__22734),
            .I(N__22729));
    InMux I__5304 (
            .O(N__22733),
            .I(N__22726));
    InMux I__5303 (
            .O(N__22732),
            .I(N__22723));
    LocalMux I__5302 (
            .O(N__22729),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__5301 (
            .O(N__22726),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__5300 (
            .O(N__22723),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__5299 (
            .O(N__22716),
            .I(N__22713));
    LocalMux I__5298 (
            .O(N__22713),
            .I(N__22710));
    Span4Mux_h I__5297 (
            .O(N__22710),
            .I(N__22707));
    Odrv4 I__5296 (
            .O(N__22707),
            .I(\ppm_encoder_1.pulses2count_9_i_1_8 ));
    InMux I__5295 (
            .O(N__22704),
            .I(N__22699));
    CascadeMux I__5294 (
            .O(N__22703),
            .I(N__22696));
    CascadeMux I__5293 (
            .O(N__22702),
            .I(N__22693));
    LocalMux I__5292 (
            .O(N__22699),
            .I(N__22689));
    InMux I__5291 (
            .O(N__22696),
            .I(N__22684));
    InMux I__5290 (
            .O(N__22693),
            .I(N__22684));
    InMux I__5289 (
            .O(N__22692),
            .I(N__22681));
    Span4Mux_v I__5288 (
            .O(N__22689),
            .I(N__22676));
    LocalMux I__5287 (
            .O(N__22684),
            .I(N__22676));
    LocalMux I__5286 (
            .O(N__22681),
            .I(N__22673));
    Span4Mux_h I__5285 (
            .O(N__22676),
            .I(N__22670));
    Span4Mux_v I__5284 (
            .O(N__22673),
            .I(N__22667));
    Span4Mux_v I__5283 (
            .O(N__22670),
            .I(N__22664));
    Span4Mux_v I__5282 (
            .O(N__22667),
            .I(N__22661));
    Odrv4 I__5281 (
            .O(N__22664),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    Odrv4 I__5280 (
            .O(N__22661),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__5279 (
            .O(N__22656),
            .I(N__22653));
    LocalMux I__5278 (
            .O(N__22653),
            .I(N__22650));
    Span4Mux_h I__5277 (
            .O(N__22650),
            .I(N__22647));
    Odrv4 I__5276 (
            .O(N__22647),
            .I(\ppm_encoder_1.pulses2count_9_i_1_4 ));
    InMux I__5275 (
            .O(N__22644),
            .I(N__22641));
    LocalMux I__5274 (
            .O(N__22641),
            .I(N__22636));
    CascadeMux I__5273 (
            .O(N__22640),
            .I(N__22633));
    InMux I__5272 (
            .O(N__22639),
            .I(N__22629));
    Span12Mux_s8_v I__5271 (
            .O(N__22636),
            .I(N__22626));
    InMux I__5270 (
            .O(N__22633),
            .I(N__22623));
    InMux I__5269 (
            .O(N__22632),
            .I(N__22620));
    LocalMux I__5268 (
            .O(N__22629),
            .I(N__22617));
    Odrv12 I__5267 (
            .O(N__22626),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__5266 (
            .O(N__22623),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__5265 (
            .O(N__22620),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    Odrv4 I__5264 (
            .O(N__22617),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__5263 (
            .O(N__22608),
            .I(N__22605));
    LocalMux I__5262 (
            .O(N__22605),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__5261 (
            .O(N__22602),
            .I(N__22599));
    LocalMux I__5260 (
            .O(N__22599),
            .I(N__22596));
    Span4Mux_h I__5259 (
            .O(N__22596),
            .I(N__22593));
    Odrv4 I__5258 (
            .O(N__22593),
            .I(\ppm_encoder_1.N_300 ));
    CascadeMux I__5257 (
            .O(N__22590),
            .I(N__22587));
    InMux I__5256 (
            .O(N__22587),
            .I(N__22584));
    LocalMux I__5255 (
            .O(N__22584),
            .I(N__22581));
    Odrv4 I__5254 (
            .O(N__22581),
            .I(\ppm_encoder_1.pulses2count_9_i_0_5 ));
    InMux I__5253 (
            .O(N__22578),
            .I(N__22573));
    CascadeMux I__5252 (
            .O(N__22577),
            .I(N__22570));
    CascadeMux I__5251 (
            .O(N__22576),
            .I(N__22566));
    LocalMux I__5250 (
            .O(N__22573),
            .I(N__22563));
    InMux I__5249 (
            .O(N__22570),
            .I(N__22560));
    InMux I__5248 (
            .O(N__22569),
            .I(N__22557));
    InMux I__5247 (
            .O(N__22566),
            .I(N__22554));
    Span4Mux_h I__5246 (
            .O(N__22563),
            .I(N__22549));
    LocalMux I__5245 (
            .O(N__22560),
            .I(N__22549));
    LocalMux I__5244 (
            .O(N__22557),
            .I(N__22544));
    LocalMux I__5243 (
            .O(N__22554),
            .I(N__22544));
    Odrv4 I__5242 (
            .O(N__22549),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    Odrv12 I__5241 (
            .O(N__22544),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    CascadeMux I__5240 (
            .O(N__22539),
            .I(N__22536));
    InMux I__5239 (
            .O(N__22536),
            .I(N__22533));
    LocalMux I__5238 (
            .O(N__22533),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    CascadeMux I__5237 (
            .O(N__22530),
            .I(N__22527));
    InMux I__5236 (
            .O(N__22527),
            .I(N__22522));
    InMux I__5235 (
            .O(N__22526),
            .I(N__22519));
    InMux I__5234 (
            .O(N__22525),
            .I(N__22516));
    LocalMux I__5233 (
            .O(N__22522),
            .I(N__22513));
    LocalMux I__5232 (
            .O(N__22519),
            .I(N__22509));
    LocalMux I__5231 (
            .O(N__22516),
            .I(N__22506));
    Span4Mux_v I__5230 (
            .O(N__22513),
            .I(N__22503));
    InMux I__5229 (
            .O(N__22512),
            .I(N__22500));
    Span4Mux_h I__5228 (
            .O(N__22509),
            .I(N__22495));
    Span4Mux_h I__5227 (
            .O(N__22506),
            .I(N__22495));
    Odrv4 I__5226 (
            .O(N__22503),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    LocalMux I__5225 (
            .O(N__22500),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__5224 (
            .O(N__22495),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__5223 (
            .O(N__22488),
            .I(N__22485));
    LocalMux I__5222 (
            .O(N__22485),
            .I(N__22482));
    Span4Mux_h I__5221 (
            .O(N__22482),
            .I(N__22479));
    Odrv4 I__5220 (
            .O(N__22479),
            .I(\ppm_encoder_1.pulses2count_9_i_1_10 ));
    InMux I__5219 (
            .O(N__22476),
            .I(N__22473));
    LocalMux I__5218 (
            .O(N__22473),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    CascadeMux I__5217 (
            .O(N__22470),
            .I(N__22465));
    CascadeMux I__5216 (
            .O(N__22469),
            .I(N__22462));
    InMux I__5215 (
            .O(N__22468),
            .I(N__22458));
    InMux I__5214 (
            .O(N__22465),
            .I(N__22455));
    InMux I__5213 (
            .O(N__22462),
            .I(N__22452));
    InMux I__5212 (
            .O(N__22461),
            .I(N__22449));
    LocalMux I__5211 (
            .O(N__22458),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__5210 (
            .O(N__22455),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__5209 (
            .O(N__22452),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__5208 (
            .O(N__22449),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    CascadeMux I__5207 (
            .O(N__22440),
            .I(N__22437));
    InMux I__5206 (
            .O(N__22437),
            .I(N__22434));
    LocalMux I__5205 (
            .O(N__22434),
            .I(N__22431));
    Odrv4 I__5204 (
            .O(N__22431),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    CascadeMux I__5203 (
            .O(N__22428),
            .I(N__22424));
    InMux I__5202 (
            .O(N__22427),
            .I(N__22420));
    InMux I__5201 (
            .O(N__22424),
            .I(N__22417));
    InMux I__5200 (
            .O(N__22423),
            .I(N__22414));
    LocalMux I__5199 (
            .O(N__22420),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__5198 (
            .O(N__22417),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__5197 (
            .O(N__22414),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__5196 (
            .O(N__22407),
            .I(N__22404));
    LocalMux I__5195 (
            .O(N__22404),
            .I(N__22401));
    Odrv4 I__5194 (
            .O(N__22401),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CascadeMux I__5193 (
            .O(N__22398),
            .I(N__22395));
    InMux I__5192 (
            .O(N__22395),
            .I(N__22392));
    LocalMux I__5191 (
            .O(N__22392),
            .I(N__22389));
    Odrv4 I__5190 (
            .O(N__22389),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__5189 (
            .O(N__22386),
            .I(N__22381));
    InMux I__5188 (
            .O(N__22385),
            .I(N__22378));
    InMux I__5187 (
            .O(N__22384),
            .I(N__22375));
    LocalMux I__5186 (
            .O(N__22381),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5185 (
            .O(N__22378),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5184 (
            .O(N__22375),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__5183 (
            .O(N__22368),
            .I(N__22363));
    InMux I__5182 (
            .O(N__22367),
            .I(N__22360));
    InMux I__5181 (
            .O(N__22366),
            .I(N__22357));
    LocalMux I__5180 (
            .O(N__22363),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__5179 (
            .O(N__22360),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__5178 (
            .O(N__22357),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    CascadeMux I__5177 (
            .O(N__22350),
            .I(N__22346));
    InMux I__5176 (
            .O(N__22349),
            .I(N__22342));
    InMux I__5175 (
            .O(N__22346),
            .I(N__22339));
    InMux I__5174 (
            .O(N__22345),
            .I(N__22336));
    LocalMux I__5173 (
            .O(N__22342),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__5172 (
            .O(N__22339),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__5171 (
            .O(N__22336),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__5170 (
            .O(N__22329),
            .I(N__22324));
    InMux I__5169 (
            .O(N__22328),
            .I(N__22321));
    InMux I__5168 (
            .O(N__22327),
            .I(N__22318));
    LocalMux I__5167 (
            .O(N__22324),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__5166 (
            .O(N__22321),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__5165 (
            .O(N__22318),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__5164 (
            .O(N__22311),
            .I(N__22307));
    CascadeMux I__5163 (
            .O(N__22310),
            .I(N__22304));
    LocalMux I__5162 (
            .O(N__22307),
            .I(N__22300));
    InMux I__5161 (
            .O(N__22304),
            .I(N__22297));
    InMux I__5160 (
            .O(N__22303),
            .I(N__22294));
    Odrv12 I__5159 (
            .O(N__22300),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    LocalMux I__5158 (
            .O(N__22297),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    LocalMux I__5157 (
            .O(N__22294),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    CascadeMux I__5156 (
            .O(N__22287),
            .I(N__22284));
    InMux I__5155 (
            .O(N__22284),
            .I(N__22280));
    CascadeMux I__5154 (
            .O(N__22283),
            .I(N__22276));
    LocalMux I__5153 (
            .O(N__22280),
            .I(N__22273));
    CascadeMux I__5152 (
            .O(N__22279),
            .I(N__22270));
    InMux I__5151 (
            .O(N__22276),
            .I(N__22266));
    Span4Mux_h I__5150 (
            .O(N__22273),
            .I(N__22263));
    InMux I__5149 (
            .O(N__22270),
            .I(N__22258));
    InMux I__5148 (
            .O(N__22269),
            .I(N__22258));
    LocalMux I__5147 (
            .O(N__22266),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__5146 (
            .O(N__22263),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    LocalMux I__5145 (
            .O(N__22258),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    CascadeMux I__5144 (
            .O(N__22251),
            .I(N__22248));
    InMux I__5143 (
            .O(N__22248),
            .I(N__22245));
    LocalMux I__5142 (
            .O(N__22245),
            .I(N__22242));
    Span4Mux_h I__5141 (
            .O(N__22242),
            .I(N__22239));
    Odrv4 I__5140 (
            .O(N__22239),
            .I(\ppm_encoder_1.pulses2count_9_i_0_7 ));
    InMux I__5139 (
            .O(N__22236),
            .I(N__22232));
    CascadeMux I__5138 (
            .O(N__22235),
            .I(N__22228));
    LocalMux I__5137 (
            .O(N__22232),
            .I(N__22225));
    InMux I__5136 (
            .O(N__22231),
            .I(N__22222));
    InMux I__5135 (
            .O(N__22228),
            .I(N__22219));
    Span4Mux_h I__5134 (
            .O(N__22225),
            .I(N__22216));
    LocalMux I__5133 (
            .O(N__22222),
            .I(N__22213));
    LocalMux I__5132 (
            .O(N__22219),
            .I(N__22210));
    Span4Mux_h I__5131 (
            .O(N__22216),
            .I(N__22207));
    Span4Mux_v I__5130 (
            .O(N__22213),
            .I(N__22204));
    Span4Mux_h I__5129 (
            .O(N__22210),
            .I(N__22201));
    Odrv4 I__5128 (
            .O(N__22207),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__5127 (
            .O(N__22204),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__5126 (
            .O(N__22201),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__5125 (
            .O(N__22194),
            .I(N__22191));
    LocalMux I__5124 (
            .O(N__22191),
            .I(N__22188));
    Span4Mux_h I__5123 (
            .O(N__22188),
            .I(N__22182));
    InMux I__5122 (
            .O(N__22187),
            .I(N__22179));
    InMux I__5121 (
            .O(N__22186),
            .I(N__22176));
    InMux I__5120 (
            .O(N__22185),
            .I(N__22173));
    Odrv4 I__5119 (
            .O(N__22182),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__5118 (
            .O(N__22179),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__5117 (
            .O(N__22176),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__5116 (
            .O(N__22173),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    CascadeMux I__5115 (
            .O(N__22164),
            .I(N__22161));
    InMux I__5114 (
            .O(N__22161),
            .I(N__22158));
    LocalMux I__5113 (
            .O(N__22158),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__5112 (
            .O(N__22155),
            .I(N__22151));
    InMux I__5111 (
            .O(N__22154),
            .I(N__22147));
    LocalMux I__5110 (
            .O(N__22151),
            .I(N__22144));
    InMux I__5109 (
            .O(N__22150),
            .I(N__22141));
    LocalMux I__5108 (
            .O(N__22147),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__5107 (
            .O(N__22144),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__5106 (
            .O(N__22141),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    CascadeMux I__5105 (
            .O(N__22134),
            .I(N__22129));
    CascadeMux I__5104 (
            .O(N__22133),
            .I(N__22126));
    InMux I__5103 (
            .O(N__22132),
            .I(N__22111));
    InMux I__5102 (
            .O(N__22129),
            .I(N__22111));
    InMux I__5101 (
            .O(N__22126),
            .I(N__22105));
    InMux I__5100 (
            .O(N__22125),
            .I(N__22105));
    InMux I__5099 (
            .O(N__22124),
            .I(N__22102));
    InMux I__5098 (
            .O(N__22123),
            .I(N__22099));
    InMux I__5097 (
            .O(N__22122),
            .I(N__22091));
    InMux I__5096 (
            .O(N__22121),
            .I(N__22091));
    InMux I__5095 (
            .O(N__22120),
            .I(N__22084));
    InMux I__5094 (
            .O(N__22119),
            .I(N__22084));
    InMux I__5093 (
            .O(N__22118),
            .I(N__22084));
    InMux I__5092 (
            .O(N__22117),
            .I(N__22079));
    InMux I__5091 (
            .O(N__22116),
            .I(N__22079));
    LocalMux I__5090 (
            .O(N__22111),
            .I(N__22076));
    InMux I__5089 (
            .O(N__22110),
            .I(N__22073));
    LocalMux I__5088 (
            .O(N__22105),
            .I(N__22069));
    LocalMux I__5087 (
            .O(N__22102),
            .I(N__22063));
    LocalMux I__5086 (
            .O(N__22099),
            .I(N__22063));
    CascadeMux I__5085 (
            .O(N__22098),
            .I(N__22060));
    InMux I__5084 (
            .O(N__22097),
            .I(N__22053));
    InMux I__5083 (
            .O(N__22096),
            .I(N__22053));
    LocalMux I__5082 (
            .O(N__22091),
            .I(N__22050));
    LocalMux I__5081 (
            .O(N__22084),
            .I(N__22045));
    LocalMux I__5080 (
            .O(N__22079),
            .I(N__22045));
    Span4Mux_v I__5079 (
            .O(N__22076),
            .I(N__22042));
    LocalMux I__5078 (
            .O(N__22073),
            .I(N__22039));
    InMux I__5077 (
            .O(N__22072),
            .I(N__22036));
    Span4Mux_h I__5076 (
            .O(N__22069),
            .I(N__22033));
    InMux I__5075 (
            .O(N__22068),
            .I(N__22030));
    Span4Mux_v I__5074 (
            .O(N__22063),
            .I(N__22027));
    InMux I__5073 (
            .O(N__22060),
            .I(N__22020));
    InMux I__5072 (
            .O(N__22059),
            .I(N__22020));
    InMux I__5071 (
            .O(N__22058),
            .I(N__22020));
    LocalMux I__5070 (
            .O(N__22053),
            .I(N__22015));
    Span4Mux_h I__5069 (
            .O(N__22050),
            .I(N__22015));
    Span4Mux_v I__5068 (
            .O(N__22045),
            .I(N__22008));
    Span4Mux_h I__5067 (
            .O(N__22042),
            .I(N__22008));
    Span4Mux_h I__5066 (
            .O(N__22039),
            .I(N__22008));
    LocalMux I__5065 (
            .O(N__22036),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__5064 (
            .O(N__22033),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__5063 (
            .O(N__22030),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__5062 (
            .O(N__22027),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__5061 (
            .O(N__22020),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__5060 (
            .O(N__22015),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__5059 (
            .O(N__22008),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__5058 (
            .O(N__21993),
            .I(N__21982));
    InMux I__5057 (
            .O(N__21992),
            .I(N__21982));
    InMux I__5056 (
            .O(N__21991),
            .I(N__21982));
    InMux I__5055 (
            .O(N__21990),
            .I(N__21968));
    InMux I__5054 (
            .O(N__21989),
            .I(N__21968));
    LocalMux I__5053 (
            .O(N__21982),
            .I(N__21961));
    InMux I__5052 (
            .O(N__21981),
            .I(N__21954));
    InMux I__5051 (
            .O(N__21980),
            .I(N__21954));
    InMux I__5050 (
            .O(N__21979),
            .I(N__21954));
    InMux I__5049 (
            .O(N__21978),
            .I(N__21951));
    InMux I__5048 (
            .O(N__21977),
            .I(N__21948));
    InMux I__5047 (
            .O(N__21976),
            .I(N__21943));
    InMux I__5046 (
            .O(N__21975),
            .I(N__21943));
    InMux I__5045 (
            .O(N__21974),
            .I(N__21939));
    InMux I__5044 (
            .O(N__21973),
            .I(N__21936));
    LocalMux I__5043 (
            .O(N__21968),
            .I(N__21933));
    InMux I__5042 (
            .O(N__21967),
            .I(N__21930));
    InMux I__5041 (
            .O(N__21966),
            .I(N__21925));
    InMux I__5040 (
            .O(N__21965),
            .I(N__21920));
    InMux I__5039 (
            .O(N__21964),
            .I(N__21920));
    Span4Mux_v I__5038 (
            .O(N__21961),
            .I(N__21915));
    LocalMux I__5037 (
            .O(N__21954),
            .I(N__21915));
    LocalMux I__5036 (
            .O(N__21951),
            .I(N__21908));
    LocalMux I__5035 (
            .O(N__21948),
            .I(N__21908));
    LocalMux I__5034 (
            .O(N__21943),
            .I(N__21908));
    InMux I__5033 (
            .O(N__21942),
            .I(N__21904));
    LocalMux I__5032 (
            .O(N__21939),
            .I(N__21901));
    LocalMux I__5031 (
            .O(N__21936),
            .I(N__21896));
    Span4Mux_v I__5030 (
            .O(N__21933),
            .I(N__21896));
    LocalMux I__5029 (
            .O(N__21930),
            .I(N__21893));
    InMux I__5028 (
            .O(N__21929),
            .I(N__21888));
    InMux I__5027 (
            .O(N__21928),
            .I(N__21888));
    LocalMux I__5026 (
            .O(N__21925),
            .I(N__21883));
    LocalMux I__5025 (
            .O(N__21920),
            .I(N__21883));
    Span4Mux_v I__5024 (
            .O(N__21915),
            .I(N__21875));
    Span4Mux_v I__5023 (
            .O(N__21908),
            .I(N__21875));
    InMux I__5022 (
            .O(N__21907),
            .I(N__21872));
    LocalMux I__5021 (
            .O(N__21904),
            .I(N__21869));
    Span4Mux_v I__5020 (
            .O(N__21901),
            .I(N__21864));
    Span4Mux_h I__5019 (
            .O(N__21896),
            .I(N__21864));
    Span4Mux_h I__5018 (
            .O(N__21893),
            .I(N__21861));
    LocalMux I__5017 (
            .O(N__21888),
            .I(N__21856));
    Span4Mux_v I__5016 (
            .O(N__21883),
            .I(N__21856));
    InMux I__5015 (
            .O(N__21882),
            .I(N__21849));
    InMux I__5014 (
            .O(N__21881),
            .I(N__21849));
    InMux I__5013 (
            .O(N__21880),
            .I(N__21849));
    Span4Mux_h I__5012 (
            .O(N__21875),
            .I(N__21844));
    LocalMux I__5011 (
            .O(N__21872),
            .I(N__21844));
    Odrv4 I__5010 (
            .O(N__21869),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__5009 (
            .O(N__21864),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__5008 (
            .O(N__21861),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__5007 (
            .O(N__21856),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__5006 (
            .O(N__21849),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__5005 (
            .O(N__21844),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    CascadeMux I__5004 (
            .O(N__21831),
            .I(N__21827));
    CascadeMux I__5003 (
            .O(N__21830),
            .I(N__21824));
    InMux I__5002 (
            .O(N__21827),
            .I(N__21821));
    InMux I__5001 (
            .O(N__21824),
            .I(N__21818));
    LocalMux I__5000 (
            .O(N__21821),
            .I(N__21814));
    LocalMux I__4999 (
            .O(N__21818),
            .I(N__21810));
    CascadeMux I__4998 (
            .O(N__21817),
            .I(N__21807));
    Span4Mux_h I__4997 (
            .O(N__21814),
            .I(N__21804));
    InMux I__4996 (
            .O(N__21813),
            .I(N__21801));
    Span4Mux_h I__4995 (
            .O(N__21810),
            .I(N__21798));
    InMux I__4994 (
            .O(N__21807),
            .I(N__21795));
    Odrv4 I__4993 (
            .O(N__21804),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__4992 (
            .O(N__21801),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    Odrv4 I__4991 (
            .O(N__21798),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__4990 (
            .O(N__21795),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    CascadeMux I__4989 (
            .O(N__21786),
            .I(N__21782));
    InMux I__4988 (
            .O(N__21785),
            .I(N__21769));
    InMux I__4987 (
            .O(N__21782),
            .I(N__21766));
    InMux I__4986 (
            .O(N__21781),
            .I(N__21763));
    InMux I__4985 (
            .O(N__21780),
            .I(N__21753));
    InMux I__4984 (
            .O(N__21779),
            .I(N__21753));
    InMux I__4983 (
            .O(N__21778),
            .I(N__21753));
    InMux I__4982 (
            .O(N__21777),
            .I(N__21744));
    InMux I__4981 (
            .O(N__21776),
            .I(N__21744));
    InMux I__4980 (
            .O(N__21775),
            .I(N__21744));
    InMux I__4979 (
            .O(N__21774),
            .I(N__21744));
    CascadeMux I__4978 (
            .O(N__21773),
            .I(N__21741));
    InMux I__4977 (
            .O(N__21772),
            .I(N__21738));
    LocalMux I__4976 (
            .O(N__21769),
            .I(N__21735));
    LocalMux I__4975 (
            .O(N__21766),
            .I(N__21730));
    LocalMux I__4974 (
            .O(N__21763),
            .I(N__21727));
    InMux I__4973 (
            .O(N__21762),
            .I(N__21722));
    InMux I__4972 (
            .O(N__21761),
            .I(N__21722));
    InMux I__4971 (
            .O(N__21760),
            .I(N__21719));
    LocalMux I__4970 (
            .O(N__21753),
            .I(N__21716));
    LocalMux I__4969 (
            .O(N__21744),
            .I(N__21713));
    InMux I__4968 (
            .O(N__21741),
            .I(N__21710));
    LocalMux I__4967 (
            .O(N__21738),
            .I(N__21707));
    Span4Mux_h I__4966 (
            .O(N__21735),
            .I(N__21704));
    CascadeMux I__4965 (
            .O(N__21734),
            .I(N__21699));
    CascadeMux I__4964 (
            .O(N__21733),
            .I(N__21696));
    Span4Mux_v I__4963 (
            .O(N__21730),
            .I(N__21691));
    Span4Mux_h I__4962 (
            .O(N__21727),
            .I(N__21691));
    LocalMux I__4961 (
            .O(N__21722),
            .I(N__21688));
    LocalMux I__4960 (
            .O(N__21719),
            .I(N__21679));
    Span4Mux_v I__4959 (
            .O(N__21716),
            .I(N__21679));
    Span4Mux_v I__4958 (
            .O(N__21713),
            .I(N__21676));
    LocalMux I__4957 (
            .O(N__21710),
            .I(N__21669));
    Span4Mux_h I__4956 (
            .O(N__21707),
            .I(N__21669));
    Span4Mux_v I__4955 (
            .O(N__21704),
            .I(N__21669));
    InMux I__4954 (
            .O(N__21703),
            .I(N__21666));
    InMux I__4953 (
            .O(N__21702),
            .I(N__21659));
    InMux I__4952 (
            .O(N__21699),
            .I(N__21659));
    InMux I__4951 (
            .O(N__21696),
            .I(N__21659));
    Span4Mux_v I__4950 (
            .O(N__21691),
            .I(N__21654));
    Span4Mux_h I__4949 (
            .O(N__21688),
            .I(N__21654));
    InMux I__4948 (
            .O(N__21687),
            .I(N__21651));
    InMux I__4947 (
            .O(N__21686),
            .I(N__21644));
    InMux I__4946 (
            .O(N__21685),
            .I(N__21644));
    InMux I__4945 (
            .O(N__21684),
            .I(N__21644));
    Span4Mux_v I__4944 (
            .O(N__21679),
            .I(N__21637));
    Span4Mux_v I__4943 (
            .O(N__21676),
            .I(N__21637));
    Span4Mux_v I__4942 (
            .O(N__21669),
            .I(N__21637));
    LocalMux I__4941 (
            .O(N__21666),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4940 (
            .O(N__21659),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__4939 (
            .O(N__21654),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4938 (
            .O(N__21651),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4937 (
            .O(N__21644),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__4936 (
            .O(N__21637),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__4935 (
            .O(N__21624),
            .I(N__21615));
    CascadeMux I__4934 (
            .O(N__21623),
            .I(N__21611));
    InMux I__4933 (
            .O(N__21622),
            .I(N__21606));
    CascadeMux I__4932 (
            .O(N__21621),
            .I(N__21603));
    CascadeMux I__4931 (
            .O(N__21620),
            .I(N__21599));
    InMux I__4930 (
            .O(N__21619),
            .I(N__21594));
    InMux I__4929 (
            .O(N__21618),
            .I(N__21594));
    InMux I__4928 (
            .O(N__21615),
            .I(N__21585));
    InMux I__4927 (
            .O(N__21614),
            .I(N__21585));
    InMux I__4926 (
            .O(N__21611),
            .I(N__21585));
    InMux I__4925 (
            .O(N__21610),
            .I(N__21585));
    CascadeMux I__4924 (
            .O(N__21609),
            .I(N__21582));
    LocalMux I__4923 (
            .O(N__21606),
            .I(N__21579));
    InMux I__4922 (
            .O(N__21603),
            .I(N__21576));
    InMux I__4921 (
            .O(N__21602),
            .I(N__21571));
    InMux I__4920 (
            .O(N__21599),
            .I(N__21571));
    LocalMux I__4919 (
            .O(N__21594),
            .I(N__21566));
    LocalMux I__4918 (
            .O(N__21585),
            .I(N__21566));
    InMux I__4917 (
            .O(N__21582),
            .I(N__21563));
    Span4Mux_s3_v I__4916 (
            .O(N__21579),
            .I(N__21558));
    LocalMux I__4915 (
            .O(N__21576),
            .I(N__21558));
    LocalMux I__4914 (
            .O(N__21571),
            .I(N__21555));
    Span4Mux_v I__4913 (
            .O(N__21566),
            .I(N__21552));
    LocalMux I__4912 (
            .O(N__21563),
            .I(N__21545));
    Span4Mux_v I__4911 (
            .O(N__21558),
            .I(N__21545));
    Span4Mux_v I__4910 (
            .O(N__21555),
            .I(N__21545));
    Odrv4 I__4909 (
            .O(N__21552),
            .I(\ppm_encoder_1.N_235 ));
    Odrv4 I__4908 (
            .O(N__21545),
            .I(\ppm_encoder_1.N_235 ));
    InMux I__4907 (
            .O(N__21540),
            .I(N__21536));
    InMux I__4906 (
            .O(N__21539),
            .I(N__21533));
    LocalMux I__4905 (
            .O(N__21536),
            .I(N__21530));
    LocalMux I__4904 (
            .O(N__21533),
            .I(N__21527));
    Span4Mux_v I__4903 (
            .O(N__21530),
            .I(N__21524));
    Span12Mux_h I__4902 (
            .O(N__21527),
            .I(N__21521));
    Span4Mux_h I__4901 (
            .O(N__21524),
            .I(N__21518));
    Odrv12 I__4900 (
            .O(N__21521),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv4 I__4899 (
            .O(N__21518),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__4898 (
            .O(N__21513),
            .I(N__21508));
    CascadeMux I__4897 (
            .O(N__21512),
            .I(N__21504));
    InMux I__4896 (
            .O(N__21511),
            .I(N__21501));
    LocalMux I__4895 (
            .O(N__21508),
            .I(N__21498));
    InMux I__4894 (
            .O(N__21507),
            .I(N__21495));
    InMux I__4893 (
            .O(N__21504),
            .I(N__21492));
    LocalMux I__4892 (
            .O(N__21501),
            .I(N__21489));
    Span4Mux_h I__4891 (
            .O(N__21498),
            .I(N__21484));
    LocalMux I__4890 (
            .O(N__21495),
            .I(N__21484));
    LocalMux I__4889 (
            .O(N__21492),
            .I(N__21481));
    Span4Mux_s3_v I__4888 (
            .O(N__21489),
            .I(N__21476));
    Span4Mux_v I__4887 (
            .O(N__21484),
            .I(N__21476));
    Odrv4 I__4886 (
            .O(N__21481),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__4885 (
            .O(N__21476),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    CascadeMux I__4884 (
            .O(N__21471),
            .I(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ));
    InMux I__4883 (
            .O(N__21468),
            .I(N__21465));
    LocalMux I__4882 (
            .O(N__21465),
            .I(N__21462));
    Span12Mux_h I__4881 (
            .O(N__21462),
            .I(N__21458));
    InMux I__4880 (
            .O(N__21461),
            .I(N__21455));
    Odrv12 I__4879 (
            .O(N__21458),
            .I(\ppm_encoder_1.N_304 ));
    LocalMux I__4878 (
            .O(N__21455),
            .I(\ppm_encoder_1.N_304 ));
    InMux I__4877 (
            .O(N__21450),
            .I(N__21446));
    InMux I__4876 (
            .O(N__21449),
            .I(N__21442));
    LocalMux I__4875 (
            .O(N__21446),
            .I(N__21439));
    InMux I__4874 (
            .O(N__21445),
            .I(N__21436));
    LocalMux I__4873 (
            .O(N__21442),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__4872 (
            .O(N__21439),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__4871 (
            .O(N__21436),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__4870 (
            .O(N__21429),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__4869 (
            .O(N__21426),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__4868 (
            .O(N__21423),
            .I(N__21414));
    SRMux I__4867 (
            .O(N__21422),
            .I(N__21414));
    SRMux I__4866 (
            .O(N__21421),
            .I(N__21414));
    GlobalMux I__4865 (
            .O(N__21414),
            .I(N__21411));
    gio2CtrlBuf I__4864 (
            .O(N__21411),
            .I(\ppm_encoder_1.N_512_g ));
    InMux I__4863 (
            .O(N__21408),
            .I(N__21404));
    InMux I__4862 (
            .O(N__21407),
            .I(N__21401));
    LocalMux I__4861 (
            .O(N__21404),
            .I(N__21398));
    LocalMux I__4860 (
            .O(N__21401),
            .I(N__21395));
    Span4Mux_v I__4859 (
            .O(N__21398),
            .I(N__21389));
    Span4Mux_h I__4858 (
            .O(N__21395),
            .I(N__21389));
    InMux I__4857 (
            .O(N__21394),
            .I(N__21386));
    Odrv4 I__4856 (
            .O(N__21389),
            .I(\ppm_encoder_1.N_247 ));
    LocalMux I__4855 (
            .O(N__21386),
            .I(\ppm_encoder_1.N_247 ));
    InMux I__4854 (
            .O(N__21381),
            .I(N__21378));
    LocalMux I__4853 (
            .O(N__21378),
            .I(\ppm_encoder_1.pulses2count_9_0_2_11 ));
    CascadeMux I__4852 (
            .O(N__21375),
            .I(N__21372));
    InMux I__4851 (
            .O(N__21372),
            .I(N__21369));
    LocalMux I__4850 (
            .O(N__21369),
            .I(\ppm_encoder_1.N_388 ));
    InMux I__4849 (
            .O(N__21366),
            .I(N__21363));
    LocalMux I__4848 (
            .O(N__21363),
            .I(N__21360));
    Span4Mux_h I__4847 (
            .O(N__21360),
            .I(N__21357));
    Span4Mux_v I__4846 (
            .O(N__21357),
            .I(N__21354));
    Odrv4 I__4845 (
            .O(N__21354),
            .I(\ppm_encoder_1.pulses2count_9_0_0_11 ));
    CascadeMux I__4844 (
            .O(N__21351),
            .I(N__21346));
    InMux I__4843 (
            .O(N__21350),
            .I(N__21343));
    InMux I__4842 (
            .O(N__21349),
            .I(N__21340));
    InMux I__4841 (
            .O(N__21346),
            .I(N__21337));
    LocalMux I__4840 (
            .O(N__21343),
            .I(N__21333));
    LocalMux I__4839 (
            .O(N__21340),
            .I(N__21330));
    LocalMux I__4838 (
            .O(N__21337),
            .I(N__21327));
    CascadeMux I__4837 (
            .O(N__21336),
            .I(N__21324));
    Span4Mux_h I__4836 (
            .O(N__21333),
            .I(N__21321));
    Sp12to4 I__4835 (
            .O(N__21330),
            .I(N__21318));
    Span4Mux_h I__4834 (
            .O(N__21327),
            .I(N__21315));
    InMux I__4833 (
            .O(N__21324),
            .I(N__21312));
    Odrv4 I__4832 (
            .O(N__21321),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv12 I__4831 (
            .O(N__21318),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__4830 (
            .O(N__21315),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__4829 (
            .O(N__21312),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    CascadeMux I__4828 (
            .O(N__21303),
            .I(N__21300));
    InMux I__4827 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__4826 (
            .O(N__21297),
            .I(\ppm_encoder_1.pulses2count_9_0_0_13 ));
    InMux I__4825 (
            .O(N__21294),
            .I(N__21291));
    LocalMux I__4824 (
            .O(N__21291),
            .I(N__21288));
    Span4Mux_v I__4823 (
            .O(N__21288),
            .I(N__21284));
    InMux I__4822 (
            .O(N__21287),
            .I(N__21281));
    Odrv4 I__4821 (
            .O(N__21284),
            .I(\ppm_encoder_1.N_303 ));
    LocalMux I__4820 (
            .O(N__21281),
            .I(\ppm_encoder_1.N_303 ));
    CascadeMux I__4819 (
            .O(N__21276),
            .I(N__21273));
    InMux I__4818 (
            .O(N__21273),
            .I(N__21268));
    CascadeMux I__4817 (
            .O(N__21272),
            .I(N__21265));
    CascadeMux I__4816 (
            .O(N__21271),
            .I(N__21262));
    LocalMux I__4815 (
            .O(N__21268),
            .I(N__21259));
    InMux I__4814 (
            .O(N__21265),
            .I(N__21256));
    InMux I__4813 (
            .O(N__21262),
            .I(N__21253));
    Span4Mux_h I__4812 (
            .O(N__21259),
            .I(N__21248));
    LocalMux I__4811 (
            .O(N__21256),
            .I(N__21248));
    LocalMux I__4810 (
            .O(N__21253),
            .I(N__21245));
    Span4Mux_h I__4809 (
            .O(N__21248),
            .I(N__21242));
    Span4Mux_h I__4808 (
            .O(N__21245),
            .I(N__21239));
    Odrv4 I__4807 (
            .O(N__21242),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__4806 (
            .O(N__21239),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__4805 (
            .O(N__21234),
            .I(N__21224));
    InMux I__4804 (
            .O(N__21233),
            .I(N__21192));
    InMux I__4803 (
            .O(N__21232),
            .I(N__21192));
    InMux I__4802 (
            .O(N__21231),
            .I(N__21192));
    InMux I__4801 (
            .O(N__21230),
            .I(N__21192));
    InMux I__4800 (
            .O(N__21229),
            .I(N__21187));
    InMux I__4799 (
            .O(N__21228),
            .I(N__21187));
    CascadeMux I__4798 (
            .O(N__21227),
            .I(N__21184));
    LocalMux I__4797 (
            .O(N__21224),
            .I(N__21181));
    InMux I__4796 (
            .O(N__21223),
            .I(N__21178));
    InMux I__4795 (
            .O(N__21222),
            .I(N__21173));
    InMux I__4794 (
            .O(N__21221),
            .I(N__21173));
    InMux I__4793 (
            .O(N__21220),
            .I(N__21170));
    InMux I__4792 (
            .O(N__21219),
            .I(N__21164));
    InMux I__4791 (
            .O(N__21218),
            .I(N__21155));
    InMux I__4790 (
            .O(N__21217),
            .I(N__21155));
    InMux I__4789 (
            .O(N__21216),
            .I(N__21155));
    InMux I__4788 (
            .O(N__21215),
            .I(N__21155));
    InMux I__4787 (
            .O(N__21214),
            .I(N__21146));
    InMux I__4786 (
            .O(N__21213),
            .I(N__21146));
    InMux I__4785 (
            .O(N__21212),
            .I(N__21146));
    InMux I__4784 (
            .O(N__21211),
            .I(N__21146));
    InMux I__4783 (
            .O(N__21210),
            .I(N__21140));
    InMux I__4782 (
            .O(N__21209),
            .I(N__21140));
    InMux I__4781 (
            .O(N__21208),
            .I(N__21131));
    InMux I__4780 (
            .O(N__21207),
            .I(N__21131));
    InMux I__4779 (
            .O(N__21206),
            .I(N__21131));
    InMux I__4778 (
            .O(N__21205),
            .I(N__21131));
    InMux I__4777 (
            .O(N__21204),
            .I(N__21123));
    InMux I__4776 (
            .O(N__21203),
            .I(N__21123));
    InMux I__4775 (
            .O(N__21202),
            .I(N__21123));
    InMux I__4774 (
            .O(N__21201),
            .I(N__21120));
    LocalMux I__4773 (
            .O(N__21192),
            .I(N__21115));
    LocalMux I__4772 (
            .O(N__21187),
            .I(N__21115));
    InMux I__4771 (
            .O(N__21184),
            .I(N__21112));
    Span4Mux_h I__4770 (
            .O(N__21181),
            .I(N__21109));
    LocalMux I__4769 (
            .O(N__21178),
            .I(N__21106));
    LocalMux I__4768 (
            .O(N__21173),
            .I(N__21101));
    LocalMux I__4767 (
            .O(N__21170),
            .I(N__21101));
    CascadeMux I__4766 (
            .O(N__21169),
            .I(N__21094));
    CascadeMux I__4765 (
            .O(N__21168),
            .I(N__21091));
    InMux I__4764 (
            .O(N__21167),
            .I(N__21080));
    LocalMux I__4763 (
            .O(N__21164),
            .I(N__21073));
    LocalMux I__4762 (
            .O(N__21155),
            .I(N__21073));
    LocalMux I__4761 (
            .O(N__21146),
            .I(N__21073));
    InMux I__4760 (
            .O(N__21145),
            .I(N__21070));
    LocalMux I__4759 (
            .O(N__21140),
            .I(N__21065));
    LocalMux I__4758 (
            .O(N__21131),
            .I(N__21065));
    CascadeMux I__4757 (
            .O(N__21130),
            .I(N__21057));
    LocalMux I__4756 (
            .O(N__21123),
            .I(N__21044));
    LocalMux I__4755 (
            .O(N__21120),
            .I(N__21044));
    Span4Mux_v I__4754 (
            .O(N__21115),
            .I(N__21044));
    LocalMux I__4753 (
            .O(N__21112),
            .I(N__21044));
    Sp12to4 I__4752 (
            .O(N__21109),
            .I(N__21041));
    Span4Mux_v I__4751 (
            .O(N__21106),
            .I(N__21038));
    Span4Mux_v I__4750 (
            .O(N__21101),
            .I(N__21035));
    InMux I__4749 (
            .O(N__21100),
            .I(N__21032));
    InMux I__4748 (
            .O(N__21099),
            .I(N__21021));
    InMux I__4747 (
            .O(N__21098),
            .I(N__21021));
    InMux I__4746 (
            .O(N__21097),
            .I(N__21021));
    InMux I__4745 (
            .O(N__21094),
            .I(N__21021));
    InMux I__4744 (
            .O(N__21091),
            .I(N__21021));
    InMux I__4743 (
            .O(N__21090),
            .I(N__21010));
    InMux I__4742 (
            .O(N__21089),
            .I(N__21010));
    InMux I__4741 (
            .O(N__21088),
            .I(N__21010));
    InMux I__4740 (
            .O(N__21087),
            .I(N__21010));
    InMux I__4739 (
            .O(N__21086),
            .I(N__21010));
    InMux I__4738 (
            .O(N__21085),
            .I(N__21005));
    InMux I__4737 (
            .O(N__21084),
            .I(N__21005));
    InMux I__4736 (
            .O(N__21083),
            .I(N__21002));
    LocalMux I__4735 (
            .O(N__21080),
            .I(N__20993));
    Span4Mux_v I__4734 (
            .O(N__21073),
            .I(N__20993));
    LocalMux I__4733 (
            .O(N__21070),
            .I(N__20993));
    Span4Mux_h I__4732 (
            .O(N__21065),
            .I(N__20993));
    InMux I__4731 (
            .O(N__21064),
            .I(N__20984));
    InMux I__4730 (
            .O(N__21063),
            .I(N__20984));
    InMux I__4729 (
            .O(N__21062),
            .I(N__20984));
    InMux I__4728 (
            .O(N__21061),
            .I(N__20984));
    InMux I__4727 (
            .O(N__21060),
            .I(N__20979));
    InMux I__4726 (
            .O(N__21057),
            .I(N__20979));
    InMux I__4725 (
            .O(N__21056),
            .I(N__20970));
    InMux I__4724 (
            .O(N__21055),
            .I(N__20970));
    InMux I__4723 (
            .O(N__21054),
            .I(N__20970));
    InMux I__4722 (
            .O(N__21053),
            .I(N__20970));
    Odrv4 I__4721 (
            .O(N__21044),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv12 I__4720 (
            .O(N__21041),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv4 I__4719 (
            .O(N__21038),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv4 I__4718 (
            .O(N__21035),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4717 (
            .O(N__21032),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4716 (
            .O(N__21021),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4715 (
            .O(N__21010),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4714 (
            .O(N__21005),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4713 (
            .O(N__21002),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    Odrv4 I__4712 (
            .O(N__20993),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4711 (
            .O(N__20984),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4710 (
            .O(N__20979),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    LocalMux I__4709 (
            .O(N__20970),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ));
    IoInMux I__4708 (
            .O(N__20943),
            .I(N__20940));
    LocalMux I__4707 (
            .O(N__20940),
            .I(N__20937));
    Span12Mux_s6_v I__4706 (
            .O(N__20937),
            .I(N__20934));
    Odrv12 I__4705 (
            .O(N__20934),
            .I(\ppm_encoder_1.N_238_i_0 ));
    CascadeMux I__4704 (
            .O(N__20931),
            .I(N__20927));
    InMux I__4703 (
            .O(N__20930),
            .I(N__20923));
    InMux I__4702 (
            .O(N__20927),
            .I(N__20920));
    CascadeMux I__4701 (
            .O(N__20926),
            .I(N__20917));
    LocalMux I__4700 (
            .O(N__20923),
            .I(N__20914));
    LocalMux I__4699 (
            .O(N__20920),
            .I(N__20911));
    InMux I__4698 (
            .O(N__20917),
            .I(N__20908));
    Span4Mux_h I__4697 (
            .O(N__20914),
            .I(N__20905));
    Span4Mux_v I__4696 (
            .O(N__20911),
            .I(N__20902));
    LocalMux I__4695 (
            .O(N__20908),
            .I(N__20899));
    Span4Mux_v I__4694 (
            .O(N__20905),
            .I(N__20894));
    Span4Mux_v I__4693 (
            .O(N__20902),
            .I(N__20894));
    Odrv4 I__4692 (
            .O(N__20899),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    Odrv4 I__4691 (
            .O(N__20894),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__4690 (
            .O(N__20889),
            .I(N__20886));
    InMux I__4689 (
            .O(N__20886),
            .I(N__20882));
    InMux I__4688 (
            .O(N__20885),
            .I(N__20879));
    LocalMux I__4687 (
            .O(N__20882),
            .I(N__20876));
    LocalMux I__4686 (
            .O(N__20879),
            .I(N__20872));
    Span4Mux_h I__4685 (
            .O(N__20876),
            .I(N__20869));
    InMux I__4684 (
            .O(N__20875),
            .I(N__20866));
    Span4Mux_v I__4683 (
            .O(N__20872),
            .I(N__20863));
    Odrv4 I__4682 (
            .O(N__20869),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__4681 (
            .O(N__20866),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__4680 (
            .O(N__20863),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__4679 (
            .O(N__20856),
            .I(bfn_11_25_0_));
    InMux I__4678 (
            .O(N__20853),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__4677 (
            .O(N__20850),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__4676 (
            .O(N__20847),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__4675 (
            .O(N__20844),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__4674 (
            .O(N__20841),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__4673 (
            .O(N__20838),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__4672 (
            .O(N__20835),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__4671 (
            .O(N__20832),
            .I(bfn_11_26_0_));
    InMux I__4670 (
            .O(N__20829),
            .I(N__20825));
    InMux I__4669 (
            .O(N__20828),
            .I(N__20822));
    LocalMux I__4668 (
            .O(N__20825),
            .I(N__20817));
    LocalMux I__4667 (
            .O(N__20822),
            .I(N__20817));
    Span4Mux_v I__4666 (
            .O(N__20817),
            .I(N__20812));
    InMux I__4665 (
            .O(N__20816),
            .I(N__20809));
    CascadeMux I__4664 (
            .O(N__20815),
            .I(N__20806));
    Span4Mux_h I__4663 (
            .O(N__20812),
            .I(N__20801));
    LocalMux I__4662 (
            .O(N__20809),
            .I(N__20801));
    InMux I__4661 (
            .O(N__20806),
            .I(N__20798));
    Odrv4 I__4660 (
            .O(N__20801),
            .I(\ppm_encoder_1.N_443 ));
    LocalMux I__4659 (
            .O(N__20798),
            .I(\ppm_encoder_1.N_443 ));
    CascadeMux I__4658 (
            .O(N__20793),
            .I(N__20790));
    InMux I__4657 (
            .O(N__20790),
            .I(N__20787));
    LocalMux I__4656 (
            .O(N__20787),
            .I(N__20784));
    Span12Mux_s8_v I__4655 (
            .O(N__20784),
            .I(N__20781));
    Odrv12 I__4654 (
            .O(N__20781),
            .I(\ppm_encoder_1.pulses2count_9_0_2_1 ));
    InMux I__4653 (
            .O(N__20778),
            .I(N__20772));
    InMux I__4652 (
            .O(N__20777),
            .I(N__20772));
    LocalMux I__4651 (
            .O(N__20772),
            .I(N__20767));
    InMux I__4650 (
            .O(N__20771),
            .I(N__20762));
    InMux I__4649 (
            .O(N__20770),
            .I(N__20762));
    Odrv4 I__4648 (
            .O(N__20767),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    LocalMux I__4647 (
            .O(N__20762),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    InMux I__4646 (
            .O(N__20757),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__4645 (
            .O(N__20754),
            .I(N__20749));
    InMux I__4644 (
            .O(N__20753),
            .I(N__20746));
    InMux I__4643 (
            .O(N__20752),
            .I(N__20743));
    LocalMux I__4642 (
            .O(N__20749),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__4641 (
            .O(N__20746),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__4640 (
            .O(N__20743),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__4639 (
            .O(N__20736),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__4638 (
            .O(N__20733),
            .I(N__20728));
    InMux I__4637 (
            .O(N__20732),
            .I(N__20725));
    InMux I__4636 (
            .O(N__20731),
            .I(N__20722));
    LocalMux I__4635 (
            .O(N__20728),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__4634 (
            .O(N__20725),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__4633 (
            .O(N__20722),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__4632 (
            .O(N__20715),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__4631 (
            .O(N__20712),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__4630 (
            .O(N__20709),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__4629 (
            .O(N__20706),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__4628 (
            .O(N__20703),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__4627 (
            .O(N__20700),
            .I(N__20697));
    LocalMux I__4626 (
            .O(N__20697),
            .I(N__20694));
    Span12Mux_h I__4625 (
            .O(N__20694),
            .I(N__20691));
    Odrv12 I__4624 (
            .O(N__20691),
            .I(\ppm_encoder_1.N_369 ));
    CascadeMux I__4623 (
            .O(N__20688),
            .I(\ppm_encoder_1.N_371_cascade_ ));
    InMux I__4622 (
            .O(N__20685),
            .I(N__20682));
    LocalMux I__4621 (
            .O(N__20682),
            .I(N__20679));
    Span4Mux_v I__4620 (
            .O(N__20679),
            .I(N__20676));
    Span4Mux_v I__4619 (
            .O(N__20676),
            .I(N__20672));
    InMux I__4618 (
            .O(N__20675),
            .I(N__20669));
    Odrv4 I__4617 (
            .O(N__20672),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    LocalMux I__4616 (
            .O(N__20669),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    InMux I__4615 (
            .O(N__20664),
            .I(N__20660));
    CascadeMux I__4614 (
            .O(N__20663),
            .I(N__20656));
    LocalMux I__4613 (
            .O(N__20660),
            .I(N__20653));
    InMux I__4612 (
            .O(N__20659),
            .I(N__20650));
    InMux I__4611 (
            .O(N__20656),
            .I(N__20647));
    Span4Mux_v I__4610 (
            .O(N__20653),
            .I(N__20644));
    LocalMux I__4609 (
            .O(N__20650),
            .I(N__20641));
    LocalMux I__4608 (
            .O(N__20647),
            .I(N__20638));
    Span4Mux_h I__4607 (
            .O(N__20644),
            .I(N__20635));
    Span4Mux_h I__4606 (
            .O(N__20641),
            .I(N__20632));
    Odrv4 I__4605 (
            .O(N__20638),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__4604 (
            .O(N__20635),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__4603 (
            .O(N__20632),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__4602 (
            .O(N__20625),
            .I(N__20622));
    LocalMux I__4601 (
            .O(N__20622),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__4600 (
            .O(N__20619),
            .I(N__20616));
    LocalMux I__4599 (
            .O(N__20616),
            .I(N__20611));
    InMux I__4598 (
            .O(N__20615),
            .I(N__20608));
    InMux I__4597 (
            .O(N__20614),
            .I(N__20605));
    Span4Mux_v I__4596 (
            .O(N__20611),
            .I(N__20602));
    LocalMux I__4595 (
            .O(N__20608),
            .I(N__20599));
    LocalMux I__4594 (
            .O(N__20605),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__4593 (
            .O(N__20602),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv12 I__4592 (
            .O(N__20599),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__4591 (
            .O(N__20592),
            .I(N__20588));
    CascadeMux I__4590 (
            .O(N__20591),
            .I(N__20583));
    LocalMux I__4589 (
            .O(N__20588),
            .I(N__20580));
    InMux I__4588 (
            .O(N__20587),
            .I(N__20577));
    InMux I__4587 (
            .O(N__20586),
            .I(N__20574));
    InMux I__4586 (
            .O(N__20583),
            .I(N__20571));
    Span4Mux_h I__4585 (
            .O(N__20580),
            .I(N__20562));
    LocalMux I__4584 (
            .O(N__20577),
            .I(N__20562));
    LocalMux I__4583 (
            .O(N__20574),
            .I(N__20562));
    LocalMux I__4582 (
            .O(N__20571),
            .I(N__20562));
    Span4Mux_v I__4581 (
            .O(N__20562),
            .I(N__20559));
    Odrv4 I__4580 (
            .O(N__20559),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__4579 (
            .O(N__20556),
            .I(N__20553));
    LocalMux I__4578 (
            .O(N__20553),
            .I(N__20550));
    Odrv4 I__4577 (
            .O(N__20550),
            .I(\ppm_encoder_1.N_360 ));
    CascadeMux I__4576 (
            .O(N__20547),
            .I(N__20544));
    InMux I__4575 (
            .O(N__20544),
            .I(N__20541));
    LocalMux I__4574 (
            .O(N__20541),
            .I(N__20536));
    InMux I__4573 (
            .O(N__20540),
            .I(N__20533));
    CascadeMux I__4572 (
            .O(N__20539),
            .I(N__20528));
    Span4Mux_v I__4571 (
            .O(N__20536),
            .I(N__20525));
    LocalMux I__4570 (
            .O(N__20533),
            .I(N__20522));
    InMux I__4569 (
            .O(N__20532),
            .I(N__20515));
    InMux I__4568 (
            .O(N__20531),
            .I(N__20515));
    InMux I__4567 (
            .O(N__20528),
            .I(N__20515));
    Span4Mux_h I__4566 (
            .O(N__20525),
            .I(N__20512));
    Span4Mux_h I__4565 (
            .O(N__20522),
            .I(N__20507));
    LocalMux I__4564 (
            .O(N__20515),
            .I(N__20507));
    Odrv4 I__4563 (
            .O(N__20512),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__4562 (
            .O(N__20507),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    CascadeMux I__4561 (
            .O(N__20502),
            .I(N__20498));
    InMux I__4560 (
            .O(N__20501),
            .I(N__20495));
    InMux I__4559 (
            .O(N__20498),
            .I(N__20492));
    LocalMux I__4558 (
            .O(N__20495),
            .I(\ppm_encoder_1.pulses2count_9_0_0_3 ));
    LocalMux I__4557 (
            .O(N__20492),
            .I(\ppm_encoder_1.pulses2count_9_0_0_3 ));
    InMux I__4556 (
            .O(N__20487),
            .I(N__20484));
    LocalMux I__4555 (
            .O(N__20484),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CascadeMux I__4554 (
            .O(N__20481),
            .I(N__20478));
    InMux I__4553 (
            .O(N__20478),
            .I(N__20475));
    LocalMux I__4552 (
            .O(N__20475),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__4551 (
            .O(N__20472),
            .I(N__20469));
    LocalMux I__4550 (
            .O(N__20469),
            .I(\ppm_encoder_1.N_365 ));
    InMux I__4549 (
            .O(N__20466),
            .I(N__20463));
    LocalMux I__4548 (
            .O(N__20463),
            .I(\ppm_encoder_1.init_pulses_RNILB4MZ0Z_0 ));
    InMux I__4547 (
            .O(N__20460),
            .I(N__20455));
    InMux I__4546 (
            .O(N__20459),
            .I(N__20450));
    InMux I__4545 (
            .O(N__20458),
            .I(N__20450));
    LocalMux I__4544 (
            .O(N__20455),
            .I(N__20444));
    LocalMux I__4543 (
            .O(N__20450),
            .I(N__20444));
    InMux I__4542 (
            .O(N__20449),
            .I(N__20441));
    Span4Mux_h I__4541 (
            .O(N__20444),
            .I(N__20435));
    LocalMux I__4540 (
            .O(N__20441),
            .I(N__20435));
    CascadeMux I__4539 (
            .O(N__20440),
            .I(N__20432));
    Span4Mux_v I__4538 (
            .O(N__20435),
            .I(N__20429));
    InMux I__4537 (
            .O(N__20432),
            .I(N__20426));
    Odrv4 I__4536 (
            .O(N__20429),
            .I(\ppm_encoder_1.N_247_i_i ));
    LocalMux I__4535 (
            .O(N__20426),
            .I(\ppm_encoder_1.N_247_i_i ));
    CascadeMux I__4534 (
            .O(N__20421),
            .I(N__20415));
    InMux I__4533 (
            .O(N__20420),
            .I(N__20409));
    InMux I__4532 (
            .O(N__20419),
            .I(N__20409));
    InMux I__4531 (
            .O(N__20418),
            .I(N__20403));
    InMux I__4530 (
            .O(N__20415),
            .I(N__20400));
    InMux I__4529 (
            .O(N__20414),
            .I(N__20392));
    LocalMux I__4528 (
            .O(N__20409),
            .I(N__20388));
    InMux I__4527 (
            .O(N__20408),
            .I(N__20381));
    InMux I__4526 (
            .O(N__20407),
            .I(N__20381));
    InMux I__4525 (
            .O(N__20406),
            .I(N__20381));
    LocalMux I__4524 (
            .O(N__20403),
            .I(N__20376));
    LocalMux I__4523 (
            .O(N__20400),
            .I(N__20376));
    InMux I__4522 (
            .O(N__20399),
            .I(N__20371));
    InMux I__4521 (
            .O(N__20398),
            .I(N__20371));
    InMux I__4520 (
            .O(N__20397),
            .I(N__20368));
    InMux I__4519 (
            .O(N__20396),
            .I(N__20363));
    InMux I__4518 (
            .O(N__20395),
            .I(N__20363));
    LocalMux I__4517 (
            .O(N__20392),
            .I(N__20359));
    InMux I__4516 (
            .O(N__20391),
            .I(N__20356));
    Span4Mux_v I__4515 (
            .O(N__20388),
            .I(N__20351));
    LocalMux I__4514 (
            .O(N__20381),
            .I(N__20351));
    Span4Mux_v I__4513 (
            .O(N__20376),
            .I(N__20337));
    LocalMux I__4512 (
            .O(N__20371),
            .I(N__20337));
    LocalMux I__4511 (
            .O(N__20368),
            .I(N__20334));
    LocalMux I__4510 (
            .O(N__20363),
            .I(N__20331));
    InMux I__4509 (
            .O(N__20362),
            .I(N__20328));
    Span4Mux_v I__4508 (
            .O(N__20359),
            .I(N__20321));
    LocalMux I__4507 (
            .O(N__20356),
            .I(N__20321));
    Span4Mux_v I__4506 (
            .O(N__20351),
            .I(N__20321));
    InMux I__4505 (
            .O(N__20350),
            .I(N__20316));
    InMux I__4504 (
            .O(N__20349),
            .I(N__20316));
    InMux I__4503 (
            .O(N__20348),
            .I(N__20311));
    InMux I__4502 (
            .O(N__20347),
            .I(N__20311));
    InMux I__4501 (
            .O(N__20346),
            .I(N__20302));
    InMux I__4500 (
            .O(N__20345),
            .I(N__20302));
    InMux I__4499 (
            .O(N__20344),
            .I(N__20302));
    InMux I__4498 (
            .O(N__20343),
            .I(N__20302));
    InMux I__4497 (
            .O(N__20342),
            .I(N__20299));
    Span4Mux_h I__4496 (
            .O(N__20337),
            .I(N__20294));
    Span4Mux_v I__4495 (
            .O(N__20334),
            .I(N__20294));
    Span4Mux_h I__4494 (
            .O(N__20331),
            .I(N__20287));
    LocalMux I__4493 (
            .O(N__20328),
            .I(N__20287));
    Span4Mux_h I__4492 (
            .O(N__20321),
            .I(N__20287));
    LocalMux I__4491 (
            .O(N__20316),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__4490 (
            .O(N__20311),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__4489 (
            .O(N__20302),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__4488 (
            .O(N__20299),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__4487 (
            .O(N__20294),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__4486 (
            .O(N__20287),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    CascadeMux I__4485 (
            .O(N__20274),
            .I(N__20269));
    CascadeMux I__4484 (
            .O(N__20273),
            .I(N__20266));
    InMux I__4483 (
            .O(N__20272),
            .I(N__20263));
    InMux I__4482 (
            .O(N__20269),
            .I(N__20258));
    InMux I__4481 (
            .O(N__20266),
            .I(N__20258));
    LocalMux I__4480 (
            .O(N__20263),
            .I(N__20250));
    LocalMux I__4479 (
            .O(N__20258),
            .I(N__20250));
    InMux I__4478 (
            .O(N__20257),
            .I(N__20247));
    InMux I__4477 (
            .O(N__20256),
            .I(N__20244));
    InMux I__4476 (
            .O(N__20255),
            .I(N__20237));
    Span4Mux_v I__4475 (
            .O(N__20250),
            .I(N__20232));
    LocalMux I__4474 (
            .O(N__20247),
            .I(N__20229));
    LocalMux I__4473 (
            .O(N__20244),
            .I(N__20226));
    InMux I__4472 (
            .O(N__20243),
            .I(N__20223));
    InMux I__4471 (
            .O(N__20242),
            .I(N__20219));
    InMux I__4470 (
            .O(N__20241),
            .I(N__20214));
    InMux I__4469 (
            .O(N__20240),
            .I(N__20211));
    LocalMux I__4468 (
            .O(N__20237),
            .I(N__20208));
    InMux I__4467 (
            .O(N__20236),
            .I(N__20203));
    InMux I__4466 (
            .O(N__20235),
            .I(N__20203));
    Span4Mux_h I__4465 (
            .O(N__20232),
            .I(N__20200));
    Span4Mux_h I__4464 (
            .O(N__20229),
            .I(N__20193));
    Span4Mux_h I__4463 (
            .O(N__20226),
            .I(N__20193));
    LocalMux I__4462 (
            .O(N__20223),
            .I(N__20193));
    InMux I__4461 (
            .O(N__20222),
            .I(N__20190));
    LocalMux I__4460 (
            .O(N__20219),
            .I(N__20187));
    InMux I__4459 (
            .O(N__20218),
            .I(N__20182));
    InMux I__4458 (
            .O(N__20217),
            .I(N__20182));
    LocalMux I__4457 (
            .O(N__20214),
            .I(N__20177));
    LocalMux I__4456 (
            .O(N__20211),
            .I(N__20177));
    Odrv4 I__4455 (
            .O(N__20208),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    LocalMux I__4454 (
            .O(N__20203),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    Odrv4 I__4453 (
            .O(N__20200),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    Odrv4 I__4452 (
            .O(N__20193),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    LocalMux I__4451 (
            .O(N__20190),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    Odrv12 I__4450 (
            .O(N__20187),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    LocalMux I__4449 (
            .O(N__20182),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    Odrv4 I__4448 (
            .O(N__20177),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ));
    InMux I__4447 (
            .O(N__20160),
            .I(N__20152));
    InMux I__4446 (
            .O(N__20159),
            .I(N__20152));
    InMux I__4445 (
            .O(N__20158),
            .I(N__20147));
    InMux I__4444 (
            .O(N__20157),
            .I(N__20144));
    LocalMux I__4443 (
            .O(N__20152),
            .I(N__20140));
    InMux I__4442 (
            .O(N__20151),
            .I(N__20137));
    InMux I__4441 (
            .O(N__20150),
            .I(N__20134));
    LocalMux I__4440 (
            .O(N__20147),
            .I(N__20129));
    LocalMux I__4439 (
            .O(N__20144),
            .I(N__20124));
    InMux I__4438 (
            .O(N__20143),
            .I(N__20121));
    Span4Mux_h I__4437 (
            .O(N__20140),
            .I(N__20116));
    LocalMux I__4436 (
            .O(N__20137),
            .I(N__20110));
    LocalMux I__4435 (
            .O(N__20134),
            .I(N__20110));
    InMux I__4434 (
            .O(N__20133),
            .I(N__20105));
    InMux I__4433 (
            .O(N__20132),
            .I(N__20105));
    Span4Mux_h I__4432 (
            .O(N__20129),
            .I(N__20100));
    InMux I__4431 (
            .O(N__20128),
            .I(N__20097));
    InMux I__4430 (
            .O(N__20127),
            .I(N__20094));
    Span4Mux_h I__4429 (
            .O(N__20124),
            .I(N__20091));
    LocalMux I__4428 (
            .O(N__20121),
            .I(N__20088));
    InMux I__4427 (
            .O(N__20120),
            .I(N__20083));
    InMux I__4426 (
            .O(N__20119),
            .I(N__20083));
    Span4Mux_v I__4425 (
            .O(N__20116),
            .I(N__20080));
    InMux I__4424 (
            .O(N__20115),
            .I(N__20077));
    Span4Mux_h I__4423 (
            .O(N__20110),
            .I(N__20072));
    LocalMux I__4422 (
            .O(N__20105),
            .I(N__20072));
    InMux I__4421 (
            .O(N__20104),
            .I(N__20067));
    InMux I__4420 (
            .O(N__20103),
            .I(N__20067));
    Span4Mux_v I__4419 (
            .O(N__20100),
            .I(N__20060));
    LocalMux I__4418 (
            .O(N__20097),
            .I(N__20060));
    LocalMux I__4417 (
            .O(N__20094),
            .I(N__20060));
    Odrv4 I__4416 (
            .O(N__20091),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    Odrv4 I__4415 (
            .O(N__20088),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    LocalMux I__4414 (
            .O(N__20083),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    Odrv4 I__4413 (
            .O(N__20080),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    LocalMux I__4412 (
            .O(N__20077),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    Odrv4 I__4411 (
            .O(N__20072),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    LocalMux I__4410 (
            .O(N__20067),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    Odrv4 I__4409 (
            .O(N__20060),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ));
    CascadeMux I__4408 (
            .O(N__20043),
            .I(N__20040));
    InMux I__4407 (
            .O(N__20040),
            .I(N__20036));
    CascadeMux I__4406 (
            .O(N__20039),
            .I(N__20033));
    LocalMux I__4405 (
            .O(N__20036),
            .I(N__20029));
    InMux I__4404 (
            .O(N__20033),
            .I(N__20026));
    InMux I__4403 (
            .O(N__20032),
            .I(N__20023));
    Span4Mux_v I__4402 (
            .O(N__20029),
            .I(N__20018));
    LocalMux I__4401 (
            .O(N__20026),
            .I(N__20018));
    LocalMux I__4400 (
            .O(N__20023),
            .I(N__20015));
    Span4Mux_h I__4399 (
            .O(N__20018),
            .I(N__20011));
    Span4Mux_h I__4398 (
            .O(N__20015),
            .I(N__20008));
    InMux I__4397 (
            .O(N__20014),
            .I(N__20005));
    Span4Mux_v I__4396 (
            .O(N__20011),
            .I(N__20002));
    Odrv4 I__4395 (
            .O(N__20008),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__4394 (
            .O(N__20005),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    Odrv4 I__4393 (
            .O(N__20002),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    CascadeMux I__4392 (
            .O(N__19995),
            .I(\ppm_encoder_1.N_441_cascade_ ));
    InMux I__4391 (
            .O(N__19992),
            .I(N__19989));
    LocalMux I__4390 (
            .O(N__19989),
            .I(N__19985));
    CascadeMux I__4389 (
            .O(N__19988),
            .I(N__19981));
    Span4Mux_h I__4388 (
            .O(N__19985),
            .I(N__19978));
    InMux I__4387 (
            .O(N__19984),
            .I(N__19973));
    InMux I__4386 (
            .O(N__19981),
            .I(N__19973));
    Odrv4 I__4385 (
            .O(N__19978),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__4384 (
            .O(N__19973),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    InMux I__4383 (
            .O(N__19968),
            .I(N__19965));
    LocalMux I__4382 (
            .O(N__19965),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_18 ));
    InMux I__4381 (
            .O(N__19962),
            .I(N__19959));
    LocalMux I__4380 (
            .O(N__19959),
            .I(N__19955));
    CascadeMux I__4379 (
            .O(N__19958),
            .I(N__19951));
    Span4Mux_h I__4378 (
            .O(N__19955),
            .I(N__19948));
    InMux I__4377 (
            .O(N__19954),
            .I(N__19945));
    InMux I__4376 (
            .O(N__19951),
            .I(N__19942));
    Span4Mux_h I__4375 (
            .O(N__19948),
            .I(N__19937));
    LocalMux I__4374 (
            .O(N__19945),
            .I(N__19937));
    LocalMux I__4373 (
            .O(N__19942),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__4372 (
            .O(N__19937),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__4371 (
            .O(N__19932),
            .I(N__19928));
    CascadeMux I__4370 (
            .O(N__19931),
            .I(N__19924));
    LocalMux I__4369 (
            .O(N__19928),
            .I(N__19921));
    InMux I__4368 (
            .O(N__19927),
            .I(N__19918));
    InMux I__4367 (
            .O(N__19924),
            .I(N__19915));
    Span12Mux_s4_v I__4366 (
            .O(N__19921),
            .I(N__19912));
    LocalMux I__4365 (
            .O(N__19918),
            .I(N__19909));
    LocalMux I__4364 (
            .O(N__19915),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv12 I__4363 (
            .O(N__19912),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__4362 (
            .O(N__19909),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__4361 (
            .O(N__19902),
            .I(N__19899));
    LocalMux I__4360 (
            .O(N__19899),
            .I(N__19896));
    Span4Mux_h I__4359 (
            .O(N__19896),
            .I(N__19893));
    Odrv4 I__4358 (
            .O(N__19893),
            .I(\ppm_encoder_1.N_383 ));
    CascadeMux I__4357 (
            .O(N__19890),
            .I(\ppm_encoder_1.N_385_cascade_ ));
    InMux I__4356 (
            .O(N__19887),
            .I(N__19884));
    LocalMux I__4355 (
            .O(N__19884),
            .I(N__19881));
    Span4Mux_v I__4354 (
            .O(N__19881),
            .I(N__19878));
    Span4Mux_v I__4353 (
            .O(N__19878),
            .I(N__19874));
    InMux I__4352 (
            .O(N__19877),
            .I(N__19871));
    Odrv4 I__4351 (
            .O(N__19874),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    LocalMux I__4350 (
            .O(N__19871),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    CascadeMux I__4349 (
            .O(N__19866),
            .I(N__19863));
    InMux I__4348 (
            .O(N__19863),
            .I(N__19855));
    InMux I__4347 (
            .O(N__19862),
            .I(N__19852));
    InMux I__4346 (
            .O(N__19861),
            .I(N__19849));
    InMux I__4345 (
            .O(N__19860),
            .I(N__19844));
    InMux I__4344 (
            .O(N__19859),
            .I(N__19844));
    InMux I__4343 (
            .O(N__19858),
            .I(N__19841));
    LocalMux I__4342 (
            .O(N__19855),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__4341 (
            .O(N__19852),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__4340 (
            .O(N__19849),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__4339 (
            .O(N__19844),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__4338 (
            .O(N__19841),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__4337 (
            .O(N__19830),
            .I(N__19827));
    LocalMux I__4336 (
            .O(N__19827),
            .I(N__19823));
    CascadeMux I__4335 (
            .O(N__19826),
            .I(N__19812));
    Span4Mux_h I__4334 (
            .O(N__19823),
            .I(N__19809));
    InMux I__4333 (
            .O(N__19822),
            .I(N__19806));
    InMux I__4332 (
            .O(N__19821),
            .I(N__19801));
    InMux I__4331 (
            .O(N__19820),
            .I(N__19801));
    InMux I__4330 (
            .O(N__19819),
            .I(N__19798));
    InMux I__4329 (
            .O(N__19818),
            .I(N__19795));
    InMux I__4328 (
            .O(N__19817),
            .I(N__19790));
    InMux I__4327 (
            .O(N__19816),
            .I(N__19790));
    InMux I__4326 (
            .O(N__19815),
            .I(N__19785));
    InMux I__4325 (
            .O(N__19812),
            .I(N__19785));
    Odrv4 I__4324 (
            .O(N__19809),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4323 (
            .O(N__19806),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4322 (
            .O(N__19801),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4321 (
            .O(N__19798),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4320 (
            .O(N__19795),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4319 (
            .O(N__19790),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__4318 (
            .O(N__19785),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__4317 (
            .O(N__19770),
            .I(N__19762));
    InMux I__4316 (
            .O(N__19769),
            .I(N__19759));
    CascadeMux I__4315 (
            .O(N__19768),
            .I(N__19756));
    CascadeMux I__4314 (
            .O(N__19767),
            .I(N__19753));
    CascadeMux I__4313 (
            .O(N__19766),
            .I(N__19750));
    CascadeMux I__4312 (
            .O(N__19765),
            .I(N__19747));
    LocalMux I__4311 (
            .O(N__19762),
            .I(N__19742));
    LocalMux I__4310 (
            .O(N__19759),
            .I(N__19739));
    InMux I__4309 (
            .O(N__19756),
            .I(N__19730));
    InMux I__4308 (
            .O(N__19753),
            .I(N__19730));
    InMux I__4307 (
            .O(N__19750),
            .I(N__19730));
    InMux I__4306 (
            .O(N__19747),
            .I(N__19730));
    InMux I__4305 (
            .O(N__19746),
            .I(N__19727));
    InMux I__4304 (
            .O(N__19745),
            .I(N__19724));
    Span4Mux_h I__4303 (
            .O(N__19742),
            .I(N__19715));
    Span4Mux_h I__4302 (
            .O(N__19739),
            .I(N__19715));
    LocalMux I__4301 (
            .O(N__19730),
            .I(N__19715));
    LocalMux I__4300 (
            .O(N__19727),
            .I(N__19715));
    LocalMux I__4299 (
            .O(N__19724),
            .I(N__19710));
    Span4Mux_v I__4298 (
            .O(N__19715),
            .I(N__19707));
    CascadeMux I__4297 (
            .O(N__19714),
            .I(N__19702));
    InMux I__4296 (
            .O(N__19713),
            .I(N__19698));
    Span4Mux_v I__4295 (
            .O(N__19710),
            .I(N__19695));
    Span4Mux_h I__4294 (
            .O(N__19707),
            .I(N__19692));
    CascadeMux I__4293 (
            .O(N__19706),
            .I(N__19683));
    InMux I__4292 (
            .O(N__19705),
            .I(N__19680));
    InMux I__4291 (
            .O(N__19702),
            .I(N__19675));
    InMux I__4290 (
            .O(N__19701),
            .I(N__19675));
    LocalMux I__4289 (
            .O(N__19698),
            .I(N__19672));
    Span4Mux_h I__4288 (
            .O(N__19695),
            .I(N__19669));
    Span4Mux_h I__4287 (
            .O(N__19692),
            .I(N__19666));
    InMux I__4286 (
            .O(N__19691),
            .I(N__19655));
    InMux I__4285 (
            .O(N__19690),
            .I(N__19655));
    InMux I__4284 (
            .O(N__19689),
            .I(N__19655));
    InMux I__4283 (
            .O(N__19688),
            .I(N__19655));
    InMux I__4282 (
            .O(N__19687),
            .I(N__19655));
    InMux I__4281 (
            .O(N__19686),
            .I(N__19650));
    InMux I__4280 (
            .O(N__19683),
            .I(N__19650));
    LocalMux I__4279 (
            .O(N__19680),
            .I(N__19643));
    LocalMux I__4278 (
            .O(N__19675),
            .I(N__19643));
    Span4Mux_h I__4277 (
            .O(N__19672),
            .I(N__19643));
    Odrv4 I__4276 (
            .O(N__19669),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv4 I__4275 (
            .O(N__19666),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    LocalMux I__4274 (
            .O(N__19655),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    LocalMux I__4273 (
            .O(N__19650),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv4 I__4272 (
            .O(N__19643),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    CascadeMux I__4271 (
            .O(N__19632),
            .I(N__19627));
    InMux I__4270 (
            .O(N__19631),
            .I(N__19615));
    InMux I__4269 (
            .O(N__19630),
            .I(N__19615));
    InMux I__4268 (
            .O(N__19627),
            .I(N__19610));
    InMux I__4267 (
            .O(N__19626),
            .I(N__19610));
    InMux I__4266 (
            .O(N__19625),
            .I(N__19607));
    InMux I__4265 (
            .O(N__19624),
            .I(N__19604));
    InMux I__4264 (
            .O(N__19623),
            .I(N__19598));
    InMux I__4263 (
            .O(N__19622),
            .I(N__19598));
    InMux I__4262 (
            .O(N__19621),
            .I(N__19594));
    CascadeMux I__4261 (
            .O(N__19620),
            .I(N__19588));
    LocalMux I__4260 (
            .O(N__19615),
            .I(N__19582));
    LocalMux I__4259 (
            .O(N__19610),
            .I(N__19582));
    LocalMux I__4258 (
            .O(N__19607),
            .I(N__19577));
    LocalMux I__4257 (
            .O(N__19604),
            .I(N__19577));
    InMux I__4256 (
            .O(N__19603),
            .I(N__19574));
    LocalMux I__4255 (
            .O(N__19598),
            .I(N__19571));
    InMux I__4254 (
            .O(N__19597),
            .I(N__19568));
    LocalMux I__4253 (
            .O(N__19594),
            .I(N__19565));
    InMux I__4252 (
            .O(N__19593),
            .I(N__19558));
    InMux I__4251 (
            .O(N__19592),
            .I(N__19558));
    InMux I__4250 (
            .O(N__19591),
            .I(N__19558));
    InMux I__4249 (
            .O(N__19588),
            .I(N__19555));
    InMux I__4248 (
            .O(N__19587),
            .I(N__19548));
    Span4Mux_v I__4247 (
            .O(N__19582),
            .I(N__19541));
    Span4Mux_v I__4246 (
            .O(N__19577),
            .I(N__19541));
    LocalMux I__4245 (
            .O(N__19574),
            .I(N__19541));
    Span4Mux_v I__4244 (
            .O(N__19571),
            .I(N__19533));
    LocalMux I__4243 (
            .O(N__19568),
            .I(N__19533));
    Span4Mux_v I__4242 (
            .O(N__19565),
            .I(N__19526));
    LocalMux I__4241 (
            .O(N__19558),
            .I(N__19526));
    LocalMux I__4240 (
            .O(N__19555),
            .I(N__19526));
    InMux I__4239 (
            .O(N__19554),
            .I(N__19521));
    InMux I__4238 (
            .O(N__19553),
            .I(N__19521));
    InMux I__4237 (
            .O(N__19552),
            .I(N__19516));
    InMux I__4236 (
            .O(N__19551),
            .I(N__19516));
    LocalMux I__4235 (
            .O(N__19548),
            .I(N__19513));
    Span4Mux_h I__4234 (
            .O(N__19541),
            .I(N__19510));
    InMux I__4233 (
            .O(N__19540),
            .I(N__19507));
    InMux I__4232 (
            .O(N__19539),
            .I(N__19502));
    InMux I__4231 (
            .O(N__19538),
            .I(N__19502));
    Span4Mux_h I__4230 (
            .O(N__19533),
            .I(N__19497));
    Span4Mux_h I__4229 (
            .O(N__19526),
            .I(N__19497));
    LocalMux I__4228 (
            .O(N__19521),
            .I(N__19492));
    LocalMux I__4227 (
            .O(N__19516),
            .I(N__19492));
    Odrv4 I__4226 (
            .O(N__19513),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__4225 (
            .O(N__19510),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__4224 (
            .O(N__19507),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__4223 (
            .O(N__19502),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__4222 (
            .O(N__19497),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv12 I__4221 (
            .O(N__19492),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    CascadeMux I__4220 (
            .O(N__19479),
            .I(N__19476));
    InMux I__4219 (
            .O(N__19476),
            .I(N__19472));
    CascadeMux I__4218 (
            .O(N__19475),
            .I(N__19468));
    LocalMux I__4217 (
            .O(N__19472),
            .I(N__19464));
    InMux I__4216 (
            .O(N__19471),
            .I(N__19461));
    InMux I__4215 (
            .O(N__19468),
            .I(N__19458));
    InMux I__4214 (
            .O(N__19467),
            .I(N__19455));
    Span4Mux_v I__4213 (
            .O(N__19464),
            .I(N__19452));
    LocalMux I__4212 (
            .O(N__19461),
            .I(N__19449));
    LocalMux I__4211 (
            .O(N__19458),
            .I(N__19444));
    LocalMux I__4210 (
            .O(N__19455),
            .I(N__19444));
    Span4Mux_s2_v I__4209 (
            .O(N__19452),
            .I(N__19441));
    Span4Mux_h I__4208 (
            .O(N__19449),
            .I(N__19436));
    Span4Mux_v I__4207 (
            .O(N__19444),
            .I(N__19436));
    Odrv4 I__4206 (
            .O(N__19441),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__4205 (
            .O(N__19436),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__4204 (
            .O(N__19431),
            .I(N__19428));
    LocalMux I__4203 (
            .O(N__19428),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    CascadeMux I__4202 (
            .O(N__19425),
            .I(N__19421));
    InMux I__4201 (
            .O(N__19424),
            .I(N__19418));
    InMux I__4200 (
            .O(N__19421),
            .I(N__19415));
    LocalMux I__4199 (
            .O(N__19418),
            .I(\ppm_encoder_1.PPM_STATE_fastZ0Z_0 ));
    LocalMux I__4198 (
            .O(N__19415),
            .I(\ppm_encoder_1.PPM_STATE_fastZ0Z_0 ));
    InMux I__4197 (
            .O(N__19410),
            .I(N__19407));
    LocalMux I__4196 (
            .O(N__19407),
            .I(N__19402));
    InMux I__4195 (
            .O(N__19406),
            .I(N__19399));
    CascadeMux I__4194 (
            .O(N__19405),
            .I(N__19396));
    Span4Mux_v I__4193 (
            .O(N__19402),
            .I(N__19393));
    LocalMux I__4192 (
            .O(N__19399),
            .I(N__19390));
    InMux I__4191 (
            .O(N__19396),
            .I(N__19387));
    Span4Mux_h I__4190 (
            .O(N__19393),
            .I(N__19384));
    Span4Mux_h I__4189 (
            .O(N__19390),
            .I(N__19381));
    LocalMux I__4188 (
            .O(N__19387),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    Odrv4 I__4187 (
            .O(N__19384),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    Odrv4 I__4186 (
            .O(N__19381),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__4185 (
            .O(N__19374),
            .I(N__19370));
    CascadeMux I__4184 (
            .O(N__19373),
            .I(N__19367));
    LocalMux I__4183 (
            .O(N__19370),
            .I(N__19364));
    InMux I__4182 (
            .O(N__19367),
            .I(N__19361));
    Span4Mux_v I__4181 (
            .O(N__19364),
            .I(N__19357));
    LocalMux I__4180 (
            .O(N__19361),
            .I(N__19354));
    InMux I__4179 (
            .O(N__19360),
            .I(N__19351));
    Span4Mux_h I__4178 (
            .O(N__19357),
            .I(N__19348));
    Span4Mux_h I__4177 (
            .O(N__19354),
            .I(N__19345));
    LocalMux I__4176 (
            .O(N__19351),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__4175 (
            .O(N__19348),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__4174 (
            .O(N__19345),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    CascadeMux I__4173 (
            .O(N__19338),
            .I(N__19333));
    CascadeMux I__4172 (
            .O(N__19337),
            .I(N__19330));
    InMux I__4171 (
            .O(N__19336),
            .I(N__19325));
    InMux I__4170 (
            .O(N__19333),
            .I(N__19325));
    InMux I__4169 (
            .O(N__19330),
            .I(N__19322));
    LocalMux I__4168 (
            .O(N__19325),
            .I(N__19319));
    LocalMux I__4167 (
            .O(N__19322),
            .I(N__19315));
    Span4Mux_h I__4166 (
            .O(N__19319),
            .I(N__19312));
    InMux I__4165 (
            .O(N__19318),
            .I(N__19309));
    Span4Mux_h I__4164 (
            .O(N__19315),
            .I(N__19306));
    Span4Mux_v I__4163 (
            .O(N__19312),
            .I(N__19303));
    LocalMux I__4162 (
            .O(N__19309),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    Odrv4 I__4161 (
            .O(N__19306),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    Odrv4 I__4160 (
            .O(N__19303),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    CascadeMux I__4159 (
            .O(N__19296),
            .I(N__19292));
    InMux I__4158 (
            .O(N__19295),
            .I(N__19289));
    InMux I__4157 (
            .O(N__19292),
            .I(N__19286));
    LocalMux I__4156 (
            .O(N__19289),
            .I(N__19283));
    LocalMux I__4155 (
            .O(N__19286),
            .I(N__19280));
    Span4Mux_h I__4154 (
            .O(N__19283),
            .I(N__19277));
    Span4Mux_v I__4153 (
            .O(N__19280),
            .I(N__19274));
    Span4Mux_h I__4152 (
            .O(N__19277),
            .I(N__19271));
    Odrv4 I__4151 (
            .O(N__19274),
            .I(\ppm_encoder_1.N_258_i_i ));
    Odrv4 I__4150 (
            .O(N__19271),
            .I(\ppm_encoder_1.N_258_i_i ));
    CascadeMux I__4149 (
            .O(N__19266),
            .I(N__19263));
    InMux I__4148 (
            .O(N__19263),
            .I(N__19259));
    InMux I__4147 (
            .O(N__19262),
            .I(N__19256));
    LocalMux I__4146 (
            .O(N__19259),
            .I(N__19253));
    LocalMux I__4145 (
            .O(N__19256),
            .I(N__19250));
    Span4Mux_h I__4144 (
            .O(N__19253),
            .I(N__19247));
    Span4Mux_h I__4143 (
            .O(N__19250),
            .I(N__19244));
    Odrv4 I__4142 (
            .O(N__19247),
            .I(\ppm_encoder_1.N_257_i_i ));
    Odrv4 I__4141 (
            .O(N__19244),
            .I(\ppm_encoder_1.N_257_i_i ));
    InMux I__4140 (
            .O(N__19239),
            .I(N__19236));
    LocalMux I__4139 (
            .O(N__19236),
            .I(N__19232));
    InMux I__4138 (
            .O(N__19235),
            .I(N__19227));
    Span4Mux_h I__4137 (
            .O(N__19232),
            .I(N__19224));
    InMux I__4136 (
            .O(N__19231),
            .I(N__19221));
    InMux I__4135 (
            .O(N__19230),
            .I(N__19218));
    LocalMux I__4134 (
            .O(N__19227),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__4133 (
            .O(N__19224),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    LocalMux I__4132 (
            .O(N__19221),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    LocalMux I__4131 (
            .O(N__19218),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__4130 (
            .O(N__19209),
            .I(N__19206));
    LocalMux I__4129 (
            .O(N__19206),
            .I(\ppm_encoder_1.pulses2count_9_0_0_6 ));
    InMux I__4128 (
            .O(N__19203),
            .I(N__19200));
    LocalMux I__4127 (
            .O(N__19200),
            .I(N__19197));
    Span4Mux_h I__4126 (
            .O(N__19197),
            .I(N__19194));
    Span4Mux_v I__4125 (
            .O(N__19194),
            .I(N__19191));
    Odrv4 I__4124 (
            .O(N__19191),
            .I(\ppm_encoder_1.N_301 ));
    CascadeMux I__4123 (
            .O(N__19188),
            .I(N__19184));
    InMux I__4122 (
            .O(N__19187),
            .I(N__19181));
    InMux I__4121 (
            .O(N__19184),
            .I(N__19177));
    LocalMux I__4120 (
            .O(N__19181),
            .I(N__19174));
    CascadeMux I__4119 (
            .O(N__19180),
            .I(N__19171));
    LocalMux I__4118 (
            .O(N__19177),
            .I(N__19167));
    Span4Mux_h I__4117 (
            .O(N__19174),
            .I(N__19164));
    InMux I__4116 (
            .O(N__19171),
            .I(N__19159));
    InMux I__4115 (
            .O(N__19170),
            .I(N__19159));
    Span4Mux_h I__4114 (
            .O(N__19167),
            .I(N__19156));
    Span4Mux_v I__4113 (
            .O(N__19164),
            .I(N__19153));
    LocalMux I__4112 (
            .O(N__19159),
            .I(N__19150));
    Odrv4 I__4111 (
            .O(N__19156),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv4 I__4110 (
            .O(N__19153),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv4 I__4109 (
            .O(N__19150),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    InMux I__4108 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__4107 (
            .O(N__19140),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__4106 (
            .O(N__19137),
            .I(N__19134));
    LocalMux I__4105 (
            .O(N__19134),
            .I(N__19131));
    Odrv12 I__4104 (
            .O(N__19131),
            .I(\ppm_encoder_1.N_302 ));
    CascadeMux I__4103 (
            .O(N__19128),
            .I(N__19125));
    InMux I__4102 (
            .O(N__19125),
            .I(N__19122));
    LocalMux I__4101 (
            .O(N__19122),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__4100 (
            .O(N__19119),
            .I(N__19116));
    LocalMux I__4099 (
            .O(N__19116),
            .I(\ppm_encoder_1.pulses2count_9_0_2_12 ));
    CascadeMux I__4098 (
            .O(N__19113),
            .I(N__19110));
    InMux I__4097 (
            .O(N__19110),
            .I(N__19107));
    LocalMux I__4096 (
            .O(N__19107),
            .I(N__19104));
    Odrv4 I__4095 (
            .O(N__19104),
            .I(\ppm_encoder_1.N_393 ));
    InMux I__4094 (
            .O(N__19101),
            .I(N__19098));
    LocalMux I__4093 (
            .O(N__19098),
            .I(N__19095));
    Odrv4 I__4092 (
            .O(N__19095),
            .I(\ppm_encoder_1.pulses2count_9_0_0_12 ));
    CascadeMux I__4091 (
            .O(N__19092),
            .I(N__19089));
    InMux I__4090 (
            .O(N__19089),
            .I(N__19085));
    CascadeMux I__4089 (
            .O(N__19088),
            .I(N__19082));
    LocalMux I__4088 (
            .O(N__19085),
            .I(N__19078));
    InMux I__4087 (
            .O(N__19082),
            .I(N__19075));
    InMux I__4086 (
            .O(N__19081),
            .I(N__19072));
    Span4Mux_v I__4085 (
            .O(N__19078),
            .I(N__19069));
    LocalMux I__4084 (
            .O(N__19075),
            .I(N__19066));
    LocalMux I__4083 (
            .O(N__19072),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    Odrv4 I__4082 (
            .O(N__19069),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    Odrv12 I__4081 (
            .O(N__19066),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    CascadeMux I__4080 (
            .O(N__19059),
            .I(N__19056));
    InMux I__4079 (
            .O(N__19056),
            .I(N__19053));
    LocalMux I__4078 (
            .O(N__19053),
            .I(N__19050));
    Odrv4 I__4077 (
            .O(N__19050),
            .I(\ppm_encoder_1.N_396 ));
    InMux I__4076 (
            .O(N__19047),
            .I(N__19044));
    LocalMux I__4075 (
            .O(N__19044),
            .I(N__19040));
    InMux I__4074 (
            .O(N__19043),
            .I(N__19037));
    Span4Mux_h I__4073 (
            .O(N__19040),
            .I(N__19033));
    LocalMux I__4072 (
            .O(N__19037),
            .I(N__19030));
    InMux I__4071 (
            .O(N__19036),
            .I(N__19027));
    Span4Mux_h I__4070 (
            .O(N__19033),
            .I(N__19024));
    Span4Mux_h I__4069 (
            .O(N__19030),
            .I(N__19021));
    LocalMux I__4068 (
            .O(N__19027),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    Odrv4 I__4067 (
            .O(N__19024),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    Odrv4 I__4066 (
            .O(N__19021),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__4065 (
            .O(N__19014),
            .I(N__19011));
    LocalMux I__4064 (
            .O(N__19011),
            .I(N__19007));
    CascadeMux I__4063 (
            .O(N__19010),
            .I(N__19004));
    Span4Mux_h I__4062 (
            .O(N__19007),
            .I(N__19001));
    InMux I__4061 (
            .O(N__19004),
            .I(N__18997));
    Span4Mux_v I__4060 (
            .O(N__19001),
            .I(N__18994));
    InMux I__4059 (
            .O(N__19000),
            .I(N__18991));
    LocalMux I__4058 (
            .O(N__18997),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__4057 (
            .O(N__18994),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    LocalMux I__4056 (
            .O(N__18991),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__4055 (
            .O(N__18984),
            .I(N__18981));
    LocalMux I__4054 (
            .O(N__18981),
            .I(N__18978));
    Span4Mux_h I__4053 (
            .O(N__18978),
            .I(N__18975));
    Odrv4 I__4052 (
            .O(N__18975),
            .I(\ppm_encoder_1.N_325 ));
    CascadeMux I__4051 (
            .O(N__18972),
            .I(\ppm_encoder_1.N_327_cascade_ ));
    InMux I__4050 (
            .O(N__18969),
            .I(N__18966));
    LocalMux I__4049 (
            .O(N__18966),
            .I(N__18962));
    CascadeMux I__4048 (
            .O(N__18965),
            .I(N__18959));
    Span4Mux_h I__4047 (
            .O(N__18962),
            .I(N__18956));
    InMux I__4046 (
            .O(N__18959),
            .I(N__18952));
    Span4Mux_h I__4045 (
            .O(N__18956),
            .I(N__18949));
    InMux I__4044 (
            .O(N__18955),
            .I(N__18946));
    LocalMux I__4043 (
            .O(N__18952),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__4042 (
            .O(N__18949),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    LocalMux I__4041 (
            .O(N__18946),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__4040 (
            .O(N__18939),
            .I(N__18936));
    LocalMux I__4039 (
            .O(N__18936),
            .I(N__18933));
    Span4Mux_h I__4038 (
            .O(N__18933),
            .I(N__18929));
    InMux I__4037 (
            .O(N__18932),
            .I(N__18926));
    Odrv4 I__4036 (
            .O(N__18929),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    LocalMux I__4035 (
            .O(N__18926),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    InMux I__4034 (
            .O(N__18921),
            .I(N__18917));
    InMux I__4033 (
            .O(N__18920),
            .I(N__18914));
    LocalMux I__4032 (
            .O(N__18917),
            .I(N__18911));
    LocalMux I__4031 (
            .O(N__18914),
            .I(N__18908));
    Odrv4 I__4030 (
            .O(N__18911),
            .I(\ppm_encoder_1.pulses2count_9_i_o2_0_5 ));
    Odrv4 I__4029 (
            .O(N__18908),
            .I(\ppm_encoder_1.pulses2count_9_i_o2_0_5 ));
    InMux I__4028 (
            .O(N__18903),
            .I(N__18894));
    InMux I__4027 (
            .O(N__18902),
            .I(N__18890));
    InMux I__4026 (
            .O(N__18901),
            .I(N__18887));
    CascadeMux I__4025 (
            .O(N__18900),
            .I(N__18882));
    InMux I__4024 (
            .O(N__18899),
            .I(N__18878));
    InMux I__4023 (
            .O(N__18898),
            .I(N__18871));
    InMux I__4022 (
            .O(N__18897),
            .I(N__18871));
    LocalMux I__4021 (
            .O(N__18894),
            .I(N__18868));
    InMux I__4020 (
            .O(N__18893),
            .I(N__18865));
    LocalMux I__4019 (
            .O(N__18890),
            .I(N__18860));
    LocalMux I__4018 (
            .O(N__18887),
            .I(N__18860));
    InMux I__4017 (
            .O(N__18886),
            .I(N__18855));
    InMux I__4016 (
            .O(N__18885),
            .I(N__18855));
    InMux I__4015 (
            .O(N__18882),
            .I(N__18851));
    CascadeMux I__4014 (
            .O(N__18881),
            .I(N__18848));
    LocalMux I__4013 (
            .O(N__18878),
            .I(N__18845));
    InMux I__4012 (
            .O(N__18877),
            .I(N__18842));
    InMux I__4011 (
            .O(N__18876),
            .I(N__18839));
    LocalMux I__4010 (
            .O(N__18871),
            .I(N__18836));
    Span4Mux_h I__4009 (
            .O(N__18868),
            .I(N__18827));
    LocalMux I__4008 (
            .O(N__18865),
            .I(N__18827));
    Span4Mux_v I__4007 (
            .O(N__18860),
            .I(N__18827));
    LocalMux I__4006 (
            .O(N__18855),
            .I(N__18827));
    InMux I__4005 (
            .O(N__18854),
            .I(N__18823));
    LocalMux I__4004 (
            .O(N__18851),
            .I(N__18820));
    InMux I__4003 (
            .O(N__18848),
            .I(N__18817));
    Span4Mux_h I__4002 (
            .O(N__18845),
            .I(N__18814));
    LocalMux I__4001 (
            .O(N__18842),
            .I(N__18805));
    LocalMux I__4000 (
            .O(N__18839),
            .I(N__18805));
    Span4Mux_v I__3999 (
            .O(N__18836),
            .I(N__18805));
    Span4Mux_h I__3998 (
            .O(N__18827),
            .I(N__18805));
    InMux I__3997 (
            .O(N__18826),
            .I(N__18802));
    LocalMux I__3996 (
            .O(N__18823),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv12 I__3995 (
            .O(N__18820),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__3994 (
            .O(N__18817),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__3993 (
            .O(N__18814),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__3992 (
            .O(N__18805),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__3991 (
            .O(N__18802),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    CascadeMux I__3990 (
            .O(N__18789),
            .I(N__18784));
    CascadeMux I__3989 (
            .O(N__18788),
            .I(N__18777));
    InMux I__3988 (
            .O(N__18787),
            .I(N__18772));
    InMux I__3987 (
            .O(N__18784),
            .I(N__18769));
    InMux I__3986 (
            .O(N__18783),
            .I(N__18764));
    InMux I__3985 (
            .O(N__18782),
            .I(N__18764));
    CascadeMux I__3984 (
            .O(N__18781),
            .I(N__18760));
    InMux I__3983 (
            .O(N__18780),
            .I(N__18756));
    InMux I__3982 (
            .O(N__18777),
            .I(N__18751));
    InMux I__3981 (
            .O(N__18776),
            .I(N__18751));
    InMux I__3980 (
            .O(N__18775),
            .I(N__18748));
    LocalMux I__3979 (
            .O(N__18772),
            .I(N__18745));
    LocalMux I__3978 (
            .O(N__18769),
            .I(N__18742));
    LocalMux I__3977 (
            .O(N__18764),
            .I(N__18736));
    InMux I__3976 (
            .O(N__18763),
            .I(N__18732));
    InMux I__3975 (
            .O(N__18760),
            .I(N__18727));
    InMux I__3974 (
            .O(N__18759),
            .I(N__18727));
    LocalMux I__3973 (
            .O(N__18756),
            .I(N__18724));
    LocalMux I__3972 (
            .O(N__18751),
            .I(N__18721));
    LocalMux I__3971 (
            .O(N__18748),
            .I(N__18716));
    Span4Mux_v I__3970 (
            .O(N__18745),
            .I(N__18716));
    Span4Mux_h I__3969 (
            .O(N__18742),
            .I(N__18713));
    InMux I__3968 (
            .O(N__18741),
            .I(N__18710));
    InMux I__3967 (
            .O(N__18740),
            .I(N__18707));
    InMux I__3966 (
            .O(N__18739),
            .I(N__18704));
    Span4Mux_h I__3965 (
            .O(N__18736),
            .I(N__18701));
    InMux I__3964 (
            .O(N__18735),
            .I(N__18698));
    LocalMux I__3963 (
            .O(N__18732),
            .I(N__18695));
    LocalMux I__3962 (
            .O(N__18727),
            .I(N__18692));
    Span4Mux_v I__3961 (
            .O(N__18724),
            .I(N__18687));
    Span4Mux_h I__3960 (
            .O(N__18721),
            .I(N__18687));
    Odrv4 I__3959 (
            .O(N__18716),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__3958 (
            .O(N__18713),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__3957 (
            .O(N__18710),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__3956 (
            .O(N__18707),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__3955 (
            .O(N__18704),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__3954 (
            .O(N__18701),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__3953 (
            .O(N__18698),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv12 I__3952 (
            .O(N__18695),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__3951 (
            .O(N__18692),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__3950 (
            .O(N__18687),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    InMux I__3949 (
            .O(N__18666),
            .I(N__18663));
    LocalMux I__3948 (
            .O(N__18663),
            .I(N__18660));
    Span4Mux_v I__3947 (
            .O(N__18660),
            .I(N__18657));
    Odrv4 I__3946 (
            .O(N__18657),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    CascadeMux I__3945 (
            .O(N__18654),
            .I(N__18650));
    CascadeMux I__3944 (
            .O(N__18653),
            .I(N__18647));
    InMux I__3943 (
            .O(N__18650),
            .I(N__18644));
    InMux I__3942 (
            .O(N__18647),
            .I(N__18641));
    LocalMux I__3941 (
            .O(N__18644),
            .I(N__18637));
    LocalMux I__3940 (
            .O(N__18641),
            .I(N__18634));
    InMux I__3939 (
            .O(N__18640),
            .I(N__18631));
    Span4Mux_v I__3938 (
            .O(N__18637),
            .I(N__18628));
    Span12Mux_h I__3937 (
            .O(N__18634),
            .I(N__18623));
    LocalMux I__3936 (
            .O(N__18631),
            .I(N__18623));
    Odrv4 I__3935 (
            .O(N__18628),
            .I(\ppm_encoder_1.N_204 ));
    Odrv12 I__3934 (
            .O(N__18623),
            .I(\ppm_encoder_1.N_204 ));
    CascadeMux I__3933 (
            .O(N__18618),
            .I(N__18615));
    InMux I__3932 (
            .O(N__18615),
            .I(N__18612));
    LocalMux I__3931 (
            .O(N__18612),
            .I(N__18608));
    InMux I__3930 (
            .O(N__18611),
            .I(N__18605));
    Span4Mux_v I__3929 (
            .O(N__18608),
            .I(N__18600));
    LocalMux I__3928 (
            .O(N__18605),
            .I(N__18600));
    Odrv4 I__3927 (
            .O(N__18600),
            .I(\ppm_encoder_1.N_255_i_i ));
    CascadeMux I__3926 (
            .O(N__18597),
            .I(\ppm_encoder_1.N_204_cascade_ ));
    InMux I__3925 (
            .O(N__18594),
            .I(N__18591));
    LocalMux I__3924 (
            .O(N__18591),
            .I(N__18586));
    InMux I__3923 (
            .O(N__18590),
            .I(N__18581));
    InMux I__3922 (
            .O(N__18589),
            .I(N__18581));
    Odrv4 I__3921 (
            .O(N__18586),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    LocalMux I__3920 (
            .O(N__18581),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__3919 (
            .O(N__18576),
            .I(N__18573));
    LocalMux I__3918 (
            .O(N__18573),
            .I(N__18568));
    InMux I__3917 (
            .O(N__18572),
            .I(N__18563));
    InMux I__3916 (
            .O(N__18571),
            .I(N__18563));
    Odrv4 I__3915 (
            .O(N__18568),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__3914 (
            .O(N__18563),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__3913 (
            .O(N__18558),
            .I(\ppm_encoder_1.N_379_cascade_ ));
    CascadeMux I__3912 (
            .O(N__18555),
            .I(N__18552));
    InMux I__3911 (
            .O(N__18552),
            .I(N__18547));
    InMux I__3910 (
            .O(N__18551),
            .I(N__18544));
    InMux I__3909 (
            .O(N__18550),
            .I(N__18541));
    LocalMux I__3908 (
            .O(N__18547),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    LocalMux I__3907 (
            .O(N__18544),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    LocalMux I__3906 (
            .O(N__18541),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    InMux I__3905 (
            .O(N__18534),
            .I(N__18529));
    InMux I__3904 (
            .O(N__18533),
            .I(N__18526));
    InMux I__3903 (
            .O(N__18532),
            .I(N__18523));
    LocalMux I__3902 (
            .O(N__18529),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    LocalMux I__3901 (
            .O(N__18526),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    LocalMux I__3900 (
            .O(N__18523),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__3899 (
            .O(N__18516),
            .I(N__18513));
    LocalMux I__3898 (
            .O(N__18513),
            .I(N__18509));
    InMux I__3897 (
            .O(N__18512),
            .I(N__18506));
    Odrv4 I__3896 (
            .O(N__18509),
            .I(\ppm_encoder_1.pulses2count_9_i_o2_0_7 ));
    LocalMux I__3895 (
            .O(N__18506),
            .I(\ppm_encoder_1.pulses2count_9_i_o2_0_7 ));
    InMux I__3894 (
            .O(N__18501),
            .I(N__18498));
    LocalMux I__3893 (
            .O(N__18498),
            .I(N__18495));
    Span4Mux_h I__3892 (
            .O(N__18495),
            .I(N__18490));
    InMux I__3891 (
            .O(N__18494),
            .I(N__18487));
    CascadeMux I__3890 (
            .O(N__18493),
            .I(N__18484));
    Span4Mux_v I__3889 (
            .O(N__18490),
            .I(N__18479));
    LocalMux I__3888 (
            .O(N__18487),
            .I(N__18479));
    InMux I__3887 (
            .O(N__18484),
            .I(N__18476));
    Span4Mux_h I__3886 (
            .O(N__18479),
            .I(N__18473));
    LocalMux I__3885 (
            .O(N__18476),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__3884 (
            .O(N__18473),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    InMux I__3883 (
            .O(N__18468),
            .I(N__18465));
    LocalMux I__3882 (
            .O(N__18465),
            .I(N__18462));
    Span4Mux_h I__3881 (
            .O(N__18462),
            .I(N__18459));
    Span4Mux_v I__3880 (
            .O(N__18459),
            .I(N__18454));
    InMux I__3879 (
            .O(N__18458),
            .I(N__18449));
    InMux I__3878 (
            .O(N__18457),
            .I(N__18449));
    Odrv4 I__3877 (
            .O(N__18454),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    LocalMux I__3876 (
            .O(N__18449),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    CascadeMux I__3875 (
            .O(N__18444),
            .I(N__18441));
    InMux I__3874 (
            .O(N__18441),
            .I(N__18438));
    LocalMux I__3873 (
            .O(N__18438),
            .I(\ppm_encoder_1.pulses2count_9_i_0_8 ));
    InMux I__3872 (
            .O(N__18435),
            .I(N__18432));
    LocalMux I__3871 (
            .O(N__18432),
            .I(N__18429));
    Span4Mux_h I__3870 (
            .O(N__18429),
            .I(N__18424));
    InMux I__3869 (
            .O(N__18428),
            .I(N__18419));
    InMux I__3868 (
            .O(N__18427),
            .I(N__18419));
    Odrv4 I__3867 (
            .O(N__18424),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    LocalMux I__3866 (
            .O(N__18419),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__3865 (
            .O(N__18414),
            .I(N__18410));
    CascadeMux I__3864 (
            .O(N__18413),
            .I(N__18407));
    LocalMux I__3863 (
            .O(N__18410),
            .I(N__18403));
    InMux I__3862 (
            .O(N__18407),
            .I(N__18400));
    InMux I__3861 (
            .O(N__18406),
            .I(N__18397));
    Span4Mux_h I__3860 (
            .O(N__18403),
            .I(N__18392));
    LocalMux I__3859 (
            .O(N__18400),
            .I(N__18392));
    LocalMux I__3858 (
            .O(N__18397),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__3857 (
            .O(N__18392),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    CascadeMux I__3856 (
            .O(N__18387),
            .I(N__18384));
    InMux I__3855 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__3854 (
            .O(N__18381),
            .I(\ppm_encoder_1.N_391 ));
    InMux I__3853 (
            .O(N__18378),
            .I(N__18375));
    LocalMux I__3852 (
            .O(N__18375),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__3851 (
            .O(N__18372),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__3850 (
            .O(N__18369),
            .I(N__18366));
    LocalMux I__3849 (
            .O(N__18366),
            .I(N__18363));
    Span4Mux_v I__3848 (
            .O(N__18363),
            .I(N__18360));
    Odrv4 I__3847 (
            .O(N__18360),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__3846 (
            .O(N__18357),
            .I(bfn_9_28_0_));
    CascadeMux I__3845 (
            .O(N__18354),
            .I(N__18351));
    InMux I__3844 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__3843 (
            .O(N__18348),
            .I(N__18345));
    Odrv4 I__3842 (
            .O(N__18345),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__3841 (
            .O(N__18342),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__3840 (
            .O(N__18339),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__3839 (
            .O(N__18336),
            .I(N__18333));
    LocalMux I__3838 (
            .O(N__18333),
            .I(N__18330));
    Odrv4 I__3837 (
            .O(N__18330),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__3836 (
            .O(N__18327),
            .I(N__18324));
    LocalMux I__3835 (
            .O(N__18324),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__3834 (
            .O(N__18321),
            .I(N__18318));
    LocalMux I__3833 (
            .O(N__18318),
            .I(N__18314));
    CascadeMux I__3832 (
            .O(N__18317),
            .I(N__18311));
    Span4Mux_h I__3831 (
            .O(N__18314),
            .I(N__18308));
    InMux I__3830 (
            .O(N__18311),
            .I(N__18305));
    Odrv4 I__3829 (
            .O(N__18308),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    LocalMux I__3828 (
            .O(N__18305),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__3827 (
            .O(N__18300),
            .I(N__18297));
    LocalMux I__3826 (
            .O(N__18297),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    CascadeMux I__3825 (
            .O(N__18294),
            .I(N__18291));
    InMux I__3824 (
            .O(N__18291),
            .I(N__18286));
    CascadeMux I__3823 (
            .O(N__18290),
            .I(N__18283));
    InMux I__3822 (
            .O(N__18289),
            .I(N__18280));
    LocalMux I__3821 (
            .O(N__18286),
            .I(N__18277));
    InMux I__3820 (
            .O(N__18283),
            .I(N__18274));
    LocalMux I__3819 (
            .O(N__18280),
            .I(N__18270));
    Span4Mux_v I__3818 (
            .O(N__18277),
            .I(N__18267));
    LocalMux I__3817 (
            .O(N__18274),
            .I(N__18264));
    CascadeMux I__3816 (
            .O(N__18273),
            .I(N__18261));
    Span4Mux_h I__3815 (
            .O(N__18270),
            .I(N__18258));
    Span4Mux_h I__3814 (
            .O(N__18267),
            .I(N__18253));
    Span4Mux_v I__3813 (
            .O(N__18264),
            .I(N__18253));
    InMux I__3812 (
            .O(N__18261),
            .I(N__18250));
    Odrv4 I__3811 (
            .O(N__18258),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    Odrv4 I__3810 (
            .O(N__18253),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    LocalMux I__3809 (
            .O(N__18250),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    InMux I__3808 (
            .O(N__18243),
            .I(N__18240));
    LocalMux I__3807 (
            .O(N__18240),
            .I(N__18237));
    Odrv4 I__3806 (
            .O(N__18237),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__3805 (
            .O(N__18234),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    CascadeMux I__3804 (
            .O(N__18231),
            .I(N__18228));
    InMux I__3803 (
            .O(N__18228),
            .I(N__18225));
    LocalMux I__3802 (
            .O(N__18225),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__3801 (
            .O(N__18222),
            .I(bfn_9_27_0_));
    InMux I__3800 (
            .O(N__18219),
            .I(N__18216));
    LocalMux I__3799 (
            .O(N__18216),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__3798 (
            .O(N__18213),
            .I(N__18210));
    LocalMux I__3797 (
            .O(N__18210),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__3796 (
            .O(N__18207),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__3795 (
            .O(N__18204),
            .I(N__18201));
    LocalMux I__3794 (
            .O(N__18201),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__3793 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__3792 (
            .O(N__18195),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__3791 (
            .O(N__18192),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    CascadeMux I__3790 (
            .O(N__18189),
            .I(N__18186));
    InMux I__3789 (
            .O(N__18186),
            .I(N__18183));
    LocalMux I__3788 (
            .O(N__18183),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__3787 (
            .O(N__18180),
            .I(N__18177));
    LocalMux I__3786 (
            .O(N__18177),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__3785 (
            .O(N__18174),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__3784 (
            .O(N__18171),
            .I(N__18168));
    LocalMux I__3783 (
            .O(N__18168),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__3782 (
            .O(N__18165),
            .I(N__18162));
    LocalMux I__3781 (
            .O(N__18162),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__3780 (
            .O(N__18159),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__3779 (
            .O(N__18156),
            .I(N__18153));
    LocalMux I__3778 (
            .O(N__18153),
            .I(N__18149));
    InMux I__3777 (
            .O(N__18152),
            .I(N__18146));
    Span4Mux_v I__3776 (
            .O(N__18149),
            .I(N__18140));
    LocalMux I__3775 (
            .O(N__18146),
            .I(N__18140));
    InMux I__3774 (
            .O(N__18145),
            .I(N__18137));
    Span4Mux_h I__3773 (
            .O(N__18140),
            .I(N__18132));
    LocalMux I__3772 (
            .O(N__18137),
            .I(N__18132));
    Span4Mux_s3_v I__3771 (
            .O(N__18132),
            .I(N__18128));
    InMux I__3770 (
            .O(N__18131),
            .I(N__18125));
    Odrv4 I__3769 (
            .O(N__18128),
            .I(\ppm_encoder_1.N_259_i_i ));
    LocalMux I__3768 (
            .O(N__18125),
            .I(\ppm_encoder_1.N_259_i_i ));
    CascadeMux I__3767 (
            .O(N__18120),
            .I(N__18117));
    InMux I__3766 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__3765 (
            .O(N__18114),
            .I(\ppm_encoder_1.init_pulses_RNIKON03Z0Z_13 ));
    InMux I__3764 (
            .O(N__18111),
            .I(N__18108));
    LocalMux I__3763 (
            .O(N__18108),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__3762 (
            .O(N__18105),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__3761 (
            .O(N__18102),
            .I(N__18099));
    LocalMux I__3760 (
            .O(N__18099),
            .I(N__18096));
    Odrv4 I__3759 (
            .O(N__18096),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO ));
    InMux I__3758 (
            .O(N__18093),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    CascadeMux I__3757 (
            .O(N__18090),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_ ));
    InMux I__3756 (
            .O(N__18087),
            .I(N__18084));
    LocalMux I__3755 (
            .O(N__18084),
            .I(N__18081));
    Span4Mux_v I__3754 (
            .O(N__18081),
            .I(N__18078));
    Odrv4 I__3753 (
            .O(N__18078),
            .I(\ppm_encoder_1.init_pulses_RNI83R42Z0Z_0 ));
    InMux I__3752 (
            .O(N__18075),
            .I(N__18072));
    LocalMux I__3751 (
            .O(N__18072),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__3750 (
            .O(N__18069),
            .I(N__18066));
    LocalMux I__3749 (
            .O(N__18066),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__3748 (
            .O(N__18063),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__3747 (
            .O(N__18060),
            .I(N__18057));
    LocalMux I__3746 (
            .O(N__18057),
            .I(\ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2 ));
    CascadeMux I__3745 (
            .O(N__18054),
            .I(N__18051));
    InMux I__3744 (
            .O(N__18051),
            .I(N__18048));
    LocalMux I__3743 (
            .O(N__18048),
            .I(N__18044));
    CascadeMux I__3742 (
            .O(N__18047),
            .I(N__18041));
    Span4Mux_h I__3741 (
            .O(N__18044),
            .I(N__18036));
    InMux I__3740 (
            .O(N__18041),
            .I(N__18033));
    InMux I__3739 (
            .O(N__18040),
            .I(N__18030));
    InMux I__3738 (
            .O(N__18039),
            .I(N__18027));
    Odrv4 I__3737 (
            .O(N__18036),
            .I(\ppm_encoder_1.N_249_i_i ));
    LocalMux I__3736 (
            .O(N__18033),
            .I(\ppm_encoder_1.N_249_i_i ));
    LocalMux I__3735 (
            .O(N__18030),
            .I(\ppm_encoder_1.N_249_i_i ));
    LocalMux I__3734 (
            .O(N__18027),
            .I(\ppm_encoder_1.N_249_i_i ));
    InMux I__3733 (
            .O(N__18018),
            .I(N__18015));
    LocalMux I__3732 (
            .O(N__18015),
            .I(N__18012));
    Span4Mux_v I__3731 (
            .O(N__18012),
            .I(N__18009));
    Odrv4 I__3730 (
            .O(N__18009),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__3729 (
            .O(N__18006),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__3728 (
            .O(N__18003),
            .I(N__18000));
    LocalMux I__3727 (
            .O(N__18000),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__3726 (
            .O(N__17997),
            .I(N__17994));
    LocalMux I__3725 (
            .O(N__17994),
            .I(N__17991));
    Odrv4 I__3724 (
            .O(N__17991),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__3723 (
            .O(N__17988),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__3722 (
            .O(N__17985),
            .I(N__17982));
    LocalMux I__3721 (
            .O(N__17982),
            .I(N__17979));
    Span4Mux_v I__3720 (
            .O(N__17979),
            .I(N__17976));
    Odrv4 I__3719 (
            .O(N__17976),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__3718 (
            .O(N__17973),
            .I(N__17970));
    LocalMux I__3717 (
            .O(N__17970),
            .I(N__17967));
    Span4Mux_h I__3716 (
            .O(N__17967),
            .I(N__17964));
    Odrv4 I__3715 (
            .O(N__17964),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__3714 (
            .O(N__17961),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__3713 (
            .O(N__17958),
            .I(N__17955));
    LocalMux I__3712 (
            .O(N__17955),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__3711 (
            .O(N__17952),
            .I(N__17949));
    LocalMux I__3710 (
            .O(N__17949),
            .I(N__17946));
    Odrv4 I__3709 (
            .O(N__17946),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__3708 (
            .O(N__17943),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__3707 (
            .O(N__17940),
            .I(N__17937));
    LocalMux I__3706 (
            .O(N__17937),
            .I(\ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6 ));
    CascadeMux I__3705 (
            .O(N__17934),
            .I(N__17930));
    InMux I__3704 (
            .O(N__17933),
            .I(N__17926));
    InMux I__3703 (
            .O(N__17930),
            .I(N__17923));
    CascadeMux I__3702 (
            .O(N__17929),
            .I(N__17920));
    LocalMux I__3701 (
            .O(N__17926),
            .I(N__17917));
    LocalMux I__3700 (
            .O(N__17923),
            .I(N__17913));
    InMux I__3699 (
            .O(N__17920),
            .I(N__17910));
    Span4Mux_v I__3698 (
            .O(N__17917),
            .I(N__17907));
    InMux I__3697 (
            .O(N__17916),
            .I(N__17904));
    Odrv4 I__3696 (
            .O(N__17913),
            .I(\ppm_encoder_1.N_253_i_i ));
    LocalMux I__3695 (
            .O(N__17910),
            .I(\ppm_encoder_1.N_253_i_i ));
    Odrv4 I__3694 (
            .O(N__17907),
            .I(\ppm_encoder_1.N_253_i_i ));
    LocalMux I__3693 (
            .O(N__17904),
            .I(\ppm_encoder_1.N_253_i_i ));
    InMux I__3692 (
            .O(N__17895),
            .I(N__17892));
    LocalMux I__3691 (
            .O(N__17892),
            .I(N__17889));
    Odrv4 I__3690 (
            .O(N__17889),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__3689 (
            .O(N__17886),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__3688 (
            .O(N__17883),
            .I(N__17880));
    LocalMux I__3687 (
            .O(N__17880),
            .I(N__17876));
    InMux I__3686 (
            .O(N__17879),
            .I(N__17873));
    Span4Mux_v I__3685 (
            .O(N__17876),
            .I(N__17866));
    LocalMux I__3684 (
            .O(N__17873),
            .I(N__17866));
    InMux I__3683 (
            .O(N__17872),
            .I(N__17861));
    InMux I__3682 (
            .O(N__17871),
            .I(N__17858));
    Span4Mux_h I__3681 (
            .O(N__17866),
            .I(N__17855));
    InMux I__3680 (
            .O(N__17865),
            .I(N__17850));
    InMux I__3679 (
            .O(N__17864),
            .I(N__17850));
    LocalMux I__3678 (
            .O(N__17861),
            .I(N__17847));
    LocalMux I__3677 (
            .O(N__17858),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    Odrv4 I__3676 (
            .O(N__17855),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__3675 (
            .O(N__17850),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    Odrv4 I__3674 (
            .O(N__17847),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__3673 (
            .O(N__17838),
            .I(N__17835));
    InMux I__3672 (
            .O(N__17835),
            .I(N__17831));
    InMux I__3671 (
            .O(N__17834),
            .I(N__17828));
    LocalMux I__3670 (
            .O(N__17831),
            .I(N__17825));
    LocalMux I__3669 (
            .O(N__17828),
            .I(N__17822));
    Odrv4 I__3668 (
            .O(N__17825),
            .I(\ppm_encoder_1.N_256_i_i ));
    Odrv12 I__3667 (
            .O(N__17822),
            .I(\ppm_encoder_1.N_256_i_i ));
    CascadeMux I__3666 (
            .O(N__17817),
            .I(N__17814));
    InMux I__3665 (
            .O(N__17814),
            .I(N__17808));
    CascadeMux I__3664 (
            .O(N__17813),
            .I(N__17799));
    InMux I__3663 (
            .O(N__17812),
            .I(N__17796));
    InMux I__3662 (
            .O(N__17811),
            .I(N__17793));
    LocalMux I__3661 (
            .O(N__17808),
            .I(N__17790));
    InMux I__3660 (
            .O(N__17807),
            .I(N__17787));
    InMux I__3659 (
            .O(N__17806),
            .I(N__17782));
    InMux I__3658 (
            .O(N__17805),
            .I(N__17782));
    InMux I__3657 (
            .O(N__17804),
            .I(N__17777));
    InMux I__3656 (
            .O(N__17803),
            .I(N__17777));
    InMux I__3655 (
            .O(N__17802),
            .I(N__17772));
    InMux I__3654 (
            .O(N__17799),
            .I(N__17772));
    LocalMux I__3653 (
            .O(N__17796),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__3652 (
            .O(N__17793),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    Odrv4 I__3651 (
            .O(N__17790),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__3650 (
            .O(N__17787),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__3649 (
            .O(N__17782),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__3648 (
            .O(N__17777),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__3647 (
            .O(N__17772),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    InMux I__3646 (
            .O(N__17757),
            .I(N__17754));
    LocalMux I__3645 (
            .O(N__17754),
            .I(N__17751));
    Odrv4 I__3644 (
            .O(N__17751),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__3643 (
            .O(N__17748),
            .I(N__17745));
    LocalMux I__3642 (
            .O(N__17745),
            .I(N__17741));
    InMux I__3641 (
            .O(N__17744),
            .I(N__17738));
    Span4Mux_h I__3640 (
            .O(N__17741),
            .I(N__17730));
    LocalMux I__3639 (
            .O(N__17738),
            .I(N__17730));
    InMux I__3638 (
            .O(N__17737),
            .I(N__17723));
    InMux I__3637 (
            .O(N__17736),
            .I(N__17723));
    InMux I__3636 (
            .O(N__17735),
            .I(N__17723));
    Odrv4 I__3635 (
            .O(N__17730),
            .I(\ppm_encoder_1.N_305 ));
    LocalMux I__3634 (
            .O(N__17723),
            .I(\ppm_encoder_1.N_305 ));
    InMux I__3633 (
            .O(N__17718),
            .I(N__17706));
    InMux I__3632 (
            .O(N__17717),
            .I(N__17700));
    InMux I__3631 (
            .O(N__17716),
            .I(N__17697));
    InMux I__3630 (
            .O(N__17715),
            .I(N__17694));
    InMux I__3629 (
            .O(N__17714),
            .I(N__17691));
    InMux I__3628 (
            .O(N__17713),
            .I(N__17688));
    InMux I__3627 (
            .O(N__17712),
            .I(N__17684));
    InMux I__3626 (
            .O(N__17711),
            .I(N__17681));
    InMux I__3625 (
            .O(N__17710),
            .I(N__17676));
    InMux I__3624 (
            .O(N__17709),
            .I(N__17676));
    LocalMux I__3623 (
            .O(N__17706),
            .I(N__17673));
    InMux I__3622 (
            .O(N__17705),
            .I(N__17670));
    CascadeMux I__3621 (
            .O(N__17704),
            .I(N__17663));
    InMux I__3620 (
            .O(N__17703),
            .I(N__17660));
    LocalMux I__3619 (
            .O(N__17700),
            .I(N__17657));
    LocalMux I__3618 (
            .O(N__17697),
            .I(N__17650));
    LocalMux I__3617 (
            .O(N__17694),
            .I(N__17650));
    LocalMux I__3616 (
            .O(N__17691),
            .I(N__17650));
    LocalMux I__3615 (
            .O(N__17688),
            .I(N__17647));
    InMux I__3614 (
            .O(N__17687),
            .I(N__17644));
    LocalMux I__3613 (
            .O(N__17684),
            .I(N__17637));
    LocalMux I__3612 (
            .O(N__17681),
            .I(N__17637));
    LocalMux I__3611 (
            .O(N__17676),
            .I(N__17637));
    Span4Mux_v I__3610 (
            .O(N__17673),
            .I(N__17632));
    LocalMux I__3609 (
            .O(N__17670),
            .I(N__17632));
    InMux I__3608 (
            .O(N__17669),
            .I(N__17629));
    InMux I__3607 (
            .O(N__17668),
            .I(N__17626));
    InMux I__3606 (
            .O(N__17667),
            .I(N__17623));
    InMux I__3605 (
            .O(N__17666),
            .I(N__17618));
    InMux I__3604 (
            .O(N__17663),
            .I(N__17618));
    LocalMux I__3603 (
            .O(N__17660),
            .I(N__17613));
    Span4Mux_h I__3602 (
            .O(N__17657),
            .I(N__17613));
    Span4Mux_v I__3601 (
            .O(N__17650),
            .I(N__17604));
    Span4Mux_h I__3600 (
            .O(N__17647),
            .I(N__17604));
    LocalMux I__3599 (
            .O(N__17644),
            .I(N__17604));
    Span4Mux_v I__3598 (
            .O(N__17637),
            .I(N__17604));
    Span4Mux_h I__3597 (
            .O(N__17632),
            .I(N__17601));
    LocalMux I__3596 (
            .O(N__17629),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    LocalMux I__3595 (
            .O(N__17626),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    LocalMux I__3594 (
            .O(N__17623),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    LocalMux I__3593 (
            .O(N__17618),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    Odrv4 I__3592 (
            .O(N__17613),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    Odrv4 I__3591 (
            .O(N__17604),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    Odrv4 I__3590 (
            .O(N__17601),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ));
    CascadeMux I__3589 (
            .O(N__17586),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_ ));
    InMux I__3588 (
            .O(N__17583),
            .I(N__17580));
    LocalMux I__3587 (
            .O(N__17580),
            .I(N__17576));
    InMux I__3586 (
            .O(N__17579),
            .I(N__17573));
    Span4Mux_v I__3585 (
            .O(N__17576),
            .I(N__17568));
    LocalMux I__3584 (
            .O(N__17573),
            .I(N__17568));
    Odrv4 I__3583 (
            .O(N__17568),
            .I(\ppm_encoder_1.N_260_i_i ));
    CascadeMux I__3582 (
            .O(N__17565),
            .I(N__17556));
    CascadeMux I__3581 (
            .O(N__17564),
            .I(N__17553));
    InMux I__3580 (
            .O(N__17563),
            .I(N__17549));
    CascadeMux I__3579 (
            .O(N__17562),
            .I(N__17545));
    CascadeMux I__3578 (
            .O(N__17561),
            .I(N__17542));
    CascadeMux I__3577 (
            .O(N__17560),
            .I(N__17536));
    CascadeMux I__3576 (
            .O(N__17559),
            .I(N__17531));
    InMux I__3575 (
            .O(N__17556),
            .I(N__17524));
    InMux I__3574 (
            .O(N__17553),
            .I(N__17524));
    CascadeMux I__3573 (
            .O(N__17552),
            .I(N__17521));
    LocalMux I__3572 (
            .O(N__17549),
            .I(N__17517));
    InMux I__3571 (
            .O(N__17548),
            .I(N__17510));
    InMux I__3570 (
            .O(N__17545),
            .I(N__17510));
    InMux I__3569 (
            .O(N__17542),
            .I(N__17510));
    CascadeMux I__3568 (
            .O(N__17541),
            .I(N__17504));
    CascadeMux I__3567 (
            .O(N__17540),
            .I(N__17501));
    InMux I__3566 (
            .O(N__17539),
            .I(N__17496));
    InMux I__3565 (
            .O(N__17536),
            .I(N__17496));
    CascadeMux I__3564 (
            .O(N__17535),
            .I(N__17493));
    InMux I__3563 (
            .O(N__17534),
            .I(N__17488));
    InMux I__3562 (
            .O(N__17531),
            .I(N__17488));
    CascadeMux I__3561 (
            .O(N__17530),
            .I(N__17480));
    CascadeMux I__3560 (
            .O(N__17529),
            .I(N__17477));
    LocalMux I__3559 (
            .O(N__17524),
            .I(N__17473));
    InMux I__3558 (
            .O(N__17521),
            .I(N__17468));
    InMux I__3557 (
            .O(N__17520),
            .I(N__17468));
    Span4Mux_h I__3556 (
            .O(N__17517),
            .I(N__17463));
    LocalMux I__3555 (
            .O(N__17510),
            .I(N__17463));
    CascadeMux I__3554 (
            .O(N__17509),
            .I(N__17455));
    InMux I__3553 (
            .O(N__17508),
            .I(N__17448));
    InMux I__3552 (
            .O(N__17507),
            .I(N__17448));
    InMux I__3551 (
            .O(N__17504),
            .I(N__17448));
    InMux I__3550 (
            .O(N__17501),
            .I(N__17445));
    LocalMux I__3549 (
            .O(N__17496),
            .I(N__17442));
    InMux I__3548 (
            .O(N__17493),
            .I(N__17439));
    LocalMux I__3547 (
            .O(N__17488),
            .I(N__17436));
    InMux I__3546 (
            .O(N__17487),
            .I(N__17429));
    InMux I__3545 (
            .O(N__17486),
            .I(N__17414));
    InMux I__3544 (
            .O(N__17485),
            .I(N__17414));
    InMux I__3543 (
            .O(N__17484),
            .I(N__17414));
    InMux I__3542 (
            .O(N__17483),
            .I(N__17414));
    InMux I__3541 (
            .O(N__17480),
            .I(N__17414));
    InMux I__3540 (
            .O(N__17477),
            .I(N__17414));
    InMux I__3539 (
            .O(N__17476),
            .I(N__17414));
    Span4Mux_s3_v I__3538 (
            .O(N__17473),
            .I(N__17411));
    LocalMux I__3537 (
            .O(N__17468),
            .I(N__17406));
    Span4Mux_v I__3536 (
            .O(N__17463),
            .I(N__17406));
    InMux I__3535 (
            .O(N__17462),
            .I(N__17403));
    CascadeMux I__3534 (
            .O(N__17461),
            .I(N__17400));
    CascadeMux I__3533 (
            .O(N__17460),
            .I(N__17397));
    InMux I__3532 (
            .O(N__17459),
            .I(N__17390));
    InMux I__3531 (
            .O(N__17458),
            .I(N__17390));
    InMux I__3530 (
            .O(N__17455),
            .I(N__17390));
    LocalMux I__3529 (
            .O(N__17448),
            .I(N__17383));
    LocalMux I__3528 (
            .O(N__17445),
            .I(N__17383));
    Span4Mux_s3_v I__3527 (
            .O(N__17442),
            .I(N__17383));
    LocalMux I__3526 (
            .O(N__17439),
            .I(N__17380));
    Span4Mux_h I__3525 (
            .O(N__17436),
            .I(N__17377));
    InMux I__3524 (
            .O(N__17435),
            .I(N__17374));
    InMux I__3523 (
            .O(N__17434),
            .I(N__17367));
    InMux I__3522 (
            .O(N__17433),
            .I(N__17367));
    InMux I__3521 (
            .O(N__17432),
            .I(N__17367));
    LocalMux I__3520 (
            .O(N__17429),
            .I(N__17364));
    LocalMux I__3519 (
            .O(N__17414),
            .I(N__17359));
    Span4Mux_h I__3518 (
            .O(N__17411),
            .I(N__17359));
    Span4Mux_h I__3517 (
            .O(N__17406),
            .I(N__17354));
    LocalMux I__3516 (
            .O(N__17403),
            .I(N__17354));
    InMux I__3515 (
            .O(N__17400),
            .I(N__17351));
    InMux I__3514 (
            .O(N__17397),
            .I(N__17348));
    LocalMux I__3513 (
            .O(N__17390),
            .I(N__17345));
    Span4Mux_v I__3512 (
            .O(N__17383),
            .I(N__17342));
    Span12Mux_h I__3511 (
            .O(N__17380),
            .I(N__17339));
    Sp12to4 I__3510 (
            .O(N__17377),
            .I(N__17336));
    LocalMux I__3509 (
            .O(N__17374),
            .I(N__17325));
    LocalMux I__3508 (
            .O(N__17367),
            .I(N__17325));
    Span4Mux_h I__3507 (
            .O(N__17364),
            .I(N__17325));
    Span4Mux_v I__3506 (
            .O(N__17359),
            .I(N__17325));
    Span4Mux_h I__3505 (
            .O(N__17354),
            .I(N__17325));
    LocalMux I__3504 (
            .O(N__17351),
            .I(scaler_1_dv));
    LocalMux I__3503 (
            .O(N__17348),
            .I(scaler_1_dv));
    Odrv12 I__3502 (
            .O(N__17345),
            .I(scaler_1_dv));
    Odrv4 I__3501 (
            .O(N__17342),
            .I(scaler_1_dv));
    Odrv12 I__3500 (
            .O(N__17339),
            .I(scaler_1_dv));
    Odrv12 I__3499 (
            .O(N__17336),
            .I(scaler_1_dv));
    Odrv4 I__3498 (
            .O(N__17325),
            .I(scaler_1_dv));
    InMux I__3497 (
            .O(N__17310),
            .I(N__17307));
    LocalMux I__3496 (
            .O(N__17307),
            .I(N__17301));
    InMux I__3495 (
            .O(N__17306),
            .I(N__17296));
    InMux I__3494 (
            .O(N__17305),
            .I(N__17296));
    InMux I__3493 (
            .O(N__17304),
            .I(N__17293));
    Span4Mux_h I__3492 (
            .O(N__17301),
            .I(N__17288));
    LocalMux I__3491 (
            .O(N__17296),
            .I(N__17288));
    LocalMux I__3490 (
            .O(N__17293),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv4 I__3489 (
            .O(N__17288),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    CascadeMux I__3488 (
            .O(N__17283),
            .I(N__17280));
    InMux I__3487 (
            .O(N__17280),
            .I(N__17277));
    LocalMux I__3486 (
            .O(N__17277),
            .I(N__17273));
    InMux I__3485 (
            .O(N__17276),
            .I(N__17270));
    Odrv4 I__3484 (
            .O(N__17273),
            .I(\ppm_encoder_1.N_248_i_i ));
    LocalMux I__3483 (
            .O(N__17270),
            .I(\ppm_encoder_1.N_248_i_i ));
    CascadeMux I__3482 (
            .O(N__17265),
            .I(N__17262));
    InMux I__3481 (
            .O(N__17262),
            .I(N__17259));
    LocalMux I__3480 (
            .O(N__17259),
            .I(N__17255));
    InMux I__3479 (
            .O(N__17258),
            .I(N__17252));
    Odrv4 I__3478 (
            .O(N__17255),
            .I(\ppm_encoder_1.N_250_i_i ));
    LocalMux I__3477 (
            .O(N__17252),
            .I(\ppm_encoder_1.N_250_i_i ));
    CascadeMux I__3476 (
            .O(N__17247),
            .I(N__17244));
    InMux I__3475 (
            .O(N__17244),
            .I(N__17241));
    LocalMux I__3474 (
            .O(N__17241),
            .I(N__17238));
    Span4Mux_v I__3473 (
            .O(N__17238),
            .I(N__17235));
    Span4Mux_h I__3472 (
            .O(N__17235),
            .I(N__17231));
    InMux I__3471 (
            .O(N__17234),
            .I(N__17228));
    Odrv4 I__3470 (
            .O(N__17231),
            .I(\ppm_encoder_1.N_254_i_i ));
    LocalMux I__3469 (
            .O(N__17228),
            .I(\ppm_encoder_1.N_254_i_i ));
    CascadeMux I__3468 (
            .O(N__17223),
            .I(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ));
    CascadeMux I__3467 (
            .O(N__17220),
            .I(N__17217));
    InMux I__3466 (
            .O(N__17217),
            .I(N__17213));
    InMux I__3465 (
            .O(N__17216),
            .I(N__17210));
    LocalMux I__3464 (
            .O(N__17213),
            .I(N__17205));
    LocalMux I__3463 (
            .O(N__17210),
            .I(N__17205));
    Odrv12 I__3462 (
            .O(N__17205),
            .I(\ppm_encoder_1.N_246_i_i ));
    CascadeMux I__3461 (
            .O(N__17202),
            .I(\ppm_encoder_1.un2_throttle_0_0_7_cascade_ ));
    InMux I__3460 (
            .O(N__17199),
            .I(N__17196));
    LocalMux I__3459 (
            .O(N__17196),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_7 ));
    InMux I__3458 (
            .O(N__17193),
            .I(N__17189));
    InMux I__3457 (
            .O(N__17192),
            .I(N__17185));
    LocalMux I__3456 (
            .O(N__17189),
            .I(N__17178));
    InMux I__3455 (
            .O(N__17188),
            .I(N__17175));
    LocalMux I__3454 (
            .O(N__17185),
            .I(N__17172));
    InMux I__3453 (
            .O(N__17184),
            .I(N__17169));
    InMux I__3452 (
            .O(N__17183),
            .I(N__17162));
    InMux I__3451 (
            .O(N__17182),
            .I(N__17162));
    InMux I__3450 (
            .O(N__17181),
            .I(N__17162));
    Odrv4 I__3449 (
            .O(N__17178),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__3448 (
            .O(N__17175),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    Odrv4 I__3447 (
            .O(N__17172),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__3446 (
            .O(N__17169),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__3445 (
            .O(N__17162),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__3444 (
            .O(N__17151),
            .I(N__17148));
    InMux I__3443 (
            .O(N__17148),
            .I(N__17144));
    InMux I__3442 (
            .O(N__17147),
            .I(N__17141));
    LocalMux I__3441 (
            .O(N__17144),
            .I(N__17138));
    LocalMux I__3440 (
            .O(N__17141),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    Odrv12 I__3439 (
            .O(N__17138),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__3438 (
            .O(N__17133),
            .I(N__17130));
    LocalMux I__3437 (
            .O(N__17130),
            .I(\ppm_encoder_1.un2_throttle_iv_0_rn_0_7 ));
    InMux I__3436 (
            .O(N__17127),
            .I(N__17124));
    LocalMux I__3435 (
            .O(N__17124),
            .I(N__17121));
    Span4Mux_v I__3434 (
            .O(N__17121),
            .I(N__17118));
    Span4Mux_h I__3433 (
            .O(N__17118),
            .I(N__17115));
    Odrv4 I__3432 (
            .O(N__17115),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__3431 (
            .O(N__17112),
            .I(N__17109));
    LocalMux I__3430 (
            .O(N__17109),
            .I(N__17106));
    Span4Mux_h I__3429 (
            .O(N__17106),
            .I(N__17102));
    InMux I__3428 (
            .O(N__17105),
            .I(N__17099));
    Span4Mux_h I__3427 (
            .O(N__17102),
            .I(N__17096));
    LocalMux I__3426 (
            .O(N__17099),
            .I(N__17093));
    Odrv4 I__3425 (
            .O(N__17096),
            .I(scaler_2_data_7));
    Odrv4 I__3424 (
            .O(N__17093),
            .I(scaler_2_data_7));
    InMux I__3423 (
            .O(N__17088),
            .I(N__17082));
    InMux I__3422 (
            .O(N__17087),
            .I(N__17082));
    LocalMux I__3421 (
            .O(N__17082),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    CascadeMux I__3420 (
            .O(N__17079),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ));
    InMux I__3419 (
            .O(N__17076),
            .I(N__17073));
    LocalMux I__3418 (
            .O(N__17073),
            .I(N__17070));
    Odrv4 I__3417 (
            .O(N__17070),
            .I(\ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1 ));
    InMux I__3416 (
            .O(N__17067),
            .I(N__17064));
    LocalMux I__3415 (
            .O(N__17064),
            .I(\ppm_encoder_1.N_426 ));
    InMux I__3414 (
            .O(N__17061),
            .I(N__17055));
    InMux I__3413 (
            .O(N__17060),
            .I(N__17052));
    InMux I__3412 (
            .O(N__17059),
            .I(N__17046));
    InMux I__3411 (
            .O(N__17058),
            .I(N__17041));
    LocalMux I__3410 (
            .O(N__17055),
            .I(N__17038));
    LocalMux I__3409 (
            .O(N__17052),
            .I(N__17033));
    InMux I__3408 (
            .O(N__17051),
            .I(N__17030));
    InMux I__3407 (
            .O(N__17050),
            .I(N__17024));
    InMux I__3406 (
            .O(N__17049),
            .I(N__17021));
    LocalMux I__3405 (
            .O(N__17046),
            .I(N__17018));
    InMux I__3404 (
            .O(N__17045),
            .I(N__17015));
    InMux I__3403 (
            .O(N__17044),
            .I(N__17012));
    LocalMux I__3402 (
            .O(N__17041),
            .I(N__17007));
    Span4Mux_v I__3401 (
            .O(N__17038),
            .I(N__17007));
    InMux I__3400 (
            .O(N__17037),
            .I(N__17002));
    InMux I__3399 (
            .O(N__17036),
            .I(N__17002));
    Span4Mux_v I__3398 (
            .O(N__17033),
            .I(N__16997));
    LocalMux I__3397 (
            .O(N__17030),
            .I(N__16997));
    InMux I__3396 (
            .O(N__17029),
            .I(N__16994));
    InMux I__3395 (
            .O(N__17028),
            .I(N__16989));
    InMux I__3394 (
            .O(N__17027),
            .I(N__16989));
    LocalMux I__3393 (
            .O(N__17024),
            .I(N__16984));
    LocalMux I__3392 (
            .O(N__17021),
            .I(N__16984));
    Span4Mux_h I__3391 (
            .O(N__17018),
            .I(N__16981));
    LocalMux I__3390 (
            .O(N__17015),
            .I(\ppm_encoder_1.N_246 ));
    LocalMux I__3389 (
            .O(N__17012),
            .I(\ppm_encoder_1.N_246 ));
    Odrv4 I__3388 (
            .O(N__17007),
            .I(\ppm_encoder_1.N_246 ));
    LocalMux I__3387 (
            .O(N__17002),
            .I(\ppm_encoder_1.N_246 ));
    Odrv4 I__3386 (
            .O(N__16997),
            .I(\ppm_encoder_1.N_246 ));
    LocalMux I__3385 (
            .O(N__16994),
            .I(\ppm_encoder_1.N_246 ));
    LocalMux I__3384 (
            .O(N__16989),
            .I(\ppm_encoder_1.N_246 ));
    Odrv4 I__3383 (
            .O(N__16984),
            .I(\ppm_encoder_1.N_246 ));
    Odrv4 I__3382 (
            .O(N__16981),
            .I(\ppm_encoder_1.N_246 ));
    CascadeMux I__3381 (
            .O(N__16962),
            .I(\ppm_encoder_1.N_426_cascade_ ));
    CascadeMux I__3380 (
            .O(N__16959),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    InMux I__3379 (
            .O(N__16956),
            .I(N__16953));
    LocalMux I__3378 (
            .O(N__16953),
            .I(N__16950));
    Odrv4 I__3377 (
            .O(N__16950),
            .I(\ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3 ));
    InMux I__3376 (
            .O(N__16947),
            .I(N__16944));
    LocalMux I__3375 (
            .O(N__16944),
            .I(N__16941));
    Span4Mux_v I__3374 (
            .O(N__16941),
            .I(N__16938));
    Odrv4 I__3373 (
            .O(N__16938),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__3372 (
            .O(N__16935),
            .I(N__16932));
    LocalMux I__3371 (
            .O(N__16932),
            .I(N__16929));
    Span4Mux_v I__3370 (
            .O(N__16929),
            .I(N__16926));
    Odrv4 I__3369 (
            .O(N__16926),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    CascadeMux I__3368 (
            .O(N__16923),
            .I(N__16915));
    CascadeMux I__3367 (
            .O(N__16922),
            .I(N__16911));
    CascadeMux I__3366 (
            .O(N__16921),
            .I(N__16907));
    CascadeMux I__3365 (
            .O(N__16920),
            .I(N__16904));
    CascadeMux I__3364 (
            .O(N__16919),
            .I(N__16901));
    InMux I__3363 (
            .O(N__16918),
            .I(N__16896));
    InMux I__3362 (
            .O(N__16915),
            .I(N__16896));
    InMux I__3361 (
            .O(N__16914),
            .I(N__16889));
    InMux I__3360 (
            .O(N__16911),
            .I(N__16889));
    InMux I__3359 (
            .O(N__16910),
            .I(N__16889));
    InMux I__3358 (
            .O(N__16907),
            .I(N__16882));
    InMux I__3357 (
            .O(N__16904),
            .I(N__16882));
    InMux I__3356 (
            .O(N__16901),
            .I(N__16882));
    LocalMux I__3355 (
            .O(N__16896),
            .I(N__16872));
    LocalMux I__3354 (
            .O(N__16889),
            .I(N__16867));
    LocalMux I__3353 (
            .O(N__16882),
            .I(N__16867));
    CascadeMux I__3352 (
            .O(N__16881),
            .I(N__16864));
    CascadeMux I__3351 (
            .O(N__16880),
            .I(N__16860));
    CascadeMux I__3350 (
            .O(N__16879),
            .I(N__16857));
    CascadeMux I__3349 (
            .O(N__16878),
            .I(N__16854));
    CascadeMux I__3348 (
            .O(N__16877),
            .I(N__16850));
    CascadeMux I__3347 (
            .O(N__16876),
            .I(N__16847));
    CascadeMux I__3346 (
            .O(N__16875),
            .I(N__16844));
    Span4Mux_v I__3345 (
            .O(N__16872),
            .I(N__16838));
    Span4Mux_h I__3344 (
            .O(N__16867),
            .I(N__16838));
    InMux I__3343 (
            .O(N__16864),
            .I(N__16833));
    InMux I__3342 (
            .O(N__16863),
            .I(N__16833));
    InMux I__3341 (
            .O(N__16860),
            .I(N__16826));
    InMux I__3340 (
            .O(N__16857),
            .I(N__16826));
    InMux I__3339 (
            .O(N__16854),
            .I(N__16826));
    InMux I__3338 (
            .O(N__16853),
            .I(N__16823));
    InMux I__3337 (
            .O(N__16850),
            .I(N__16816));
    InMux I__3336 (
            .O(N__16847),
            .I(N__16816));
    InMux I__3335 (
            .O(N__16844),
            .I(N__16816));
    InMux I__3334 (
            .O(N__16843),
            .I(N__16813));
    Odrv4 I__3333 (
            .O(N__16838),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__3332 (
            .O(N__16833),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__3331 (
            .O(N__16826),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__3330 (
            .O(N__16823),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__3329 (
            .O(N__16816),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__3328 (
            .O(N__16813),
            .I(\ppm_encoder_1.N_241 ));
    CascadeMux I__3327 (
            .O(N__16800),
            .I(N__16783));
    InMux I__3326 (
            .O(N__16799),
            .I(N__16767));
    InMux I__3325 (
            .O(N__16798),
            .I(N__16767));
    InMux I__3324 (
            .O(N__16797),
            .I(N__16767));
    InMux I__3323 (
            .O(N__16796),
            .I(N__16767));
    InMux I__3322 (
            .O(N__16795),
            .I(N__16767));
    InMux I__3321 (
            .O(N__16794),
            .I(N__16767));
    InMux I__3320 (
            .O(N__16793),
            .I(N__16762));
    InMux I__3319 (
            .O(N__16792),
            .I(N__16762));
    InMux I__3318 (
            .O(N__16791),
            .I(N__16759));
    InMux I__3317 (
            .O(N__16790),
            .I(N__16748));
    InMux I__3316 (
            .O(N__16789),
            .I(N__16748));
    InMux I__3315 (
            .O(N__16788),
            .I(N__16748));
    InMux I__3314 (
            .O(N__16787),
            .I(N__16748));
    InMux I__3313 (
            .O(N__16786),
            .I(N__16748));
    InMux I__3312 (
            .O(N__16783),
            .I(N__16739));
    InMux I__3311 (
            .O(N__16782),
            .I(N__16739));
    InMux I__3310 (
            .O(N__16781),
            .I(N__16739));
    InMux I__3309 (
            .O(N__16780),
            .I(N__16739));
    LocalMux I__3308 (
            .O(N__16767),
            .I(N__16736));
    LocalMux I__3307 (
            .O(N__16762),
            .I(N__16733));
    LocalMux I__3306 (
            .O(N__16759),
            .I(\ppm_encoder_1.N_348 ));
    LocalMux I__3305 (
            .O(N__16748),
            .I(\ppm_encoder_1.N_348 ));
    LocalMux I__3304 (
            .O(N__16739),
            .I(\ppm_encoder_1.N_348 ));
    Odrv4 I__3303 (
            .O(N__16736),
            .I(\ppm_encoder_1.N_348 ));
    Odrv12 I__3302 (
            .O(N__16733),
            .I(\ppm_encoder_1.N_348 ));
    InMux I__3301 (
            .O(N__16722),
            .I(N__16719));
    LocalMux I__3300 (
            .O(N__16719),
            .I(N__16716));
    Span4Mux_v I__3299 (
            .O(N__16716),
            .I(N__16713));
    Odrv4 I__3298 (
            .O(N__16713),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__3297 (
            .O(N__16710),
            .I(N__16707));
    LocalMux I__3296 (
            .O(N__16707),
            .I(N__16704));
    Span12Mux_v I__3295 (
            .O(N__16704),
            .I(N__16701));
    Odrv12 I__3294 (
            .O(N__16701),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__3293 (
            .O(N__16698),
            .I(N__16695));
    LocalMux I__3292 (
            .O(N__16695),
            .I(N__16692));
    Span4Mux_h I__3291 (
            .O(N__16692),
            .I(N__16689));
    Span4Mux_v I__3290 (
            .O(N__16689),
            .I(N__16685));
    InMux I__3289 (
            .O(N__16688),
            .I(N__16682));
    Span4Mux_h I__3288 (
            .O(N__16685),
            .I(N__16677));
    LocalMux I__3287 (
            .O(N__16682),
            .I(N__16677));
    Odrv4 I__3286 (
            .O(N__16677),
            .I(scaler_4_data_8));
    InMux I__3285 (
            .O(N__16674),
            .I(N__16671));
    LocalMux I__3284 (
            .O(N__16671),
            .I(N__16668));
    Span4Mux_h I__3283 (
            .O(N__16668),
            .I(N__16665));
    Span4Mux_v I__3282 (
            .O(N__16665),
            .I(N__16662));
    Span4Mux_v I__3281 (
            .O(N__16662),
            .I(N__16659));
    Odrv4 I__3280 (
            .O(N__16659),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__3279 (
            .O(N__16656),
            .I(N__16653));
    LocalMux I__3278 (
            .O(N__16653),
            .I(N__16650));
    Span12Mux_v I__3277 (
            .O(N__16650),
            .I(N__16646));
    InMux I__3276 (
            .O(N__16649),
            .I(N__16643));
    Odrv12 I__3275 (
            .O(N__16646),
            .I(scaler_1_data_7));
    LocalMux I__3274 (
            .O(N__16643),
            .I(scaler_1_data_7));
    InMux I__3273 (
            .O(N__16638),
            .I(N__16635));
    LocalMux I__3272 (
            .O(N__16635),
            .I(N__16632));
    Sp12to4 I__3271 (
            .O(N__16632),
            .I(N__16629));
    Span12Mux_v I__3270 (
            .O(N__16629),
            .I(N__16626));
    Odrv12 I__3269 (
            .O(N__16626),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__3268 (
            .O(N__16623),
            .I(N__16620));
    LocalMux I__3267 (
            .O(N__16620),
            .I(N__16617));
    Span4Mux_h I__3266 (
            .O(N__16617),
            .I(N__16614));
    Span4Mux_v I__3265 (
            .O(N__16614),
            .I(N__16610));
    InMux I__3264 (
            .O(N__16613),
            .I(N__16607));
    Span4Mux_h I__3263 (
            .O(N__16610),
            .I(N__16602));
    LocalMux I__3262 (
            .O(N__16607),
            .I(N__16602));
    Odrv4 I__3261 (
            .O(N__16602),
            .I(scaler_4_data_7));
    CascadeMux I__3260 (
            .O(N__16599),
            .I(\ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_ ));
    InMux I__3259 (
            .O(N__16596),
            .I(N__16593));
    LocalMux I__3258 (
            .O(N__16593),
            .I(N__16590));
    Odrv4 I__3257 (
            .O(N__16590),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__3256 (
            .O(N__16587),
            .I(N__16584));
    LocalMux I__3255 (
            .O(N__16584),
            .I(N__16581));
    Odrv4 I__3254 (
            .O(N__16581),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__3253 (
            .O(N__16578),
            .I(N__16575));
    LocalMux I__3252 (
            .O(N__16575),
            .I(N__16572));
    Odrv4 I__3251 (
            .O(N__16572),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__3250 (
            .O(N__16569),
            .I(N__16566));
    LocalMux I__3249 (
            .O(N__16566),
            .I(N__16563));
    Span4Mux_v I__3248 (
            .O(N__16563),
            .I(N__16560));
    Odrv4 I__3247 (
            .O(N__16560),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    CascadeMux I__3246 (
            .O(N__16557),
            .I(N__16554));
    InMux I__3245 (
            .O(N__16554),
            .I(N__16551));
    LocalMux I__3244 (
            .O(N__16551),
            .I(N__16548));
    Span4Mux_v I__3243 (
            .O(N__16548),
            .I(N__16545));
    Odrv4 I__3242 (
            .O(N__16545),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__3241 (
            .O(N__16542),
            .I(N__16539));
    LocalMux I__3240 (
            .O(N__16539),
            .I(N__16536));
    Span4Mux_v I__3239 (
            .O(N__16536),
            .I(N__16533));
    Odrv4 I__3238 (
            .O(N__16533),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__3237 (
            .O(N__16530),
            .I(N__16527));
    LocalMux I__3236 (
            .O(N__16527),
            .I(N__16524));
    Span4Mux_v I__3235 (
            .O(N__16524),
            .I(N__16521));
    Odrv4 I__3234 (
            .O(N__16521),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_13 ));
    InMux I__3233 (
            .O(N__16518),
            .I(N__16515));
    LocalMux I__3232 (
            .O(N__16515),
            .I(N__16512));
    Odrv4 I__3231 (
            .O(N__16512),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__3230 (
            .O(N__16509),
            .I(N__16506));
    LocalMux I__3229 (
            .O(N__16506),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__3228 (
            .O(N__16503),
            .I(N__16500));
    LocalMux I__3227 (
            .O(N__16500),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__3226 (
            .O(N__16497),
            .I(N__16494));
    LocalMux I__3225 (
            .O(N__16494),
            .I(N__16491));
    Span4Mux_v I__3224 (
            .O(N__16491),
            .I(N__16488));
    Odrv4 I__3223 (
            .O(N__16488),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__3222 (
            .O(N__16485),
            .I(N__16482));
    LocalMux I__3221 (
            .O(N__16482),
            .I(N__16479));
    Odrv4 I__3220 (
            .O(N__16479),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__3219 (
            .O(N__16476),
            .I(N__16473));
    LocalMux I__3218 (
            .O(N__16473),
            .I(N__16469));
    InMux I__3217 (
            .O(N__16472),
            .I(N__16466));
    Odrv4 I__3216 (
            .O(N__16469),
            .I(\ppm_encoder_1.N_245_i_i ));
    LocalMux I__3215 (
            .O(N__16466),
            .I(\ppm_encoder_1.N_245_i_i ));
    InMux I__3214 (
            .O(N__16461),
            .I(N__16458));
    LocalMux I__3213 (
            .O(N__16458),
            .I(N__16455));
    Span4Mux_v I__3212 (
            .O(N__16455),
            .I(N__16452));
    Odrv4 I__3211 (
            .O(N__16452),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__3210 (
            .O(N__16449),
            .I(N__16445));
    CascadeMux I__3209 (
            .O(N__16448),
            .I(N__16442));
    LocalMux I__3208 (
            .O(N__16445),
            .I(N__16439));
    InMux I__3207 (
            .O(N__16442),
            .I(N__16436));
    Span4Mux_h I__3206 (
            .O(N__16439),
            .I(N__16433));
    LocalMux I__3205 (
            .O(N__16436),
            .I(\ppm_encoder_1.N_251_i_i ));
    Odrv4 I__3204 (
            .O(N__16433),
            .I(\ppm_encoder_1.N_251_i_i ));
    InMux I__3203 (
            .O(N__16428),
            .I(N__16425));
    LocalMux I__3202 (
            .O(N__16425),
            .I(N__16422));
    Odrv12 I__3201 (
            .O(N__16422),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CascadeMux I__3200 (
            .O(N__16419),
            .I(N__16416));
    InMux I__3199 (
            .O(N__16416),
            .I(N__16413));
    LocalMux I__3198 (
            .O(N__16413),
            .I(N__16410));
    Span4Mux_h I__3197 (
            .O(N__16410),
            .I(N__16407));
    Odrv4 I__3196 (
            .O(N__16407),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    InMux I__3195 (
            .O(N__16404),
            .I(N__16401));
    LocalMux I__3194 (
            .O(N__16401),
            .I(\ppm_encoder_1.pulses2count_9_i_o2_0_14 ));
    InMux I__3193 (
            .O(N__16398),
            .I(N__16395));
    LocalMux I__3192 (
            .O(N__16395),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_12 ));
    CascadeMux I__3191 (
            .O(N__16392),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ));
    InMux I__3190 (
            .O(N__16389),
            .I(N__16386));
    LocalMux I__3189 (
            .O(N__16386),
            .I(\ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12 ));
    CascadeMux I__3188 (
            .O(N__16383),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_ ));
    InMux I__3187 (
            .O(N__16380),
            .I(N__16377));
    LocalMux I__3186 (
            .O(N__16377),
            .I(\ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7 ));
    CascadeMux I__3185 (
            .O(N__16374),
            .I(N__16371));
    InMux I__3184 (
            .O(N__16371),
            .I(N__16367));
    InMux I__3183 (
            .O(N__16370),
            .I(N__16364));
    LocalMux I__3182 (
            .O(N__16367),
            .I(N__16360));
    LocalMux I__3181 (
            .O(N__16364),
            .I(N__16357));
    CascadeMux I__3180 (
            .O(N__16363),
            .I(N__16354));
    Span4Mux_h I__3179 (
            .O(N__16360),
            .I(N__16351));
    Span4Mux_v I__3178 (
            .O(N__16357),
            .I(N__16348));
    InMux I__3177 (
            .O(N__16354),
            .I(N__16345));
    Odrv4 I__3176 (
            .O(N__16351),
            .I(\ppm_encoder_1.N_114 ));
    Odrv4 I__3175 (
            .O(N__16348),
            .I(\ppm_encoder_1.N_114 ));
    LocalMux I__3174 (
            .O(N__16345),
            .I(\ppm_encoder_1.N_114 ));
    InMux I__3173 (
            .O(N__16338),
            .I(N__16335));
    LocalMux I__3172 (
            .O(N__16335),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_12 ));
    CascadeMux I__3171 (
            .O(N__16332),
            .I(\ppm_encoder_1.N_407_cascade_ ));
    CascadeMux I__3170 (
            .O(N__16329),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_ ));
    CascadeMux I__3169 (
            .O(N__16326),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    InMux I__3168 (
            .O(N__16323),
            .I(N__16320));
    LocalMux I__3167 (
            .O(N__16320),
            .I(\ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2 ));
    InMux I__3166 (
            .O(N__16317),
            .I(N__16314));
    LocalMux I__3165 (
            .O(N__16314),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_14 ));
    CascadeMux I__3164 (
            .O(N__16311),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ));
    InMux I__3163 (
            .O(N__16308),
            .I(N__16305));
    LocalMux I__3162 (
            .O(N__16305),
            .I(\ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5 ));
    InMux I__3161 (
            .O(N__16302),
            .I(N__16299));
    LocalMux I__3160 (
            .O(N__16299),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0 ));
    InMux I__3159 (
            .O(N__16296),
            .I(N__16293));
    LocalMux I__3158 (
            .O(N__16293),
            .I(N__16290));
    Odrv12 I__3157 (
            .O(N__16290),
            .I(scaler_2_data_5));
    InMux I__3156 (
            .O(N__16287),
            .I(N__16284));
    LocalMux I__3155 (
            .O(N__16284),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__3154 (
            .O(N__16281),
            .I(N__16278));
    LocalMux I__3153 (
            .O(N__16278),
            .I(N__16275));
    Span4Mux_h I__3152 (
            .O(N__16275),
            .I(N__16272));
    Span4Mux_h I__3151 (
            .O(N__16272),
            .I(N__16269));
    Odrv4 I__3150 (
            .O(N__16269),
            .I(scaler_4_data_5));
    CEMux I__3149 (
            .O(N__16266),
            .I(N__16263));
    LocalMux I__3148 (
            .O(N__16263),
            .I(N__16258));
    CEMux I__3147 (
            .O(N__16262),
            .I(N__16255));
    CEMux I__3146 (
            .O(N__16261),
            .I(N__16250));
    IoSpan4Mux I__3145 (
            .O(N__16258),
            .I(N__16245));
    LocalMux I__3144 (
            .O(N__16255),
            .I(N__16245));
    CEMux I__3143 (
            .O(N__16254),
            .I(N__16240));
    CEMux I__3142 (
            .O(N__16253),
            .I(N__16237));
    LocalMux I__3141 (
            .O(N__16250),
            .I(N__16234));
    Span4Mux_s1_v I__3140 (
            .O(N__16245),
            .I(N__16231));
    CEMux I__3139 (
            .O(N__16244),
            .I(N__16228));
    CEMux I__3138 (
            .O(N__16243),
            .I(N__16225));
    LocalMux I__3137 (
            .O(N__16240),
            .I(N__16222));
    LocalMux I__3136 (
            .O(N__16237),
            .I(N__16215));
    Span4Mux_v I__3135 (
            .O(N__16234),
            .I(N__16215));
    Span4Mux_v I__3134 (
            .O(N__16231),
            .I(N__16215));
    LocalMux I__3133 (
            .O(N__16228),
            .I(N__16212));
    LocalMux I__3132 (
            .O(N__16225),
            .I(N__16209));
    Span4Mux_v I__3131 (
            .O(N__16222),
            .I(N__16206));
    Span4Mux_h I__3130 (
            .O(N__16215),
            .I(N__16203));
    Span4Mux_v I__3129 (
            .O(N__16212),
            .I(N__16200));
    Span4Mux_h I__3128 (
            .O(N__16209),
            .I(N__16193));
    Span4Mux_h I__3127 (
            .O(N__16206),
            .I(N__16193));
    Span4Mux_v I__3126 (
            .O(N__16203),
            .I(N__16193));
    Odrv4 I__3125 (
            .O(N__16200),
            .I(\ppm_encoder_1.scaler_1_dv_0 ));
    Odrv4 I__3124 (
            .O(N__16193),
            .I(\ppm_encoder_1.scaler_1_dv_0 ));
    CascadeMux I__3123 (
            .O(N__16188),
            .I(N__16185));
    InMux I__3122 (
            .O(N__16185),
            .I(N__16181));
    InMux I__3121 (
            .O(N__16184),
            .I(N__16178));
    LocalMux I__3120 (
            .O(N__16181),
            .I(\ppm_encoder_1.N_252_i_i ));
    LocalMux I__3119 (
            .O(N__16178),
            .I(\ppm_encoder_1.N_252_i_i ));
    InMux I__3118 (
            .O(N__16173),
            .I(N__16170));
    LocalMux I__3117 (
            .O(N__16170),
            .I(N__16167));
    Odrv4 I__3116 (
            .O(N__16167),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_8 ));
    InMux I__3115 (
            .O(N__16164),
            .I(N__16161));
    LocalMux I__3114 (
            .O(N__16161),
            .I(\ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8 ));
    CascadeMux I__3113 (
            .O(N__16158),
            .I(\ppm_encoder_1.N_235_cascade_ ));
    InMux I__3112 (
            .O(N__16155),
            .I(N__16152));
    LocalMux I__3111 (
            .O(N__16152),
            .I(N__16149));
    Span4Mux_h I__3110 (
            .O(N__16149),
            .I(N__16146));
    Span4Mux_v I__3109 (
            .O(N__16146),
            .I(N__16143));
    Odrv4 I__3108 (
            .O(N__16143),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__3107 (
            .O(N__16140),
            .I(N__16137));
    LocalMux I__3106 (
            .O(N__16137),
            .I(N__16134));
    Span4Mux_v I__3105 (
            .O(N__16134),
            .I(N__16130));
    InMux I__3104 (
            .O(N__16133),
            .I(N__16127));
    Span4Mux_v I__3103 (
            .O(N__16130),
            .I(N__16124));
    LocalMux I__3102 (
            .O(N__16127),
            .I(N__16121));
    Span4Mux_h I__3101 (
            .O(N__16124),
            .I(N__16116));
    Span4Mux_v I__3100 (
            .O(N__16121),
            .I(N__16116));
    Odrv4 I__3099 (
            .O(N__16116),
            .I(scaler_3_data_8));
    InMux I__3098 (
            .O(N__16113),
            .I(N__16110));
    LocalMux I__3097 (
            .O(N__16110),
            .I(N__16107));
    Span4Mux_h I__3096 (
            .O(N__16107),
            .I(N__16104));
    Span4Mux_h I__3095 (
            .O(N__16104),
            .I(N__16101));
    Odrv4 I__3094 (
            .O(N__16101),
            .I(scaler_3_data_5));
    InMux I__3093 (
            .O(N__16098),
            .I(N__16095));
    LocalMux I__3092 (
            .O(N__16095),
            .I(N__16092));
    Span4Mux_h I__3091 (
            .O(N__16092),
            .I(N__16088));
    CascadeMux I__3090 (
            .O(N__16091),
            .I(N__16085));
    Span4Mux_h I__3089 (
            .O(N__16088),
            .I(N__16082));
    InMux I__3088 (
            .O(N__16085),
            .I(N__16079));
    Odrv4 I__3087 (
            .O(N__16082),
            .I(scaler_4_data_4));
    LocalMux I__3086 (
            .O(N__16079),
            .I(scaler_4_data_4));
    InMux I__3085 (
            .O(N__16074),
            .I(N__16071));
    LocalMux I__3084 (
            .O(N__16071),
            .I(N__16068));
    Span4Mux_h I__3083 (
            .O(N__16068),
            .I(N__16064));
    CascadeMux I__3082 (
            .O(N__16067),
            .I(N__16061));
    Span4Mux_h I__3081 (
            .O(N__16064),
            .I(N__16058));
    InMux I__3080 (
            .O(N__16061),
            .I(N__16055));
    Odrv4 I__3079 (
            .O(N__16058),
            .I(scaler_1_data_4));
    LocalMux I__3078 (
            .O(N__16055),
            .I(scaler_1_data_4));
    InMux I__3077 (
            .O(N__16050),
            .I(N__16047));
    LocalMux I__3076 (
            .O(N__16047),
            .I(N__16044));
    Span12Mux_h I__3075 (
            .O(N__16044),
            .I(N__16041));
    Odrv12 I__3074 (
            .O(N__16041),
            .I(scaler_1_data_5));
    CascadeMux I__3073 (
            .O(N__16038),
            .I(N__16035));
    InMux I__3072 (
            .O(N__16035),
            .I(N__16032));
    LocalMux I__3071 (
            .O(N__16032),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    CascadeMux I__3070 (
            .O(N__16029),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_ ));
    CascadeMux I__3069 (
            .O(N__16026),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_ ));
    InMux I__3068 (
            .O(N__16023),
            .I(N__16020));
    LocalMux I__3067 (
            .O(N__16020),
            .I(N__16017));
    Span4Mux_h I__3066 (
            .O(N__16017),
            .I(N__16013));
    InMux I__3065 (
            .O(N__16016),
            .I(N__16010));
    Odrv4 I__3064 (
            .O(N__16013),
            .I(scaler_1_data_11));
    LocalMux I__3063 (
            .O(N__16010),
            .I(scaler_1_data_11));
    InMux I__3062 (
            .O(N__16005),
            .I(N__16002));
    LocalMux I__3061 (
            .O(N__16002),
            .I(N__15999));
    Odrv4 I__3060 (
            .O(N__15999),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__3059 (
            .O(N__15996),
            .I(N__15993));
    LocalMux I__3058 (
            .O(N__15993),
            .I(N__15989));
    CascadeMux I__3057 (
            .O(N__15992),
            .I(N__15986));
    Span4Mux_v I__3056 (
            .O(N__15989),
            .I(N__15983));
    InMux I__3055 (
            .O(N__15986),
            .I(N__15980));
    Span4Mux_h I__3054 (
            .O(N__15983),
            .I(N__15975));
    LocalMux I__3053 (
            .O(N__15980),
            .I(N__15975));
    Odrv4 I__3052 (
            .O(N__15975),
            .I(scaler_2_data_12));
    InMux I__3051 (
            .O(N__15972),
            .I(N__15969));
    LocalMux I__3050 (
            .O(N__15969),
            .I(N__15966));
    Span4Mux_v I__3049 (
            .O(N__15966),
            .I(N__15963));
    Span4Mux_h I__3048 (
            .O(N__15963),
            .I(N__15960));
    Odrv4 I__3047 (
            .O(N__15960),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__3046 (
            .O(N__15957),
            .I(N__15954));
    LocalMux I__3045 (
            .O(N__15954),
            .I(\ppm_encoder_1.N_418 ));
    CascadeMux I__3044 (
            .O(N__15951),
            .I(\ppm_encoder_1.N_417_cascade_ ));
    CascadeMux I__3043 (
            .O(N__15948),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_ ));
    InMux I__3042 (
            .O(N__15945),
            .I(N__15942));
    LocalMux I__3041 (
            .O(N__15942),
            .I(N__15939));
    Span4Mux_h I__3040 (
            .O(N__15939),
            .I(N__15936));
    Odrv4 I__3039 (
            .O(N__15936),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__3038 (
            .O(N__15933),
            .I(N__15930));
    LocalMux I__3037 (
            .O(N__15930),
            .I(N__15926));
    InMux I__3036 (
            .O(N__15929),
            .I(N__15923));
    Span12Mux_h I__3035 (
            .O(N__15926),
            .I(N__15920));
    LocalMux I__3034 (
            .O(N__15923),
            .I(N__15917));
    Odrv12 I__3033 (
            .O(N__15920),
            .I(scaler_2_data_8));
    Odrv4 I__3032 (
            .O(N__15917),
            .I(scaler_2_data_8));
    InMux I__3031 (
            .O(N__15912),
            .I(N__15909));
    LocalMux I__3030 (
            .O(N__15909),
            .I(N__15906));
    Span4Mux_h I__3029 (
            .O(N__15906),
            .I(N__15903));
    Span4Mux_v I__3028 (
            .O(N__15903),
            .I(N__15900));
    Span4Mux_v I__3027 (
            .O(N__15900),
            .I(N__15897));
    Odrv4 I__3026 (
            .O(N__15897),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    CascadeMux I__3025 (
            .O(N__15894),
            .I(N__15891));
    InMux I__3024 (
            .O(N__15891),
            .I(N__15888));
    LocalMux I__3023 (
            .O(N__15888),
            .I(N__15885));
    Span4Mux_h I__3022 (
            .O(N__15885),
            .I(N__15882));
    Span4Mux_v I__3021 (
            .O(N__15882),
            .I(N__15879));
    Span4Mux_h I__3020 (
            .O(N__15879),
            .I(N__15875));
    InMux I__3019 (
            .O(N__15878),
            .I(N__15872));
    Odrv4 I__3018 (
            .O(N__15875),
            .I(scaler_1_data_8));
    LocalMux I__3017 (
            .O(N__15872),
            .I(scaler_1_data_8));
    CascadeMux I__3016 (
            .O(N__15867),
            .I(N__15863));
    InMux I__3015 (
            .O(N__15866),
            .I(N__15860));
    InMux I__3014 (
            .O(N__15863),
            .I(N__15857));
    LocalMux I__3013 (
            .O(N__15860),
            .I(N__15854));
    LocalMux I__3012 (
            .O(N__15857),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__3011 (
            .O(N__15854),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    CascadeMux I__3010 (
            .O(N__15849),
            .I(\ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_ ));
    InMux I__3009 (
            .O(N__15846),
            .I(N__15843));
    LocalMux I__3008 (
            .O(N__15843),
            .I(N__15840));
    Span4Mux_v I__3007 (
            .O(N__15840),
            .I(N__15836));
    InMux I__3006 (
            .O(N__15839),
            .I(N__15833));
    Span4Mux_h I__3005 (
            .O(N__15836),
            .I(N__15830));
    LocalMux I__3004 (
            .O(N__15833),
            .I(N__15827));
    Odrv4 I__3003 (
            .O(N__15830),
            .I(scaler_2_data_13));
    Odrv4 I__3002 (
            .O(N__15827),
            .I(scaler_2_data_13));
    InMux I__3001 (
            .O(N__15822),
            .I(N__15819));
    LocalMux I__3000 (
            .O(N__15819),
            .I(N__15816));
    Span4Mux_s3_v I__2999 (
            .O(N__15816),
            .I(N__15813));
    Span4Mux_h I__2998 (
            .O(N__15813),
            .I(N__15810));
    Odrv4 I__2997 (
            .O(N__15810),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__2996 (
            .O(N__15807),
            .I(N__15801));
    InMux I__2995 (
            .O(N__15806),
            .I(N__15801));
    LocalMux I__2994 (
            .O(N__15801),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    CascadeMux I__2993 (
            .O(N__15798),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ));
    CascadeMux I__2992 (
            .O(N__15795),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ));
    CascadeMux I__2991 (
            .O(N__15792),
            .I(N__15789));
    InMux I__2990 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__2989 (
            .O(N__15786),
            .I(N__15783));
    Odrv12 I__2988 (
            .O(N__15783),
            .I(\ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13 ));
    InMux I__2987 (
            .O(N__15780),
            .I(N__15777));
    LocalMux I__2986 (
            .O(N__15777),
            .I(N__15773));
    InMux I__2985 (
            .O(N__15776),
            .I(N__15770));
    Span4Mux_h I__2984 (
            .O(N__15773),
            .I(N__15767));
    LocalMux I__2983 (
            .O(N__15770),
            .I(N__15764));
    Span4Mux_h I__2982 (
            .O(N__15767),
            .I(N__15761));
    Span4Mux_h I__2981 (
            .O(N__15764),
            .I(N__15758));
    Odrv4 I__2980 (
            .O(N__15761),
            .I(scaler_3_data_13));
    Odrv4 I__2979 (
            .O(N__15758),
            .I(scaler_3_data_13));
    InMux I__2978 (
            .O(N__15753),
            .I(N__15750));
    LocalMux I__2977 (
            .O(N__15750),
            .I(N__15747));
    Span4Mux_h I__2976 (
            .O(N__15747),
            .I(N__15744));
    Odrv4 I__2975 (
            .O(N__15744),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    CascadeMux I__2974 (
            .O(N__15741),
            .I(N__15737));
    InMux I__2973 (
            .O(N__15740),
            .I(N__15732));
    InMux I__2972 (
            .O(N__15737),
            .I(N__15732));
    LocalMux I__2971 (
            .O(N__15732),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__2970 (
            .O(N__15729),
            .I(N__15726));
    LocalMux I__2969 (
            .O(N__15726),
            .I(N__15723));
    Odrv12 I__2968 (
            .O(N__15723),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_11 ));
    InMux I__2967 (
            .O(N__15720),
            .I(N__15717));
    LocalMux I__2966 (
            .O(N__15717),
            .I(N__15713));
    InMux I__2965 (
            .O(N__15716),
            .I(N__15710));
    Span4Mux_h I__2964 (
            .O(N__15713),
            .I(N__15707));
    LocalMux I__2963 (
            .O(N__15710),
            .I(N__15704));
    Span4Mux_v I__2962 (
            .O(N__15707),
            .I(N__15701));
    Span4Mux_h I__2961 (
            .O(N__15704),
            .I(N__15698));
    Odrv4 I__2960 (
            .O(N__15701),
            .I(scaler_3_data_11));
    Odrv4 I__2959 (
            .O(N__15698),
            .I(scaler_3_data_11));
    CascadeMux I__2958 (
            .O(N__15693),
            .I(N__15690));
    InMux I__2957 (
            .O(N__15690),
            .I(N__15687));
    LocalMux I__2956 (
            .O(N__15687),
            .I(N__15684));
    Span4Mux_s3_v I__2955 (
            .O(N__15684),
            .I(N__15681));
    Odrv4 I__2954 (
            .O(N__15681),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    CascadeMux I__2953 (
            .O(N__15678),
            .I(\ppm_encoder_1.N_114_cascade_ ));
    InMux I__2952 (
            .O(N__15675),
            .I(N__15670));
    InMux I__2951 (
            .O(N__15674),
            .I(N__15667));
    InMux I__2950 (
            .O(N__15673),
            .I(N__15664));
    LocalMux I__2949 (
            .O(N__15670),
            .I(N__15661));
    LocalMux I__2948 (
            .O(N__15667),
            .I(N__15658));
    LocalMux I__2947 (
            .O(N__15664),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__2946 (
            .O(N__15661),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__2945 (
            .O(N__15658),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    CascadeMux I__2944 (
            .O(N__15651),
            .I(N__15646));
    CascadeMux I__2943 (
            .O(N__15650),
            .I(N__15643));
    InMux I__2942 (
            .O(N__15649),
            .I(N__15640));
    InMux I__2941 (
            .O(N__15646),
            .I(N__15637));
    InMux I__2940 (
            .O(N__15643),
            .I(N__15634));
    LocalMux I__2939 (
            .O(N__15640),
            .I(N__15629));
    LocalMux I__2938 (
            .O(N__15637),
            .I(N__15629));
    LocalMux I__2937 (
            .O(N__15634),
            .I(N__15626));
    Odrv4 I__2936 (
            .O(N__15629),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__2935 (
            .O(N__15626),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    CascadeMux I__2934 (
            .O(N__15621),
            .I(\ppm_encoder_1.N_348_cascade_ ));
    InMux I__2933 (
            .O(N__15618),
            .I(N__15615));
    LocalMux I__2932 (
            .O(N__15615),
            .I(N__15612));
    Odrv4 I__2931 (
            .O(N__15612),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    CascadeMux I__2930 (
            .O(N__15609),
            .I(\ppm_encoder_1.init_pulses_18_i_0_14_cascade_ ));
    InMux I__2929 (
            .O(N__15606),
            .I(N__15603));
    LocalMux I__2928 (
            .O(N__15603),
            .I(\ppm_encoder_1.init_pulses_18_i_a2_0_14 ));
    InMux I__2927 (
            .O(N__15600),
            .I(N__15597));
    LocalMux I__2926 (
            .O(N__15597),
            .I(N__15594));
    Odrv4 I__2925 (
            .O(N__15594),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    CascadeMux I__2924 (
            .O(N__15591),
            .I(\ppm_encoder_1.N_241_cascade_ ));
    CascadeMux I__2923 (
            .O(N__15588),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ));
    CascadeMux I__2922 (
            .O(N__15585),
            .I(N__15582));
    InMux I__2921 (
            .O(N__15582),
            .I(N__15579));
    LocalMux I__2920 (
            .O(N__15579),
            .I(\ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14 ));
    CascadeMux I__2919 (
            .O(N__15576),
            .I(N__15573));
    InMux I__2918 (
            .O(N__15573),
            .I(N__15570));
    LocalMux I__2917 (
            .O(N__15570),
            .I(N__15567));
    Odrv4 I__2916 (
            .O(N__15567),
            .I(\ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15 ));
    InMux I__2915 (
            .O(N__15564),
            .I(N__15561));
    LocalMux I__2914 (
            .O(N__15561),
            .I(N__15558));
    Span4Mux_v I__2913 (
            .O(N__15558),
            .I(N__15555));
    Odrv4 I__2912 (
            .O(N__15555),
            .I(\ppm_encoder_1.N_403 ));
    CascadeMux I__2911 (
            .O(N__15552),
            .I(N__15549));
    InMux I__2910 (
            .O(N__15549),
            .I(N__15546));
    LocalMux I__2909 (
            .O(N__15546),
            .I(N__15543));
    Span4Mux_h I__2908 (
            .O(N__15543),
            .I(N__15540));
    Odrv4 I__2907 (
            .O(N__15540),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    InMux I__2906 (
            .O(N__15537),
            .I(N__15534));
    LocalMux I__2905 (
            .O(N__15534),
            .I(N__15531));
    Odrv12 I__2904 (
            .O(N__15531),
            .I(\ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10 ));
    InMux I__2903 (
            .O(N__15528),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__2902 (
            .O(N__15525),
            .I(N__15522));
    LocalMux I__2901 (
            .O(N__15522),
            .I(N__15519));
    Odrv12 I__2900 (
            .O(N__15519),
            .I(\ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11 ));
    InMux I__2899 (
            .O(N__15516),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__2898 (
            .O(N__15513),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__2897 (
            .O(N__15510),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__2896 (
            .O(N__15507),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__2895 (
            .O(N__15504),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__2894 (
            .O(N__15501),
            .I(bfn_7_25_0_));
    InMux I__2893 (
            .O(N__15498),
            .I(N__15495));
    LocalMux I__2892 (
            .O(N__15495),
            .I(N__15492));
    Odrv12 I__2891 (
            .O(N__15492),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__2890 (
            .O(N__15489),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__2889 (
            .O(N__15486),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__2888 (
            .O(N__15483),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__2887 (
            .O(N__15480),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__2886 (
            .O(N__15477),
            .I(N__15474));
    LocalMux I__2885 (
            .O(N__15474),
            .I(\ppm_encoder_1.init_pulses_RNI398E4Z0Z_4 ));
    InMux I__2884 (
            .O(N__15471),
            .I(N__15468));
    LocalMux I__2883 (
            .O(N__15468),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__2882 (
            .O(N__15465),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__2881 (
            .O(N__15462),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__2880 (
            .O(N__15459),
            .I(N__15456));
    LocalMux I__2879 (
            .O(N__15456),
            .I(N__15453));
    Odrv4 I__2878 (
            .O(N__15453),
            .I(\ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6 ));
    InMux I__2877 (
            .O(N__15450),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__2876 (
            .O(N__15447),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__2875 (
            .O(N__15444),
            .I(bfn_7_24_0_));
    InMux I__2874 (
            .O(N__15441),
            .I(N__15438));
    LocalMux I__2873 (
            .O(N__15438),
            .I(N__15435));
    Odrv4 I__2872 (
            .O(N__15435),
            .I(\ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9 ));
    InMux I__2871 (
            .O(N__15432),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    CascadeMux I__2870 (
            .O(N__15429),
            .I(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ));
    InMux I__2869 (
            .O(N__15426),
            .I(N__15423));
    LocalMux I__2868 (
            .O(N__15423),
            .I(\ppm_encoder_1.un2_throttle_iv_i_i_1_4 ));
    CascadeMux I__2867 (
            .O(N__15420),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ));
    InMux I__2866 (
            .O(N__15417),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__2865 (
            .O(N__15414),
            .I(N__15411));
    LocalMux I__2864 (
            .O(N__15411),
            .I(N__15407));
    IoInMux I__2863 (
            .O(N__15410),
            .I(N__15404));
    Span4Mux_h I__2862 (
            .O(N__15407),
            .I(N__15401));
    LocalMux I__2861 (
            .O(N__15404),
            .I(N__15398));
    Span4Mux_v I__2860 (
            .O(N__15401),
            .I(N__15395));
    IoSpan4Mux I__2859 (
            .O(N__15398),
            .I(N__15392));
    Odrv4 I__2858 (
            .O(N__15395),
            .I(uart_input_c));
    Odrv4 I__2857 (
            .O(N__15392),
            .I(uart_input_c));
    InMux I__2856 (
            .O(N__15387),
            .I(N__15384));
    LocalMux I__2855 (
            .O(N__15384),
            .I(N__15381));
    Span4Mux_v I__2854 (
            .O(N__15381),
            .I(N__15378));
    Odrv4 I__2853 (
            .O(N__15378),
            .I(\uart_sync.aux_0__0_Z0Z_0 ));
    InMux I__2852 (
            .O(N__15375),
            .I(N__15372));
    LocalMux I__2851 (
            .O(N__15372),
            .I(N__15368));
    InMux I__2850 (
            .O(N__15371),
            .I(N__15364));
    Span4Mux_h I__2849 (
            .O(N__15368),
            .I(N__15361));
    InMux I__2848 (
            .O(N__15367),
            .I(N__15358));
    LocalMux I__2847 (
            .O(N__15364),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__2846 (
            .O(N__15361),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    LocalMux I__2845 (
            .O(N__15358),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    CascadeMux I__2844 (
            .O(N__15351),
            .I(N__15348));
    InMux I__2843 (
            .O(N__15348),
            .I(N__15345));
    LocalMux I__2842 (
            .O(N__15345),
            .I(N__15342));
    Span4Mux_h I__2841 (
            .O(N__15342),
            .I(N__15339));
    Odrv4 I__2840 (
            .O(N__15339),
            .I(\ppm_encoder_1.pulses2count_9_0_o2_0_6 ));
    CascadeMux I__2839 (
            .O(N__15336),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ));
    InMux I__2838 (
            .O(N__15333),
            .I(N__15330));
    LocalMux I__2837 (
            .O(N__15330),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_11 ));
    CascadeMux I__2836 (
            .O(N__15327),
            .I(\ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_ ));
    InMux I__2835 (
            .O(N__15324),
            .I(N__15321));
    LocalMux I__2834 (
            .O(N__15321),
            .I(N__15318));
    Odrv4 I__2833 (
            .O(N__15318),
            .I(\ppm_encoder_1.N_462 ));
    InMux I__2832 (
            .O(N__15315),
            .I(N__15312));
    LocalMux I__2831 (
            .O(N__15312),
            .I(N__15307));
    InMux I__2830 (
            .O(N__15311),
            .I(N__15302));
    InMux I__2829 (
            .O(N__15310),
            .I(N__15302));
    Odrv4 I__2828 (
            .O(N__15307),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__2827 (
            .O(N__15302),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    InMux I__2826 (
            .O(N__15297),
            .I(N__15294));
    LocalMux I__2825 (
            .O(N__15294),
            .I(N__15291));
    Odrv4 I__2824 (
            .O(N__15291),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__2823 (
            .O(N__15288),
            .I(N__15285));
    LocalMux I__2822 (
            .O(N__15285),
            .I(N__15281));
    InMux I__2821 (
            .O(N__15284),
            .I(N__15278));
    Span4Mux_v I__2820 (
            .O(N__15281),
            .I(N__15275));
    LocalMux I__2819 (
            .O(N__15278),
            .I(N__15272));
    Odrv4 I__2818 (
            .O(N__15275),
            .I(scaler_4_data_9));
    Odrv4 I__2817 (
            .O(N__15272),
            .I(scaler_4_data_9));
    InMux I__2816 (
            .O(N__15267),
            .I(N__15263));
    InMux I__2815 (
            .O(N__15266),
            .I(N__15260));
    LocalMux I__2814 (
            .O(N__15263),
            .I(N__15257));
    LocalMux I__2813 (
            .O(N__15260),
            .I(N__15254));
    Span4Mux_v I__2812 (
            .O(N__15257),
            .I(N__15251));
    Span4Mux_h I__2811 (
            .O(N__15254),
            .I(N__15248));
    Odrv4 I__2810 (
            .O(N__15251),
            .I(scaler_3_data_10));
    Odrv4 I__2809 (
            .O(N__15248),
            .I(scaler_3_data_10));
    InMux I__2808 (
            .O(N__15243),
            .I(N__15240));
    LocalMux I__2807 (
            .O(N__15240),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__2806 (
            .O(N__15237),
            .I(N__15234));
    LocalMux I__2805 (
            .O(N__15234),
            .I(N__15231));
    Span4Mux_v I__2804 (
            .O(N__15231),
            .I(N__15226));
    InMux I__2803 (
            .O(N__15230),
            .I(N__15223));
    InMux I__2802 (
            .O(N__15229),
            .I(N__15219));
    Span4Mux_v I__2801 (
            .O(N__15226),
            .I(N__15214));
    LocalMux I__2800 (
            .O(N__15223),
            .I(N__15214));
    CascadeMux I__2799 (
            .O(N__15222),
            .I(N__15211));
    LocalMux I__2798 (
            .O(N__15219),
            .I(N__15208));
    Span4Mux_h I__2797 (
            .O(N__15214),
            .I(N__15205));
    InMux I__2796 (
            .O(N__15211),
            .I(N__15202));
    Odrv4 I__2795 (
            .O(N__15208),
            .I(frame_decoder_OFF2data_0));
    Odrv4 I__2794 (
            .O(N__15205),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__2793 (
            .O(N__15202),
            .I(frame_decoder_OFF2data_0));
    InMux I__2792 (
            .O(N__15195),
            .I(N__15191));
    InMux I__2791 (
            .O(N__15194),
            .I(N__15188));
    LocalMux I__2790 (
            .O(N__15191),
            .I(N__15185));
    LocalMux I__2789 (
            .O(N__15188),
            .I(N__15181));
    Span4Mux_v I__2788 (
            .O(N__15185),
            .I(N__15178));
    InMux I__2787 (
            .O(N__15184),
            .I(N__15175));
    Span4Mux_h I__2786 (
            .O(N__15181),
            .I(N__15171));
    Span4Mux_h I__2785 (
            .O(N__15178),
            .I(N__15168));
    LocalMux I__2784 (
            .O(N__15175),
            .I(N__15165));
    InMux I__2783 (
            .O(N__15174),
            .I(N__15162));
    Odrv4 I__2782 (
            .O(N__15171),
            .I(frame_decoder_CH2data_0));
    Odrv4 I__2781 (
            .O(N__15168),
            .I(frame_decoder_CH2data_0));
    Odrv12 I__2780 (
            .O(N__15165),
            .I(frame_decoder_CH2data_0));
    LocalMux I__2779 (
            .O(N__15162),
            .I(frame_decoder_CH2data_0));
    InMux I__2778 (
            .O(N__15153),
            .I(N__15149));
    CascadeMux I__2777 (
            .O(N__15152),
            .I(N__15146));
    LocalMux I__2776 (
            .O(N__15149),
            .I(N__15143));
    InMux I__2775 (
            .O(N__15146),
            .I(N__15140));
    Odrv12 I__2774 (
            .O(N__15143),
            .I(scaler_2_data_4));
    LocalMux I__2773 (
            .O(N__15140),
            .I(scaler_2_data_4));
    InMux I__2772 (
            .O(N__15135),
            .I(N__15131));
    InMux I__2771 (
            .O(N__15134),
            .I(N__15128));
    LocalMux I__2770 (
            .O(N__15131),
            .I(N__15123));
    LocalMux I__2769 (
            .O(N__15128),
            .I(N__15123));
    Span4Mux_h I__2768 (
            .O(N__15123),
            .I(N__15120));
    Odrv4 I__2767 (
            .O(N__15120),
            .I(scaler_4_data_12));
    InMux I__2766 (
            .O(N__15117),
            .I(N__15114));
    LocalMux I__2765 (
            .O(N__15114),
            .I(N__15111));
    Odrv4 I__2764 (
            .O(N__15111),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__2763 (
            .O(N__15108),
            .I(N__15102));
    InMux I__2762 (
            .O(N__15107),
            .I(N__15099));
    InMux I__2761 (
            .O(N__15106),
            .I(N__15096));
    InMux I__2760 (
            .O(N__15105),
            .I(N__15090));
    LocalMux I__2759 (
            .O(N__15102),
            .I(N__15083));
    LocalMux I__2758 (
            .O(N__15099),
            .I(N__15083));
    LocalMux I__2757 (
            .O(N__15096),
            .I(N__15083));
    InMux I__2756 (
            .O(N__15095),
            .I(N__15080));
    InMux I__2755 (
            .O(N__15094),
            .I(N__15077));
    InMux I__2754 (
            .O(N__15093),
            .I(N__15074));
    LocalMux I__2753 (
            .O(N__15090),
            .I(N__15070));
    Span4Mux_v I__2752 (
            .O(N__15083),
            .I(N__15061));
    LocalMux I__2751 (
            .O(N__15080),
            .I(N__15061));
    LocalMux I__2750 (
            .O(N__15077),
            .I(N__15061));
    LocalMux I__2749 (
            .O(N__15074),
            .I(N__15061));
    InMux I__2748 (
            .O(N__15073),
            .I(N__15058));
    Span4Mux_v I__2747 (
            .O(N__15070),
            .I(N__15053));
    Span4Mux_v I__2746 (
            .O(N__15061),
            .I(N__15048));
    LocalMux I__2745 (
            .O(N__15058),
            .I(N__15048));
    InMux I__2744 (
            .O(N__15057),
            .I(N__15045));
    InMux I__2743 (
            .O(N__15056),
            .I(N__15042));
    Odrv4 I__2742 (
            .O(N__15053),
            .I(uart_data_4));
    Odrv4 I__2741 (
            .O(N__15048),
            .I(uart_data_4));
    LocalMux I__2740 (
            .O(N__15045),
            .I(uart_data_4));
    LocalMux I__2739 (
            .O(N__15042),
            .I(uart_data_4));
    InMux I__2738 (
            .O(N__15033),
            .I(N__15030));
    LocalMux I__2737 (
            .O(N__15030),
            .I(N__15027));
    Odrv4 I__2736 (
            .O(N__15027),
            .I(frame_decoder_CH1data_4));
    CEMux I__2735 (
            .O(N__15024),
            .I(N__15021));
    LocalMux I__2734 (
            .O(N__15021),
            .I(N__15018));
    Span4Mux_v I__2733 (
            .O(N__15018),
            .I(N__15014));
    CEMux I__2732 (
            .O(N__15017),
            .I(N__15011));
    Span4Mux_h I__2731 (
            .O(N__15014),
            .I(N__15008));
    LocalMux I__2730 (
            .O(N__15011),
            .I(N__15005));
    Odrv4 I__2729 (
            .O(N__15008),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa_0 ));
    Odrv12 I__2728 (
            .O(N__15005),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa_0 ));
    InMux I__2727 (
            .O(N__15000),
            .I(N__14997));
    LocalMux I__2726 (
            .O(N__14997),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__2725 (
            .O(N__14994),
            .I(N__14991));
    LocalMux I__2724 (
            .O(N__14991),
            .I(N__14987));
    InMux I__2723 (
            .O(N__14990),
            .I(N__14984));
    Odrv12 I__2722 (
            .O(N__14987),
            .I(scaler_1_data_12));
    LocalMux I__2721 (
            .O(N__14984),
            .I(scaler_1_data_12));
    InMux I__2720 (
            .O(N__14979),
            .I(N__14976));
    LocalMux I__2719 (
            .O(N__14976),
            .I(N__14973));
    Span4Mux_v I__2718 (
            .O(N__14973),
            .I(N__14969));
    InMux I__2717 (
            .O(N__14972),
            .I(N__14966));
    Odrv4 I__2716 (
            .O(N__14969),
            .I(scaler_1_data_13));
    LocalMux I__2715 (
            .O(N__14966),
            .I(scaler_1_data_13));
    InMux I__2714 (
            .O(N__14961),
            .I(N__14958));
    LocalMux I__2713 (
            .O(N__14958),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    IoInMux I__2712 (
            .O(N__14955),
            .I(N__14952));
    LocalMux I__2711 (
            .O(N__14952),
            .I(N__14949));
    Span12Mux_s8_v I__2710 (
            .O(N__14949),
            .I(N__14943));
    InMux I__2709 (
            .O(N__14948),
            .I(N__14940));
    InMux I__2708 (
            .O(N__14947),
            .I(N__14934));
    InMux I__2707 (
            .O(N__14946),
            .I(N__14934));
    Span12Mux_h I__2706 (
            .O(N__14943),
            .I(N__14929));
    LocalMux I__2705 (
            .O(N__14940),
            .I(N__14926));
    InMux I__2704 (
            .O(N__14939),
            .I(N__14923));
    LocalMux I__2703 (
            .O(N__14934),
            .I(N__14920));
    InMux I__2702 (
            .O(N__14933),
            .I(N__14917));
    CascadeMux I__2701 (
            .O(N__14932),
            .I(N__14913));
    Span12Mux_v I__2700 (
            .O(N__14929),
            .I(N__14906));
    Sp12to4 I__2699 (
            .O(N__14926),
            .I(N__14906));
    LocalMux I__2698 (
            .O(N__14923),
            .I(N__14906));
    Span4Mux_h I__2697 (
            .O(N__14920),
            .I(N__14901));
    LocalMux I__2696 (
            .O(N__14917),
            .I(N__14901));
    InMux I__2695 (
            .O(N__14916),
            .I(N__14896));
    InMux I__2694 (
            .O(N__14913),
            .I(N__14896));
    Span12Mux_s9_v I__2693 (
            .O(N__14906),
            .I(N__14893));
    Odrv4 I__2692 (
            .O(N__14901),
            .I(frame_decoder_dv_c));
    LocalMux I__2691 (
            .O(N__14896),
            .I(frame_decoder_dv_c));
    Odrv12 I__2690 (
            .O(N__14893),
            .I(frame_decoder_dv_c));
    IoInMux I__2689 (
            .O(N__14886),
            .I(N__14883));
    LocalMux I__2688 (
            .O(N__14883),
            .I(frame_decoder_dv_c_0));
    InMux I__2687 (
            .O(N__14880),
            .I(N__14877));
    LocalMux I__2686 (
            .O(N__14877),
            .I(\ppm_encoder_1.N_415 ));
    CascadeMux I__2685 (
            .O(N__14874),
            .I(\ppm_encoder_1.N_414_cascade_ ));
    CascadeMux I__2684 (
            .O(N__14871),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_ ));
    CascadeMux I__2683 (
            .O(N__14868),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ));
    CascadeMux I__2682 (
            .O(N__14865),
            .I(N__14861));
    CascadeMux I__2681 (
            .O(N__14864),
            .I(N__14858));
    InMux I__2680 (
            .O(N__14861),
            .I(N__14855));
    InMux I__2679 (
            .O(N__14858),
            .I(N__14851));
    LocalMux I__2678 (
            .O(N__14855),
            .I(N__14848));
    InMux I__2677 (
            .O(N__14854),
            .I(N__14845));
    LocalMux I__2676 (
            .O(N__14851),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    Odrv12 I__2675 (
            .O(N__14848),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__2674 (
            .O(N__14845),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__2673 (
            .O(N__14838),
            .I(N__14835));
    LocalMux I__2672 (
            .O(N__14835),
            .I(\ppm_encoder_1.N_412 ));
    CascadeMux I__2671 (
            .O(N__14832),
            .I(\ppm_encoder_1.N_411_cascade_ ));
    CascadeMux I__2670 (
            .O(N__14829),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_ ));
    InMux I__2669 (
            .O(N__14826),
            .I(N__14823));
    LocalMux I__2668 (
            .O(N__14823),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_9 ));
    InMux I__2667 (
            .O(N__14820),
            .I(N__14817));
    LocalMux I__2666 (
            .O(N__14817),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__2665 (
            .O(N__14814),
            .I(N__14811));
    LocalMux I__2664 (
            .O(N__14811),
            .I(N__14807));
    InMux I__2663 (
            .O(N__14810),
            .I(N__14804));
    Span4Mux_v I__2662 (
            .O(N__14807),
            .I(N__14801));
    LocalMux I__2661 (
            .O(N__14804),
            .I(N__14798));
    Odrv4 I__2660 (
            .O(N__14801),
            .I(scaler_2_data_9));
    Odrv4 I__2659 (
            .O(N__14798),
            .I(scaler_2_data_9));
    InMux I__2658 (
            .O(N__14793),
            .I(N__14789));
    InMux I__2657 (
            .O(N__14792),
            .I(N__14786));
    LocalMux I__2656 (
            .O(N__14789),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    LocalMux I__2655 (
            .O(N__14786),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__2654 (
            .O(N__14781),
            .I(N__14777));
    InMux I__2653 (
            .O(N__14780),
            .I(N__14774));
    LocalMux I__2652 (
            .O(N__14777),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    LocalMux I__2651 (
            .O(N__14774),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__2650 (
            .O(N__14769),
            .I(N__14766));
    LocalMux I__2649 (
            .O(N__14766),
            .I(N__14762));
    InMux I__2648 (
            .O(N__14765),
            .I(N__14759));
    Span4Mux_h I__2647 (
            .O(N__14762),
            .I(N__14754));
    LocalMux I__2646 (
            .O(N__14759),
            .I(N__14754));
    Span4Mux_v I__2645 (
            .O(N__14754),
            .I(N__14751));
    Odrv4 I__2644 (
            .O(N__14751),
            .I(scaler_2_data_6));
    InMux I__2643 (
            .O(N__14748),
            .I(N__14742));
    InMux I__2642 (
            .O(N__14747),
            .I(N__14742));
    LocalMux I__2641 (
            .O(N__14742),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    CascadeMux I__2640 (
            .O(N__14739),
            .I(N__14736));
    InMux I__2639 (
            .O(N__14736),
            .I(N__14732));
    InMux I__2638 (
            .O(N__14735),
            .I(N__14729));
    LocalMux I__2637 (
            .O(N__14732),
            .I(N__14726));
    LocalMux I__2636 (
            .O(N__14729),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    Odrv4 I__2635 (
            .O(N__14726),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    CascadeMux I__2634 (
            .O(N__14721),
            .I(\ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_ ));
    InMux I__2633 (
            .O(N__14718),
            .I(N__14715));
    LocalMux I__2632 (
            .O(N__14715),
            .I(\ppm_encoder_1.un2_throttle_iv_0_rn_0_6 ));
    CascadeMux I__2631 (
            .O(N__14712),
            .I(\ppm_encoder_1.un2_throttle_0_6_cascade_ ));
    CascadeMux I__2630 (
            .O(N__14709),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ));
    InMux I__2629 (
            .O(N__14706),
            .I(N__14703));
    LocalMux I__2628 (
            .O(N__14703),
            .I(\ppm_encoder_1.un2_throttle_iv_0_sn_6 ));
    InMux I__2627 (
            .O(N__14700),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__2626 (
            .O(N__14697),
            .I(N__14691));
    InMux I__2625 (
            .O(N__14696),
            .I(N__14691));
    LocalMux I__2624 (
            .O(N__14691),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__2623 (
            .O(N__14688),
            .I(N__14684));
    InMux I__2622 (
            .O(N__14687),
            .I(N__14681));
    LocalMux I__2621 (
            .O(N__14684),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__2620 (
            .O(N__14681),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__2619 (
            .O(N__14676),
            .I(N__14672));
    InMux I__2618 (
            .O(N__14675),
            .I(N__14667));
    InMux I__2617 (
            .O(N__14672),
            .I(N__14667));
    LocalMux I__2616 (
            .O(N__14667),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__2615 (
            .O(N__14664),
            .I(N__14660));
    InMux I__2614 (
            .O(N__14663),
            .I(N__14657));
    LocalMux I__2613 (
            .O(N__14660),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__2612 (
            .O(N__14657),
            .I(\reset_module_System.countZ0Z_13 ));
    CascadeMux I__2611 (
            .O(N__14652),
            .I(N__14649));
    InMux I__2610 (
            .O(N__14649),
            .I(N__14641));
    InMux I__2609 (
            .O(N__14648),
            .I(N__14641));
    InMux I__2608 (
            .O(N__14647),
            .I(N__14636));
    InMux I__2607 (
            .O(N__14646),
            .I(N__14636));
    LocalMux I__2606 (
            .O(N__14641),
            .I(N__14631));
    LocalMux I__2605 (
            .O(N__14636),
            .I(N__14631));
    Odrv4 I__2604 (
            .O(N__14631),
            .I(\reset_module_System.reset6_15 ));
    InMux I__2603 (
            .O(N__14628),
            .I(N__14625));
    LocalMux I__2602 (
            .O(N__14625),
            .I(N__14621));
    CascadeMux I__2601 (
            .O(N__14624),
            .I(N__14618));
    Span4Mux_v I__2600 (
            .O(N__14621),
            .I(N__14615));
    InMux I__2599 (
            .O(N__14618),
            .I(N__14612));
    Odrv4 I__2598 (
            .O(N__14615),
            .I(scaler_3_data_4));
    LocalMux I__2597 (
            .O(N__14612),
            .I(scaler_3_data_4));
    InMux I__2596 (
            .O(N__14607),
            .I(N__14603));
    CascadeMux I__2595 (
            .O(N__14606),
            .I(N__14599));
    LocalMux I__2594 (
            .O(N__14603),
            .I(N__14595));
    InMux I__2593 (
            .O(N__14602),
            .I(N__14592));
    InMux I__2592 (
            .O(N__14599),
            .I(N__14587));
    InMux I__2591 (
            .O(N__14598),
            .I(N__14587));
    Odrv4 I__2590 (
            .O(N__14595),
            .I(\scaler_2.un2_source_data_0 ));
    LocalMux I__2589 (
            .O(N__14592),
            .I(\scaler_2.un2_source_data_0 ));
    LocalMux I__2588 (
            .O(N__14587),
            .I(\scaler_2.un2_source_data_0 ));
    CascadeMux I__2587 (
            .O(N__14580),
            .I(N__14577));
    InMux I__2586 (
            .O(N__14577),
            .I(N__14574));
    LocalMux I__2585 (
            .O(N__14574),
            .I(N__14571));
    Odrv4 I__2584 (
            .O(N__14571),
            .I(\scaler_2.un2_source_data_0_cry_1_c_RNO_0 ));
    InMux I__2583 (
            .O(N__14568),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__2582 (
            .O(N__14565),
            .I(N__14561));
    InMux I__2581 (
            .O(N__14564),
            .I(N__14558));
    LocalMux I__2580 (
            .O(N__14561),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__2579 (
            .O(N__14558),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__2578 (
            .O(N__14553),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__2577 (
            .O(N__14550),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__2576 (
            .O(N__14547),
            .I(N__14543));
    InMux I__2575 (
            .O(N__14546),
            .I(N__14540));
    LocalMux I__2574 (
            .O(N__14543),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__2573 (
            .O(N__14540),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__2572 (
            .O(N__14535),
            .I(\reset_module_System.count_1_cry_15 ));
    CascadeMux I__2571 (
            .O(N__14532),
            .I(N__14528));
    InMux I__2570 (
            .O(N__14531),
            .I(N__14525));
    InMux I__2569 (
            .O(N__14528),
            .I(N__14522));
    LocalMux I__2568 (
            .O(N__14525),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__2567 (
            .O(N__14522),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__2566 (
            .O(N__14517),
            .I(bfn_5_19_0_));
    CascadeMux I__2565 (
            .O(N__14514),
            .I(N__14511));
    InMux I__2564 (
            .O(N__14511),
            .I(N__14507));
    InMux I__2563 (
            .O(N__14510),
            .I(N__14504));
    LocalMux I__2562 (
            .O(N__14507),
            .I(N__14501));
    LocalMux I__2561 (
            .O(N__14504),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__2560 (
            .O(N__14501),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__2559 (
            .O(N__14496),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__2558 (
            .O(N__14493),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__2557 (
            .O(N__14490),
            .I(N__14487));
    InMux I__2556 (
            .O(N__14487),
            .I(N__14483));
    InMux I__2555 (
            .O(N__14486),
            .I(N__14480));
    LocalMux I__2554 (
            .O(N__14483),
            .I(N__14477));
    LocalMux I__2553 (
            .O(N__14480),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__2552 (
            .O(N__14477),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__2551 (
            .O(N__14472),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__2550 (
            .O(N__14469),
            .I(N__14465));
    InMux I__2549 (
            .O(N__14468),
            .I(N__14462));
    LocalMux I__2548 (
            .O(N__14465),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__2547 (
            .O(N__14462),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__2546 (
            .O(N__14457),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__2545 (
            .O(N__14454),
            .I(N__14450));
    InMux I__2544 (
            .O(N__14453),
            .I(N__14447));
    LocalMux I__2543 (
            .O(N__14450),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__2542 (
            .O(N__14447),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__2541 (
            .O(N__14442),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__2540 (
            .O(N__14439),
            .I(N__14435));
    InMux I__2539 (
            .O(N__14438),
            .I(N__14432));
    LocalMux I__2538 (
            .O(N__14435),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__2537 (
            .O(N__14432),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__2536 (
            .O(N__14427),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__2535 (
            .O(N__14424),
            .I(N__14420));
    InMux I__2534 (
            .O(N__14423),
            .I(N__14417));
    LocalMux I__2533 (
            .O(N__14420),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__2532 (
            .O(N__14417),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__2531 (
            .O(N__14412),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__2530 (
            .O(N__14409),
            .I(N__14405));
    InMux I__2529 (
            .O(N__14408),
            .I(N__14402));
    LocalMux I__2528 (
            .O(N__14405),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__2527 (
            .O(N__14402),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__2526 (
            .O(N__14397),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__2525 (
            .O(N__14394),
            .I(N__14390));
    InMux I__2524 (
            .O(N__14393),
            .I(N__14387));
    InMux I__2523 (
            .O(N__14390),
            .I(N__14384));
    LocalMux I__2522 (
            .O(N__14387),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__2521 (
            .O(N__14384),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__2520 (
            .O(N__14379),
            .I(bfn_5_18_0_));
    InMux I__2519 (
            .O(N__14376),
            .I(N__14372));
    InMux I__2518 (
            .O(N__14375),
            .I(N__14369));
    LocalMux I__2517 (
            .O(N__14372),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__2516 (
            .O(N__14369),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__2515 (
            .O(N__14364),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__2514 (
            .O(N__14361),
            .I(N__14357));
    InMux I__2513 (
            .O(N__14360),
            .I(N__14354));
    LocalMux I__2512 (
            .O(N__14357),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__2511 (
            .O(N__14354),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__2510 (
            .O(N__14349),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__2509 (
            .O(N__14346),
            .I(N__14342));
    InMux I__2508 (
            .O(N__14345),
            .I(N__14339));
    LocalMux I__2507 (
            .O(N__14342),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__2506 (
            .O(N__14339),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__2505 (
            .O(N__14334),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__2504 (
            .O(N__14331),
            .I(\uart.un4_timer_Count_1_cry_3 ));
    CascadeMux I__2503 (
            .O(N__14328),
            .I(N__14321));
    InMux I__2502 (
            .O(N__14327),
            .I(N__14318));
    InMux I__2501 (
            .O(N__14326),
            .I(N__14311));
    InMux I__2500 (
            .O(N__14325),
            .I(N__14311));
    InMux I__2499 (
            .O(N__14324),
            .I(N__14311));
    InMux I__2498 (
            .O(N__14321),
            .I(N__14308));
    LocalMux I__2497 (
            .O(N__14318),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__2496 (
            .O(N__14311),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__2495 (
            .O(N__14308),
            .I(\uart.timer_CountZ0Z_5 ));
    InMux I__2494 (
            .O(N__14301),
            .I(\uart.un4_timer_Count_1_cry_4 ));
    InMux I__2493 (
            .O(N__14298),
            .I(N__14292));
    InMux I__2492 (
            .O(N__14297),
            .I(N__14292));
    LocalMux I__2491 (
            .O(N__14292),
            .I(N__14286));
    CascadeMux I__2490 (
            .O(N__14291),
            .I(N__14283));
    CascadeMux I__2489 (
            .O(N__14290),
            .I(N__14280));
    InMux I__2488 (
            .O(N__14289),
            .I(N__14276));
    Span4Mux_v I__2487 (
            .O(N__14286),
            .I(N__14273));
    InMux I__2486 (
            .O(N__14283),
            .I(N__14268));
    InMux I__2485 (
            .O(N__14280),
            .I(N__14268));
    InMux I__2484 (
            .O(N__14279),
            .I(N__14265));
    LocalMux I__2483 (
            .O(N__14276),
            .I(\uart.timer_CountZ0Z_6 ));
    Odrv4 I__2482 (
            .O(N__14273),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__2481 (
            .O(N__14268),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__2480 (
            .O(N__14265),
            .I(\uart.timer_CountZ0Z_6 ));
    InMux I__2479 (
            .O(N__14256),
            .I(\uart.un4_timer_Count_1_cry_5 ));
    InMux I__2478 (
            .O(N__14253),
            .I(\uart.un4_timer_Count_1_cry_6 ));
    InMux I__2477 (
            .O(N__14250),
            .I(N__14244));
    InMux I__2476 (
            .O(N__14249),
            .I(N__14241));
    InMux I__2475 (
            .O(N__14248),
            .I(N__14237));
    InMux I__2474 (
            .O(N__14247),
            .I(N__14234));
    LocalMux I__2473 (
            .O(N__14244),
            .I(N__14228));
    LocalMux I__2472 (
            .O(N__14241),
            .I(N__14228));
    InMux I__2471 (
            .O(N__14240),
            .I(N__14224));
    LocalMux I__2470 (
            .O(N__14237),
            .I(N__14219));
    LocalMux I__2469 (
            .O(N__14234),
            .I(N__14219));
    InMux I__2468 (
            .O(N__14233),
            .I(N__14214));
    Span4Mux_v I__2467 (
            .O(N__14228),
            .I(N__14211));
    InMux I__2466 (
            .O(N__14227),
            .I(N__14208));
    LocalMux I__2465 (
            .O(N__14224),
            .I(N__14205));
    Span4Mux_h I__2464 (
            .O(N__14219),
            .I(N__14202));
    InMux I__2463 (
            .O(N__14218),
            .I(N__14197));
    InMux I__2462 (
            .O(N__14217),
            .I(N__14197));
    LocalMux I__2461 (
            .O(N__14214),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__2460 (
            .O(N__14211),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__2459 (
            .O(N__14208),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__2458 (
            .O(N__14205),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__2457 (
            .O(N__14202),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__2456 (
            .O(N__14197),
            .I(\uart.timer_CountZ0Z_7 ));
    SRMux I__2455 (
            .O(N__14184),
            .I(N__14180));
    SRMux I__2454 (
            .O(N__14183),
            .I(N__14177));
    LocalMux I__2453 (
            .O(N__14180),
            .I(N__14173));
    LocalMux I__2452 (
            .O(N__14177),
            .I(N__14170));
    SRMux I__2451 (
            .O(N__14176),
            .I(N__14167));
    Span4Mux_v I__2450 (
            .O(N__14173),
            .I(N__14164));
    Span4Mux_v I__2449 (
            .O(N__14170),
            .I(N__14159));
    LocalMux I__2448 (
            .O(N__14167),
            .I(N__14159));
    Span4Mux_h I__2447 (
            .O(N__14164),
            .I(N__14156));
    Span4Mux_h I__2446 (
            .O(N__14159),
            .I(N__14153));
    Odrv4 I__2445 (
            .O(N__14156),
            .I(\uart.timer_Count_1_sqmuxa_i ));
    Odrv4 I__2444 (
            .O(N__14153),
            .I(\uart.timer_Count_1_sqmuxa_i ));
    CascadeMux I__2443 (
            .O(N__14148),
            .I(N__14145));
    InMux I__2442 (
            .O(N__14145),
            .I(N__14139));
    InMux I__2441 (
            .O(N__14144),
            .I(N__14136));
    InMux I__2440 (
            .O(N__14143),
            .I(N__14133));
    InMux I__2439 (
            .O(N__14142),
            .I(N__14130));
    LocalMux I__2438 (
            .O(N__14139),
            .I(N__14125));
    LocalMux I__2437 (
            .O(N__14136),
            .I(N__14125));
    LocalMux I__2436 (
            .O(N__14133),
            .I(\uart.timer_CountZ0Z_0 ));
    LocalMux I__2435 (
            .O(N__14130),
            .I(\uart.timer_CountZ0Z_0 ));
    Odrv4 I__2434 (
            .O(N__14125),
            .I(\uart.timer_CountZ0Z_0 ));
    InMux I__2433 (
            .O(N__14118),
            .I(N__14111));
    InMux I__2432 (
            .O(N__14117),
            .I(N__14108));
    InMux I__2431 (
            .O(N__14116),
            .I(N__14103));
    InMux I__2430 (
            .O(N__14115),
            .I(N__14103));
    InMux I__2429 (
            .O(N__14114),
            .I(N__14100));
    LocalMux I__2428 (
            .O(N__14111),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__2427 (
            .O(N__14108),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__2426 (
            .O(N__14103),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__2425 (
            .O(N__14100),
            .I(\uart.timer_CountZ0Z_4 ));
    InMux I__2424 (
            .O(N__14091),
            .I(N__14088));
    LocalMux I__2423 (
            .O(N__14088),
            .I(\uart.un1_state_2_0_a3_0 ));
    InMux I__2422 (
            .O(N__14085),
            .I(N__14082));
    LocalMux I__2421 (
            .O(N__14082),
            .I(N__14076));
    InMux I__2420 (
            .O(N__14081),
            .I(N__14073));
    InMux I__2419 (
            .O(N__14080),
            .I(N__14070));
    InMux I__2418 (
            .O(N__14079),
            .I(N__14067));
    Odrv4 I__2417 (
            .O(N__14076),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__2416 (
            .O(N__14073),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__2415 (
            .O(N__14070),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__2414 (
            .O(N__14067),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__2413 (
            .O(N__14058),
            .I(N__14053));
    CascadeMux I__2412 (
            .O(N__14057),
            .I(N__14050));
    InMux I__2411 (
            .O(N__14056),
            .I(N__14047));
    LocalMux I__2410 (
            .O(N__14053),
            .I(N__14044));
    InMux I__2409 (
            .O(N__14050),
            .I(N__14041));
    LocalMux I__2408 (
            .O(N__14047),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv12 I__2407 (
            .O(N__14044),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__2406 (
            .O(N__14041),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__2405 (
            .O(N__14034),
            .I(N__14030));
    InMux I__2404 (
            .O(N__14033),
            .I(N__14027));
    LocalMux I__2403 (
            .O(N__14030),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__2402 (
            .O(N__14027),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__2401 (
            .O(N__14022),
            .I(N__14019));
    LocalMux I__2400 (
            .O(N__14019),
            .I(\reset_module_System.count_1_2 ));
    InMux I__2399 (
            .O(N__14016),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__2398 (
            .O(N__14013),
            .I(N__14009));
    InMux I__2397 (
            .O(N__14012),
            .I(N__14006));
    LocalMux I__2396 (
            .O(N__14009),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__2395 (
            .O(N__14006),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__2394 (
            .O(N__14001),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__2393 (
            .O(N__13998),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__2392 (
            .O(N__13995),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__2391 (
            .O(N__13992),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__2390 (
            .O(N__13989),
            .I(N__13986));
    LocalMux I__2389 (
            .O(N__13986),
            .I(scaler_1_data_14));
    InMux I__2388 (
            .O(N__13983),
            .I(bfn_4_30_0_));
    InMux I__2387 (
            .O(N__13980),
            .I(N__13977));
    LocalMux I__2386 (
            .O(N__13977),
            .I(\uart_sync.aux_1__0_Z0Z_0 ));
    InMux I__2385 (
            .O(N__13974),
            .I(N__13969));
    InMux I__2384 (
            .O(N__13973),
            .I(N__13966));
    InMux I__2383 (
            .O(N__13972),
            .I(N__13963));
    LocalMux I__2382 (
            .O(N__13969),
            .I(N__13960));
    LocalMux I__2381 (
            .O(N__13966),
            .I(N__13957));
    LocalMux I__2380 (
            .O(N__13963),
            .I(\uart.timer_CountZ0Z_1 ));
    Odrv4 I__2379 (
            .O(N__13960),
            .I(\uart.timer_CountZ0Z_1 ));
    Odrv4 I__2378 (
            .O(N__13957),
            .I(\uart.timer_CountZ0Z_1 ));
    InMux I__2377 (
            .O(N__13950),
            .I(N__13944));
    InMux I__2376 (
            .O(N__13949),
            .I(N__13941));
    InMux I__2375 (
            .O(N__13948),
            .I(N__13936));
    InMux I__2374 (
            .O(N__13947),
            .I(N__13936));
    LocalMux I__2373 (
            .O(N__13944),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__2372 (
            .O(N__13941),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__2371 (
            .O(N__13936),
            .I(\uart.timer_CountZ0Z_2 ));
    InMux I__2370 (
            .O(N__13929),
            .I(\uart.un4_timer_Count_1_cry_1 ));
    CascadeMux I__2369 (
            .O(N__13926),
            .I(N__13921));
    InMux I__2368 (
            .O(N__13925),
            .I(N__13917));
    InMux I__2367 (
            .O(N__13924),
            .I(N__13914));
    InMux I__2366 (
            .O(N__13921),
            .I(N__13909));
    InMux I__2365 (
            .O(N__13920),
            .I(N__13909));
    LocalMux I__2364 (
            .O(N__13917),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__2363 (
            .O(N__13914),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__2362 (
            .O(N__13909),
            .I(\uart.timer_CountZ0Z_3 ));
    InMux I__2361 (
            .O(N__13902),
            .I(\uart.un4_timer_Count_1_cry_2 ));
    InMux I__2360 (
            .O(N__13899),
            .I(N__13895));
    InMux I__2359 (
            .O(N__13898),
            .I(N__13892));
    LocalMux I__2358 (
            .O(N__13895),
            .I(N__13889));
    LocalMux I__2357 (
            .O(N__13892),
            .I(N__13886));
    Span4Mux_h I__2356 (
            .O(N__13889),
            .I(N__13883));
    Span4Mux_h I__2355 (
            .O(N__13886),
            .I(N__13880));
    Odrv4 I__2354 (
            .O(N__13883),
            .I(scaler_3_data_12));
    Odrv4 I__2353 (
            .O(N__13880),
            .I(scaler_3_data_12));
    InMux I__2352 (
            .O(N__13875),
            .I(N__13872));
    LocalMux I__2351 (
            .O(N__13872),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__2350 (
            .O(N__13869),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__2349 (
            .O(N__13866),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__2348 (
            .O(N__13863),
            .I(N__13860));
    LocalMux I__2347 (
            .O(N__13860),
            .I(N__13857));
    Span4Mux_v I__2346 (
            .O(N__13857),
            .I(N__13854));
    Odrv4 I__2345 (
            .O(N__13854),
            .I(scaler_3_data_14));
    InMux I__2344 (
            .O(N__13851),
            .I(bfn_4_28_0_));
    InMux I__2343 (
            .O(N__13848),
            .I(N__13845));
    LocalMux I__2342 (
            .O(N__13845),
            .I(N__13842));
    Span4Mux_v I__2341 (
            .O(N__13842),
            .I(N__13838));
    InMux I__2340 (
            .O(N__13841),
            .I(N__13835));
    Odrv4 I__2339 (
            .O(N__13838),
            .I(scaler_1_data_6));
    LocalMux I__2338 (
            .O(N__13835),
            .I(scaler_1_data_6));
    InMux I__2337 (
            .O(N__13830),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__2336 (
            .O(N__13827),
            .I(\ppm_encoder_1.un1_throttle_cry_7 ));
    InMux I__2335 (
            .O(N__13824),
            .I(N__13821));
    LocalMux I__2334 (
            .O(N__13821),
            .I(N__13817));
    InMux I__2333 (
            .O(N__13820),
            .I(N__13814));
    Odrv4 I__2332 (
            .O(N__13817),
            .I(scaler_1_data_9));
    LocalMux I__2331 (
            .O(N__13814),
            .I(scaler_1_data_9));
    InMux I__2330 (
            .O(N__13809),
            .I(N__13806));
    LocalMux I__2329 (
            .O(N__13806),
            .I(N__13803));
    Odrv4 I__2328 (
            .O(N__13803),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__2327 (
            .O(N__13800),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__2326 (
            .O(N__13797),
            .I(N__13794));
    LocalMux I__2325 (
            .O(N__13794),
            .I(N__13790));
    InMux I__2324 (
            .O(N__13793),
            .I(N__13787));
    Odrv4 I__2323 (
            .O(N__13790),
            .I(scaler_1_data_10));
    LocalMux I__2322 (
            .O(N__13787),
            .I(scaler_1_data_10));
    InMux I__2321 (
            .O(N__13782),
            .I(N__13779));
    LocalMux I__2320 (
            .O(N__13779),
            .I(N__13776));
    Odrv4 I__2319 (
            .O(N__13776),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__2318 (
            .O(N__13773),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__2317 (
            .O(N__13770),
            .I(N__13766));
    InMux I__2316 (
            .O(N__13769),
            .I(N__13763));
    LocalMux I__2315 (
            .O(N__13766),
            .I(N__13760));
    LocalMux I__2314 (
            .O(N__13763),
            .I(N__13757));
    Span4Mux_h I__2313 (
            .O(N__13760),
            .I(N__13752));
    Span4Mux_h I__2312 (
            .O(N__13757),
            .I(N__13752));
    Odrv4 I__2311 (
            .O(N__13752),
            .I(scaler_3_data_6));
    InMux I__2310 (
            .O(N__13749),
            .I(N__13745));
    InMux I__2309 (
            .O(N__13748),
            .I(N__13742));
    LocalMux I__2308 (
            .O(N__13745),
            .I(N__13739));
    LocalMux I__2307 (
            .O(N__13742),
            .I(N__13736));
    Span4Mux_v I__2306 (
            .O(N__13739),
            .I(N__13731));
    Span4Mux_v I__2305 (
            .O(N__13736),
            .I(N__13731));
    Odrv4 I__2304 (
            .O(N__13731),
            .I(scaler_3_data_7));
    InMux I__2303 (
            .O(N__13728),
            .I(N__13725));
    LocalMux I__2302 (
            .O(N__13725),
            .I(N__13722));
    Odrv12 I__2301 (
            .O(N__13722),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__2300 (
            .O(N__13719),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__2299 (
            .O(N__13716),
            .I(\ppm_encoder_1.un1_elevator_cry_7 ));
    InMux I__2298 (
            .O(N__13713),
            .I(N__13710));
    LocalMux I__2297 (
            .O(N__13710),
            .I(N__13706));
    InMux I__2296 (
            .O(N__13709),
            .I(N__13703));
    Span4Mux_v I__2295 (
            .O(N__13706),
            .I(N__13698));
    LocalMux I__2294 (
            .O(N__13703),
            .I(N__13698));
    Span4Mux_h I__2293 (
            .O(N__13698),
            .I(N__13695));
    Odrv4 I__2292 (
            .O(N__13695),
            .I(scaler_3_data_9));
    InMux I__2291 (
            .O(N__13692),
            .I(N__13689));
    LocalMux I__2290 (
            .O(N__13689),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__2289 (
            .O(N__13686),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__2288 (
            .O(N__13683),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__2287 (
            .O(N__13680),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__2286 (
            .O(N__13677),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__2285 (
            .O(N__13674),
            .I(N__13670));
    InMux I__2284 (
            .O(N__13673),
            .I(N__13667));
    LocalMux I__2283 (
            .O(N__13670),
            .I(N__13662));
    LocalMux I__2282 (
            .O(N__13667),
            .I(N__13662));
    Span4Mux_v I__2281 (
            .O(N__13662),
            .I(N__13659));
    Odrv4 I__2280 (
            .O(N__13659),
            .I(scaler_2_data_11));
    InMux I__2279 (
            .O(N__13656),
            .I(N__13653));
    LocalMux I__2278 (
            .O(N__13653),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__2277 (
            .O(N__13650),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__2276 (
            .O(N__13647),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__2275 (
            .O(N__13644),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__2274 (
            .O(N__13641),
            .I(N__13638));
    LocalMux I__2273 (
            .O(N__13638),
            .I(N__13635));
    Span4Mux_v I__2272 (
            .O(N__13635),
            .I(N__13632));
    Odrv4 I__2271 (
            .O(N__13632),
            .I(scaler_2_data_14));
    InMux I__2270 (
            .O(N__13629),
            .I(bfn_4_25_0_));
    InMux I__2269 (
            .O(N__13626),
            .I(N__13623));
    LocalMux I__2268 (
            .O(N__13623),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__2267 (
            .O(N__13620),
            .I(N__13617));
    LocalMux I__2266 (
            .O(N__13617),
            .I(N__13613));
    CascadeMux I__2265 (
            .O(N__13616),
            .I(N__13610));
    Span4Mux_v I__2264 (
            .O(N__13613),
            .I(N__13607));
    InMux I__2263 (
            .O(N__13610),
            .I(N__13604));
    Span4Mux_s1_v I__2262 (
            .O(N__13607),
            .I(N__13601));
    LocalMux I__2261 (
            .O(N__13604),
            .I(N__13598));
    Odrv4 I__2260 (
            .O(N__13601),
            .I(scaler_4_data_10));
    Odrv4 I__2259 (
            .O(N__13598),
            .I(scaler_4_data_10));
    InMux I__2258 (
            .O(N__13593),
            .I(N__13590));
    LocalMux I__2257 (
            .O(N__13590),
            .I(N__13586));
    InMux I__2256 (
            .O(N__13589),
            .I(N__13583));
    Span4Mux_v I__2255 (
            .O(N__13586),
            .I(N__13580));
    LocalMux I__2254 (
            .O(N__13583),
            .I(N__13577));
    Odrv4 I__2253 (
            .O(N__13580),
            .I(scaler_2_data_10));
    Odrv4 I__2252 (
            .O(N__13577),
            .I(scaler_2_data_10));
    InMux I__2251 (
            .O(N__13572),
            .I(N__13569));
    LocalMux I__2250 (
            .O(N__13569),
            .I(N__13566));
    Odrv4 I__2249 (
            .O(N__13566),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__2248 (
            .O(N__13563),
            .I(N__13560));
    LocalMux I__2247 (
            .O(N__13560),
            .I(N__13556));
    InMux I__2246 (
            .O(N__13559),
            .I(N__13553));
    Span4Mux_h I__2245 (
            .O(N__13556),
            .I(N__13550));
    LocalMux I__2244 (
            .O(N__13553),
            .I(N__13547));
    Span4Mux_s2_h I__2243 (
            .O(N__13550),
            .I(N__13542));
    Span4Mux_h I__2242 (
            .O(N__13547),
            .I(N__13542));
    Odrv4 I__2241 (
            .O(N__13542),
            .I(scaler_4_data_13));
    InMux I__2240 (
            .O(N__13539),
            .I(N__13536));
    LocalMux I__2239 (
            .O(N__13536),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    InMux I__2238 (
            .O(N__13533),
            .I(N__13530));
    LocalMux I__2237 (
            .O(N__13530),
            .I(N__13527));
    Span4Mux_h I__2236 (
            .O(N__13527),
            .I(N__13523));
    InMux I__2235 (
            .O(N__13526),
            .I(N__13520));
    Span4Mux_v I__2234 (
            .O(N__13523),
            .I(N__13517));
    LocalMux I__2233 (
            .O(N__13520),
            .I(N__13514));
    Odrv4 I__2232 (
            .O(N__13517),
            .I(scaler_4_data_6));
    Odrv4 I__2231 (
            .O(N__13514),
            .I(scaler_4_data_6));
    InMux I__2230 (
            .O(N__13509),
            .I(N__13506));
    LocalMux I__2229 (
            .O(N__13506),
            .I(N__13500));
    InMux I__2228 (
            .O(N__13505),
            .I(N__13497));
    InMux I__2227 (
            .O(N__13504),
            .I(N__13494));
    CascadeMux I__2226 (
            .O(N__13503),
            .I(N__13491));
    Span4Mux_v I__2225 (
            .O(N__13500),
            .I(N__13486));
    LocalMux I__2224 (
            .O(N__13497),
            .I(N__13486));
    LocalMux I__2223 (
            .O(N__13494),
            .I(N__13483));
    InMux I__2222 (
            .O(N__13491),
            .I(N__13480));
    Odrv4 I__2221 (
            .O(N__13486),
            .I(frame_decoder_OFF3data_0));
    Odrv4 I__2220 (
            .O(N__13483),
            .I(frame_decoder_OFF3data_0));
    LocalMux I__2219 (
            .O(N__13480),
            .I(frame_decoder_OFF3data_0));
    InMux I__2218 (
            .O(N__13473),
            .I(N__13469));
    InMux I__2217 (
            .O(N__13472),
            .I(N__13466));
    LocalMux I__2216 (
            .O(N__13469),
            .I(N__13461));
    LocalMux I__2215 (
            .O(N__13466),
            .I(N__13461));
    Span4Mux_v I__2214 (
            .O(N__13461),
            .I(N__13456));
    InMux I__2213 (
            .O(N__13460),
            .I(N__13453));
    InMux I__2212 (
            .O(N__13459),
            .I(N__13450));
    Odrv4 I__2211 (
            .O(N__13456),
            .I(frame_decoder_CH3data_0));
    LocalMux I__2210 (
            .O(N__13453),
            .I(frame_decoder_CH3data_0));
    LocalMux I__2209 (
            .O(N__13450),
            .I(frame_decoder_CH3data_0));
    InMux I__2208 (
            .O(N__13443),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__2207 (
            .O(N__13440),
            .I(\ppm_encoder_1.un1_aileron_cry_7 ));
    InMux I__2206 (
            .O(N__13437),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__2205 (
            .O(N__13434),
            .I(N__13431));
    LocalMux I__2204 (
            .O(N__13431),
            .I(N__13427));
    InMux I__2203 (
            .O(N__13430),
            .I(N__13424));
    Span4Mux_h I__2202 (
            .O(N__13427),
            .I(N__13421));
    LocalMux I__2201 (
            .O(N__13424),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    Odrv4 I__2200 (
            .O(N__13421),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    InMux I__2199 (
            .O(N__13416),
            .I(N__13413));
    LocalMux I__2198 (
            .O(N__13413),
            .I(N__13410));
    Span4Mux_h I__2197 (
            .O(N__13410),
            .I(N__13407));
    Odrv4 I__2196 (
            .O(N__13407),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa ));
    CascadeMux I__2195 (
            .O(N__13404),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_ ));
    CEMux I__2194 (
            .O(N__13401),
            .I(N__13398));
    LocalMux I__2193 (
            .O(N__13398),
            .I(N__13395));
    Span4Mux_h I__2192 (
            .O(N__13395),
            .I(N__13392));
    Span4Mux_v I__2191 (
            .O(N__13392),
            .I(N__13389));
    Odrv4 I__2190 (
            .O(N__13389),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa_0 ));
    InMux I__2189 (
            .O(N__13386),
            .I(N__13368));
    InMux I__2188 (
            .O(N__13385),
            .I(N__13368));
    InMux I__2187 (
            .O(N__13384),
            .I(N__13368));
    InMux I__2186 (
            .O(N__13383),
            .I(N__13368));
    InMux I__2185 (
            .O(N__13382),
            .I(N__13368));
    InMux I__2184 (
            .O(N__13381),
            .I(N__13361));
    InMux I__2183 (
            .O(N__13380),
            .I(N__13361));
    InMux I__2182 (
            .O(N__13379),
            .I(N__13361));
    LocalMux I__2181 (
            .O(N__13368),
            .I(N__13355));
    LocalMux I__2180 (
            .O(N__13361),
            .I(N__13355));
    InMux I__2179 (
            .O(N__13360),
            .I(N__13352));
    Odrv4 I__2178 (
            .O(N__13355),
            .I(\uart.data_rdyc_1 ));
    LocalMux I__2177 (
            .O(N__13352),
            .I(\uart.data_rdyc_1 ));
    InMux I__2176 (
            .O(N__13347),
            .I(N__13343));
    CascadeMux I__2175 (
            .O(N__13346),
            .I(N__13340));
    LocalMux I__2174 (
            .O(N__13343),
            .I(N__13337));
    InMux I__2173 (
            .O(N__13340),
            .I(N__13334));
    Odrv4 I__2172 (
            .O(N__13337),
            .I(\uart.data_AuxZ0Z_4 ));
    LocalMux I__2171 (
            .O(N__13334),
            .I(\uart.data_AuxZ0Z_4 ));
    SRMux I__2170 (
            .O(N__13329),
            .I(N__13326));
    LocalMux I__2169 (
            .O(N__13326),
            .I(N__13322));
    SRMux I__2168 (
            .O(N__13325),
            .I(N__13319));
    Span4Mux_h I__2167 (
            .O(N__13322),
            .I(N__13316));
    LocalMux I__2166 (
            .O(N__13319),
            .I(N__13313));
    Odrv4 I__2165 (
            .O(N__13316),
            .I(\uart.state_RNIQABT2Z0Z_4 ));
    Odrv12 I__2164 (
            .O(N__13313),
            .I(\uart.state_RNIQABT2Z0Z_4 ));
    InMux I__2163 (
            .O(N__13308),
            .I(N__13305));
    LocalMux I__2162 (
            .O(N__13305),
            .I(N__13302));
    Span4Mux_h I__2161 (
            .O(N__13302),
            .I(N__13298));
    InMux I__2160 (
            .O(N__13301),
            .I(N__13295));
    Odrv4 I__2159 (
            .O(N__13298),
            .I(\uart_frame_decoder.state_1_ns_0_i_o2_0_10 ));
    LocalMux I__2158 (
            .O(N__13295),
            .I(\uart_frame_decoder.state_1_ns_0_i_o2_0_10 ));
    CascadeMux I__2157 (
            .O(N__13290),
            .I(N__13286));
    InMux I__2156 (
            .O(N__13289),
            .I(N__13283));
    InMux I__2155 (
            .O(N__13286),
            .I(N__13280));
    LocalMux I__2154 (
            .O(N__13283),
            .I(N__13277));
    LocalMux I__2153 (
            .O(N__13280),
            .I(N__13274));
    Span4Mux_v I__2152 (
            .O(N__13277),
            .I(N__13271));
    Odrv4 I__2151 (
            .O(N__13274),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa ));
    Odrv4 I__2150 (
            .O(N__13271),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa ));
    InMux I__2149 (
            .O(N__13266),
            .I(N__13254));
    InMux I__2148 (
            .O(N__13265),
            .I(N__13254));
    InMux I__2147 (
            .O(N__13264),
            .I(N__13254));
    InMux I__2146 (
            .O(N__13263),
            .I(N__13254));
    LocalMux I__2145 (
            .O(N__13254),
            .I(N__13250));
    InMux I__2144 (
            .O(N__13253),
            .I(N__13247));
    Span4Mux_v I__2143 (
            .O(N__13250),
            .I(N__13241));
    LocalMux I__2142 (
            .O(N__13247),
            .I(N__13241));
    InMux I__2141 (
            .O(N__13246),
            .I(N__13238));
    Span4Mux_v I__2140 (
            .O(N__13241),
            .I(N__13231));
    LocalMux I__2139 (
            .O(N__13238),
            .I(N__13228));
    InMux I__2138 (
            .O(N__13237),
            .I(N__13225));
    InMux I__2137 (
            .O(N__13236),
            .I(N__13218));
    InMux I__2136 (
            .O(N__13235),
            .I(N__13218));
    InMux I__2135 (
            .O(N__13234),
            .I(N__13218));
    Odrv4 I__2134 (
            .O(N__13231),
            .I(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ));
    Odrv4 I__2133 (
            .O(N__13228),
            .I(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ));
    LocalMux I__2132 (
            .O(N__13225),
            .I(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ));
    LocalMux I__2131 (
            .O(N__13218),
            .I(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ));
    InMux I__2130 (
            .O(N__13209),
            .I(N__13205));
    InMux I__2129 (
            .O(N__13208),
            .I(N__13202));
    LocalMux I__2128 (
            .O(N__13205),
            .I(N__13199));
    LocalMux I__2127 (
            .O(N__13202),
            .I(N__13196));
    Span12Mux_v I__2126 (
            .O(N__13199),
            .I(N__13193));
    Span4Mux_h I__2125 (
            .O(N__13196),
            .I(N__13190));
    Odrv12 I__2124 (
            .O(N__13193),
            .I(scaler_4_data_11));
    Odrv4 I__2123 (
            .O(N__13190),
            .I(scaler_4_data_11));
    InMux I__2122 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__2121 (
            .O(N__13182),
            .I(N__13179));
    Span4Mux_v I__2120 (
            .O(N__13179),
            .I(N__13176));
    Odrv4 I__2119 (
            .O(N__13176),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    CascadeMux I__2118 (
            .O(N__13173),
            .I(N__13169));
    InMux I__2117 (
            .O(N__13172),
            .I(N__13165));
    InMux I__2116 (
            .O(N__13169),
            .I(N__13162));
    CascadeMux I__2115 (
            .O(N__13168),
            .I(N__13158));
    LocalMux I__2114 (
            .O(N__13165),
            .I(N__13149));
    LocalMux I__2113 (
            .O(N__13162),
            .I(N__13149));
    InMux I__2112 (
            .O(N__13161),
            .I(N__13140));
    InMux I__2111 (
            .O(N__13158),
            .I(N__13140));
    InMux I__2110 (
            .O(N__13157),
            .I(N__13140));
    InMux I__2109 (
            .O(N__13156),
            .I(N__13140));
    InMux I__2108 (
            .O(N__13155),
            .I(N__13137));
    InMux I__2107 (
            .O(N__13154),
            .I(N__13134));
    Span4Mux_v I__2106 (
            .O(N__13149),
            .I(N__13131));
    LocalMux I__2105 (
            .O(N__13140),
            .I(N__13128));
    LocalMux I__2104 (
            .O(N__13137),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__2103 (
            .O(N__13134),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    Odrv4 I__2102 (
            .O(N__13131),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    Odrv4 I__2101 (
            .O(N__13128),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    CascadeMux I__2100 (
            .O(N__13119),
            .I(N__13113));
    InMux I__2099 (
            .O(N__13118),
            .I(N__13107));
    InMux I__2098 (
            .O(N__13117),
            .I(N__13103));
    InMux I__2097 (
            .O(N__13116),
            .I(N__13100));
    InMux I__2096 (
            .O(N__13113),
            .I(N__13094));
    InMux I__2095 (
            .O(N__13112),
            .I(N__13094));
    InMux I__2094 (
            .O(N__13111),
            .I(N__13084));
    InMux I__2093 (
            .O(N__13110),
            .I(N__13084));
    LocalMux I__2092 (
            .O(N__13107),
            .I(N__13081));
    InMux I__2091 (
            .O(N__13106),
            .I(N__13078));
    LocalMux I__2090 (
            .O(N__13103),
            .I(N__13075));
    LocalMux I__2089 (
            .O(N__13100),
            .I(N__13072));
    InMux I__2088 (
            .O(N__13099),
            .I(N__13069));
    LocalMux I__2087 (
            .O(N__13094),
            .I(N__13066));
    InMux I__2086 (
            .O(N__13093),
            .I(N__13063));
    InMux I__2085 (
            .O(N__13092),
            .I(N__13054));
    InMux I__2084 (
            .O(N__13091),
            .I(N__13054));
    InMux I__2083 (
            .O(N__13090),
            .I(N__13054));
    InMux I__2082 (
            .O(N__13089),
            .I(N__13051));
    LocalMux I__2081 (
            .O(N__13084),
            .I(N__13044));
    Span4Mux_s3_h I__2080 (
            .O(N__13081),
            .I(N__13044));
    LocalMux I__2079 (
            .O(N__13078),
            .I(N__13044));
    Span4Mux_v I__2078 (
            .O(N__13075),
            .I(N__13039));
    Span4Mux_v I__2077 (
            .O(N__13072),
            .I(N__13039));
    LocalMux I__2076 (
            .O(N__13069),
            .I(N__13032));
    Span4Mux_h I__2075 (
            .O(N__13066),
            .I(N__13032));
    LocalMux I__2074 (
            .O(N__13063),
            .I(N__13032));
    InMux I__2073 (
            .O(N__13062),
            .I(N__13027));
    InMux I__2072 (
            .O(N__13061),
            .I(N__13027));
    LocalMux I__2071 (
            .O(N__13054),
            .I(N__13020));
    LocalMux I__2070 (
            .O(N__13051),
            .I(N__13020));
    Span4Mux_v I__2069 (
            .O(N__13044),
            .I(N__13020));
    Odrv4 I__2068 (
            .O(N__13039),
            .I(uart_data_rdy));
    Odrv4 I__2067 (
            .O(N__13032),
            .I(uart_data_rdy));
    LocalMux I__2066 (
            .O(N__13027),
            .I(uart_data_rdy));
    Odrv4 I__2065 (
            .O(N__13020),
            .I(uart_data_rdy));
    InMux I__2064 (
            .O(N__13011),
            .I(N__13008));
    LocalMux I__2063 (
            .O(N__13008),
            .I(N__13005));
    Span4Mux_v I__2062 (
            .O(N__13005),
            .I(N__13001));
    InMux I__2061 (
            .O(N__13004),
            .I(N__12998));
    Odrv4 I__2060 (
            .O(N__13001),
            .I(\uart_frame_decoder.count8_THRU_CO ));
    LocalMux I__2059 (
            .O(N__12998),
            .I(\uart_frame_decoder.count8_THRU_CO ));
    InMux I__2058 (
            .O(N__12993),
            .I(N__12987));
    InMux I__2057 (
            .O(N__12992),
            .I(N__12987));
    LocalMux I__2056 (
            .O(N__12987),
            .I(N__12982));
    CascadeMux I__2055 (
            .O(N__12986),
            .I(N__12978));
    InMux I__2054 (
            .O(N__12985),
            .I(N__12970));
    Span4Mux_h I__2053 (
            .O(N__12982),
            .I(N__12967));
    InMux I__2052 (
            .O(N__12981),
            .I(N__12964));
    InMux I__2051 (
            .O(N__12978),
            .I(N__12961));
    InMux I__2050 (
            .O(N__12977),
            .I(N__12950));
    InMux I__2049 (
            .O(N__12976),
            .I(N__12950));
    InMux I__2048 (
            .O(N__12975),
            .I(N__12950));
    InMux I__2047 (
            .O(N__12974),
            .I(N__12950));
    InMux I__2046 (
            .O(N__12973),
            .I(N__12950));
    LocalMux I__2045 (
            .O(N__12970),
            .I(\uart.bit_CountZ0Z_2 ));
    Odrv4 I__2044 (
            .O(N__12967),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__2043 (
            .O(N__12964),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__2042 (
            .O(N__12961),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__2041 (
            .O(N__12950),
            .I(\uart.bit_CountZ0Z_2 ));
    CascadeMux I__2040 (
            .O(N__12939),
            .I(N__12936));
    InMux I__2039 (
            .O(N__12936),
            .I(N__12930));
    InMux I__2038 (
            .O(N__12935),
            .I(N__12930));
    LocalMux I__2037 (
            .O(N__12930),
            .I(N__12926));
    InMux I__2036 (
            .O(N__12929),
            .I(N__12915));
    Span4Mux_h I__2035 (
            .O(N__12926),
            .I(N__12912));
    InMux I__2034 (
            .O(N__12925),
            .I(N__12907));
    InMux I__2033 (
            .O(N__12924),
            .I(N__12907));
    InMux I__2032 (
            .O(N__12923),
            .I(N__12904));
    InMux I__2031 (
            .O(N__12922),
            .I(N__12899));
    InMux I__2030 (
            .O(N__12921),
            .I(N__12899));
    InMux I__2029 (
            .O(N__12920),
            .I(N__12892));
    InMux I__2028 (
            .O(N__12919),
            .I(N__12892));
    InMux I__2027 (
            .O(N__12918),
            .I(N__12892));
    LocalMux I__2026 (
            .O(N__12915),
            .I(\uart.bit_CountZ0Z_1 ));
    Odrv4 I__2025 (
            .O(N__12912),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__2024 (
            .O(N__12907),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__2023 (
            .O(N__12904),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__2022 (
            .O(N__12899),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__2021 (
            .O(N__12892),
            .I(\uart.bit_CountZ0Z_1 ));
    InMux I__2020 (
            .O(N__12879),
            .I(N__12871));
    InMux I__2019 (
            .O(N__12878),
            .I(N__12871));
    InMux I__2018 (
            .O(N__12877),
            .I(N__12866));
    InMux I__2017 (
            .O(N__12876),
            .I(N__12866));
    LocalMux I__2016 (
            .O(N__12871),
            .I(N__12863));
    LocalMux I__2015 (
            .O(N__12866),
            .I(N__12850));
    Span4Mux_v I__2014 (
            .O(N__12863),
            .I(N__12850));
    InMux I__2013 (
            .O(N__12862),
            .I(N__12847));
    InMux I__2012 (
            .O(N__12861),
            .I(N__12842));
    InMux I__2011 (
            .O(N__12860),
            .I(N__12842));
    InMux I__2010 (
            .O(N__12859),
            .I(N__12831));
    InMux I__2009 (
            .O(N__12858),
            .I(N__12831));
    InMux I__2008 (
            .O(N__12857),
            .I(N__12831));
    InMux I__2007 (
            .O(N__12856),
            .I(N__12831));
    InMux I__2006 (
            .O(N__12855),
            .I(N__12831));
    Odrv4 I__2005 (
            .O(N__12850),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__2004 (
            .O(N__12847),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__2003 (
            .O(N__12842),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__2002 (
            .O(N__12831),
            .I(\uart.bit_CountZ0Z_0 ));
    InMux I__2001 (
            .O(N__12822),
            .I(N__12819));
    LocalMux I__2000 (
            .O(N__12819),
            .I(\uart.data_Auxce_0_0_2 ));
    InMux I__1999 (
            .O(N__12816),
            .I(N__12813));
    LocalMux I__1998 (
            .O(N__12813),
            .I(N__12810));
    Odrv4 I__1997 (
            .O(N__12810),
            .I(\reset_module_System.reset6_13 ));
    InMux I__1996 (
            .O(N__12807),
            .I(N__12804));
    LocalMux I__1995 (
            .O(N__12804),
            .I(\reset_module_System.reset6_3 ));
    InMux I__1994 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__1993 (
            .O(N__12798),
            .I(N__12795));
    Odrv4 I__1992 (
            .O(N__12795),
            .I(\reset_module_System.reset6_17 ));
    InMux I__1991 (
            .O(N__12792),
            .I(N__12789));
    LocalMux I__1990 (
            .O(N__12789),
            .I(N__12783));
    InMux I__1989 (
            .O(N__12788),
            .I(N__12780));
    InMux I__1988 (
            .O(N__12787),
            .I(N__12774));
    InMux I__1987 (
            .O(N__12786),
            .I(N__12771));
    Span4Mux_s1_v I__1986 (
            .O(N__12783),
            .I(N__12766));
    LocalMux I__1985 (
            .O(N__12780),
            .I(N__12766));
    InMux I__1984 (
            .O(N__12779),
            .I(N__12763));
    InMux I__1983 (
            .O(N__12778),
            .I(N__12760));
    InMux I__1982 (
            .O(N__12777),
            .I(N__12757));
    LocalMux I__1981 (
            .O(N__12774),
            .I(N__12752));
    LocalMux I__1980 (
            .O(N__12771),
            .I(N__12752));
    Span4Mux_v I__1979 (
            .O(N__12766),
            .I(N__12745));
    LocalMux I__1978 (
            .O(N__12763),
            .I(N__12745));
    LocalMux I__1977 (
            .O(N__12760),
            .I(N__12745));
    LocalMux I__1976 (
            .O(N__12757),
            .I(N__12742));
    Span12Mux_s10_v I__1975 (
            .O(N__12752),
            .I(N__12736));
    Span4Mux_v I__1974 (
            .O(N__12745),
            .I(N__12731));
    Span4Mux_s3_h I__1973 (
            .O(N__12742),
            .I(N__12731));
    InMux I__1972 (
            .O(N__12741),
            .I(N__12728));
    InMux I__1971 (
            .O(N__12740),
            .I(N__12725));
    InMux I__1970 (
            .O(N__12739),
            .I(N__12722));
    Odrv12 I__1969 (
            .O(N__12736),
            .I(uart_data_1));
    Odrv4 I__1968 (
            .O(N__12731),
            .I(uart_data_1));
    LocalMux I__1967 (
            .O(N__12728),
            .I(uart_data_1));
    LocalMux I__1966 (
            .O(N__12725),
            .I(uart_data_1));
    LocalMux I__1965 (
            .O(N__12722),
            .I(uart_data_1));
    CascadeMux I__1964 (
            .O(N__12711),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ));
    CascadeMux I__1963 (
            .O(N__12708),
            .I(N__12705));
    InMux I__1962 (
            .O(N__12705),
            .I(N__12699));
    InMux I__1961 (
            .O(N__12704),
            .I(N__12699));
    LocalMux I__1960 (
            .O(N__12699),
            .I(N__12695));
    InMux I__1959 (
            .O(N__12698),
            .I(N__12692));
    Span4Mux_h I__1958 (
            .O(N__12695),
            .I(N__12689));
    LocalMux I__1957 (
            .O(N__12692),
            .I(N__12686));
    Odrv4 I__1956 (
            .O(N__12689),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ));
    Odrv4 I__1955 (
            .O(N__12686),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ));
    InMux I__1954 (
            .O(N__12681),
            .I(N__12677));
    InMux I__1953 (
            .O(N__12680),
            .I(N__12674));
    LocalMux I__1952 (
            .O(N__12677),
            .I(N__12671));
    LocalMux I__1951 (
            .O(N__12674),
            .I(\uart.stateZ0Z_0 ));
    Odrv4 I__1950 (
            .O(N__12671),
            .I(\uart.stateZ0Z_0 ));
    CascadeMux I__1949 (
            .O(N__12666),
            .I(N__12663));
    InMux I__1948 (
            .O(N__12663),
            .I(N__12660));
    LocalMux I__1947 (
            .O(N__12660),
            .I(N__12655));
    InMux I__1946 (
            .O(N__12659),
            .I(N__12652));
    InMux I__1945 (
            .O(N__12658),
            .I(N__12649));
    Sp12to4 I__1944 (
            .O(N__12655),
            .I(N__12644));
    LocalMux I__1943 (
            .O(N__12652),
            .I(N__12644));
    LocalMux I__1942 (
            .O(N__12649),
            .I(\uart.stateZ0Z_1 ));
    Odrv12 I__1941 (
            .O(N__12644),
            .I(\uart.stateZ0Z_1 ));
    CascadeMux I__1940 (
            .O(N__12639),
            .I(N__12634));
    CascadeMux I__1939 (
            .O(N__12638),
            .I(N__12623));
    CascadeMux I__1938 (
            .O(N__12637),
            .I(N__12620));
    InMux I__1937 (
            .O(N__12634),
            .I(N__12603));
    InMux I__1936 (
            .O(N__12633),
            .I(N__12603));
    InMux I__1935 (
            .O(N__12632),
            .I(N__12603));
    InMux I__1934 (
            .O(N__12631),
            .I(N__12603));
    InMux I__1933 (
            .O(N__12630),
            .I(N__12603));
    InMux I__1932 (
            .O(N__12629),
            .I(N__12603));
    InMux I__1931 (
            .O(N__12628),
            .I(N__12603));
    InMux I__1930 (
            .O(N__12627),
            .I(N__12603));
    InMux I__1929 (
            .O(N__12626),
            .I(N__12600));
    InMux I__1928 (
            .O(N__12623),
            .I(N__12596));
    InMux I__1927 (
            .O(N__12620),
            .I(N__12592));
    LocalMux I__1926 (
            .O(N__12603),
            .I(N__12587));
    LocalMux I__1925 (
            .O(N__12600),
            .I(N__12587));
    InMux I__1924 (
            .O(N__12599),
            .I(N__12584));
    LocalMux I__1923 (
            .O(N__12596),
            .I(N__12581));
    InMux I__1922 (
            .O(N__12595),
            .I(N__12578));
    LocalMux I__1921 (
            .O(N__12592),
            .I(N__12571));
    Sp12to4 I__1920 (
            .O(N__12587),
            .I(N__12571));
    LocalMux I__1919 (
            .O(N__12584),
            .I(N__12571));
    Odrv4 I__1918 (
            .O(N__12581),
            .I(uart_input_sync));
    LocalMux I__1917 (
            .O(N__12578),
            .I(uart_input_sync));
    Odrv12 I__1916 (
            .O(N__12571),
            .I(uart_input_sync));
    InMux I__1915 (
            .O(N__12564),
            .I(N__12560));
    CascadeMux I__1914 (
            .O(N__12563),
            .I(N__12557));
    LocalMux I__1913 (
            .O(N__12560),
            .I(N__12554));
    InMux I__1912 (
            .O(N__12557),
            .I(N__12551));
    Odrv4 I__1911 (
            .O(N__12554),
            .I(\uart.data_AuxZ0Z_3 ));
    LocalMux I__1910 (
            .O(N__12551),
            .I(\uart.data_AuxZ0Z_3 ));
    InMux I__1909 (
            .O(N__12546),
            .I(N__12540));
    InMux I__1908 (
            .O(N__12545),
            .I(N__12537));
    InMux I__1907 (
            .O(N__12544),
            .I(N__12534));
    InMux I__1906 (
            .O(N__12543),
            .I(N__12531));
    LocalMux I__1905 (
            .O(N__12540),
            .I(N__12519));
    LocalMux I__1904 (
            .O(N__12537),
            .I(N__12519));
    LocalMux I__1903 (
            .O(N__12534),
            .I(N__12519));
    LocalMux I__1902 (
            .O(N__12531),
            .I(N__12519));
    InMux I__1901 (
            .O(N__12530),
            .I(N__12516));
    InMux I__1900 (
            .O(N__12529),
            .I(N__12513));
    InMux I__1899 (
            .O(N__12528),
            .I(N__12510));
    Span4Mux_v I__1898 (
            .O(N__12519),
            .I(N__12500));
    LocalMux I__1897 (
            .O(N__12516),
            .I(N__12500));
    LocalMux I__1896 (
            .O(N__12513),
            .I(N__12500));
    LocalMux I__1895 (
            .O(N__12510),
            .I(N__12500));
    InMux I__1894 (
            .O(N__12509),
            .I(N__12497));
    Span4Mux_v I__1893 (
            .O(N__12500),
            .I(N__12490));
    LocalMux I__1892 (
            .O(N__12497),
            .I(N__12490));
    InMux I__1891 (
            .O(N__12496),
            .I(N__12487));
    InMux I__1890 (
            .O(N__12495),
            .I(N__12484));
    Odrv4 I__1889 (
            .O(N__12490),
            .I(uart_data_3));
    LocalMux I__1888 (
            .O(N__12487),
            .I(uart_data_3));
    LocalMux I__1887 (
            .O(N__12484),
            .I(uart_data_3));
    InMux I__1886 (
            .O(N__12477),
            .I(N__12474));
    LocalMux I__1885 (
            .O(N__12474),
            .I(N__12471));
    Span4Mux_v I__1884 (
            .O(N__12471),
            .I(N__12467));
    InMux I__1883 (
            .O(N__12470),
            .I(N__12464));
    Odrv4 I__1882 (
            .O(N__12467),
            .I(\uart.data_AuxZ0Z_6 ));
    LocalMux I__1881 (
            .O(N__12464),
            .I(\uart.data_AuxZ0Z_6 ));
    InMux I__1880 (
            .O(N__12459),
            .I(N__12452));
    InMux I__1879 (
            .O(N__12458),
            .I(N__12449));
    InMux I__1878 (
            .O(N__12457),
            .I(N__12446));
    InMux I__1877 (
            .O(N__12456),
            .I(N__12443));
    InMux I__1876 (
            .O(N__12455),
            .I(N__12440));
    LocalMux I__1875 (
            .O(N__12452),
            .I(N__12435));
    LocalMux I__1874 (
            .O(N__12449),
            .I(N__12432));
    LocalMux I__1873 (
            .O(N__12446),
            .I(N__12427));
    LocalMux I__1872 (
            .O(N__12443),
            .I(N__12427));
    LocalMux I__1871 (
            .O(N__12440),
            .I(N__12424));
    InMux I__1870 (
            .O(N__12439),
            .I(N__12421));
    InMux I__1869 (
            .O(N__12438),
            .I(N__12418));
    Span4Mux_v I__1868 (
            .O(N__12435),
            .I(N__12414));
    Span4Mux_h I__1867 (
            .O(N__12432),
            .I(N__12411));
    Span4Mux_v I__1866 (
            .O(N__12427),
            .I(N__12402));
    Span4Mux_h I__1865 (
            .O(N__12424),
            .I(N__12402));
    LocalMux I__1864 (
            .O(N__12421),
            .I(N__12402));
    LocalMux I__1863 (
            .O(N__12418),
            .I(N__12402));
    InMux I__1862 (
            .O(N__12417),
            .I(N__12399));
    Span4Mux_v I__1861 (
            .O(N__12414),
            .I(N__12394));
    Span4Mux_v I__1860 (
            .O(N__12411),
            .I(N__12391));
    Span4Mux_v I__1859 (
            .O(N__12402),
            .I(N__12386));
    LocalMux I__1858 (
            .O(N__12399),
            .I(N__12386));
    InMux I__1857 (
            .O(N__12398),
            .I(N__12383));
    InMux I__1856 (
            .O(N__12397),
            .I(N__12380));
    Odrv4 I__1855 (
            .O(N__12394),
            .I(uart_data_6));
    Odrv4 I__1854 (
            .O(N__12391),
            .I(uart_data_6));
    Odrv4 I__1853 (
            .O(N__12386),
            .I(uart_data_6));
    LocalMux I__1852 (
            .O(N__12383),
            .I(uart_data_6));
    LocalMux I__1851 (
            .O(N__12380),
            .I(uart_data_6));
    CascadeMux I__1850 (
            .O(N__12369),
            .I(\reset_module_System.reset6_11_cascade_ ));
    InMux I__1849 (
            .O(N__12366),
            .I(N__12361));
    InMux I__1848 (
            .O(N__12365),
            .I(N__12356));
    InMux I__1847 (
            .O(N__12364),
            .I(N__12356));
    LocalMux I__1846 (
            .O(N__12361),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__1845 (
            .O(N__12356),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__1844 (
            .O(N__12351),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__1843 (
            .O(N__12348),
            .I(N__12345));
    LocalMux I__1842 (
            .O(N__12345),
            .I(\uart.data_Auxce_0_0_4 ));
    InMux I__1841 (
            .O(N__12342),
            .I(N__12334));
    InMux I__1840 (
            .O(N__12341),
            .I(N__12334));
    InMux I__1839 (
            .O(N__12340),
            .I(N__12329));
    InMux I__1838 (
            .O(N__12339),
            .I(N__12329));
    LocalMux I__1837 (
            .O(N__12334),
            .I(N__12326));
    LocalMux I__1836 (
            .O(N__12329),
            .I(\reset_module_System.reset6_14 ));
    Odrv4 I__1835 (
            .O(N__12326),
            .I(\reset_module_System.reset6_14 ));
    SRMux I__1834 (
            .O(N__12321),
            .I(N__12318));
    LocalMux I__1833 (
            .O(N__12318),
            .I(N__12315));
    Odrv12 I__1832 (
            .O(N__12315),
            .I(\uart.state_RNIAFHLZ0Z_3 ));
    InMux I__1831 (
            .O(N__12312),
            .I(N__12306));
    InMux I__1830 (
            .O(N__12311),
            .I(N__12303));
    InMux I__1829 (
            .O(N__12310),
            .I(N__12300));
    InMux I__1828 (
            .O(N__12309),
            .I(N__12297));
    LocalMux I__1827 (
            .O(N__12306),
            .I(N__12292));
    LocalMux I__1826 (
            .O(N__12303),
            .I(N__12292));
    LocalMux I__1825 (
            .O(N__12300),
            .I(\uart.N_153_0 ));
    LocalMux I__1824 (
            .O(N__12297),
            .I(\uart.N_153_0 ));
    Odrv4 I__1823 (
            .O(N__12292),
            .I(\uart.N_153_0 ));
    InMux I__1822 (
            .O(N__12285),
            .I(N__12281));
    InMux I__1821 (
            .O(N__12284),
            .I(N__12278));
    LocalMux I__1820 (
            .O(N__12281),
            .I(N__12267));
    LocalMux I__1819 (
            .O(N__12278),
            .I(N__12267));
    InMux I__1818 (
            .O(N__12277),
            .I(N__12264));
    InMux I__1817 (
            .O(N__12276),
            .I(N__12261));
    InMux I__1816 (
            .O(N__12275),
            .I(N__12258));
    InMux I__1815 (
            .O(N__12274),
            .I(N__12255));
    InMux I__1814 (
            .O(N__12273),
            .I(N__12250));
    InMux I__1813 (
            .O(N__12272),
            .I(N__12250));
    Odrv4 I__1812 (
            .O(N__12267),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__1811 (
            .O(N__12264),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__1810 (
            .O(N__12261),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__1809 (
            .O(N__12258),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__1808 (
            .O(N__12255),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__1807 (
            .O(N__12250),
            .I(\uart.stateZ0Z_3 ));
    CascadeMux I__1806 (
            .O(N__12237),
            .I(N__12234));
    InMux I__1805 (
            .O(N__12234),
            .I(N__12231));
    LocalMux I__1804 (
            .O(N__12231),
            .I(N__12228));
    Odrv4 I__1803 (
            .O(N__12228),
            .I(\uart.N_168_1 ));
    InMux I__1802 (
            .O(N__12225),
            .I(N__12222));
    LocalMux I__1801 (
            .O(N__12222),
            .I(N__12219));
    Odrv4 I__1800 (
            .O(N__12219),
            .I(\uart.N_167 ));
    CascadeMux I__1799 (
            .O(N__12216),
            .I(N__12210));
    CascadeMux I__1798 (
            .O(N__12215),
            .I(N__12203));
    InMux I__1797 (
            .O(N__12214),
            .I(N__12197));
    InMux I__1796 (
            .O(N__12213),
            .I(N__12197));
    InMux I__1795 (
            .O(N__12210),
            .I(N__12192));
    InMux I__1794 (
            .O(N__12209),
            .I(N__12192));
    InMux I__1793 (
            .O(N__12208),
            .I(N__12189));
    InMux I__1792 (
            .O(N__12207),
            .I(N__12186));
    InMux I__1791 (
            .O(N__12206),
            .I(N__12183));
    InMux I__1790 (
            .O(N__12203),
            .I(N__12180));
    InMux I__1789 (
            .O(N__12202),
            .I(N__12177));
    LocalMux I__1788 (
            .O(N__12197),
            .I(N__12174));
    LocalMux I__1787 (
            .O(N__12192),
            .I(N__12171));
    LocalMux I__1786 (
            .O(N__12189),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1785 (
            .O(N__12186),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1784 (
            .O(N__12183),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1783 (
            .O(N__12180),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__1782 (
            .O(N__12177),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__1781 (
            .O(N__12174),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__1780 (
            .O(N__12171),
            .I(\uart.stateZ0Z_4 ));
    CascadeMux I__1779 (
            .O(N__12156),
            .I(\reset_module_System.count_1_1_cascade_ ));
    CascadeMux I__1778 (
            .O(N__12153),
            .I(\uart.N_153_0_cascade_ ));
    CascadeMux I__1777 (
            .O(N__12150),
            .I(\uart.state_srsts_i_a3_0_0_3_cascade_ ));
    InMux I__1776 (
            .O(N__12147),
            .I(N__12144));
    LocalMux I__1775 (
            .O(N__12144),
            .I(\uart.N_170 ));
    InMux I__1774 (
            .O(N__12141),
            .I(N__12138));
    LocalMux I__1773 (
            .O(N__12138),
            .I(\uart.un1_state_2_0_a3_2 ));
    InMux I__1772 (
            .O(N__12135),
            .I(N__12132));
    LocalMux I__1771 (
            .O(N__12132),
            .I(N__12128));
    InMux I__1770 (
            .O(N__12131),
            .I(N__12125));
    Odrv4 I__1769 (
            .O(N__12128),
            .I(\uart.N_146_0 ));
    LocalMux I__1768 (
            .O(N__12125),
            .I(\uart.N_146_0 ));
    InMux I__1767 (
            .O(N__12120),
            .I(N__12096));
    InMux I__1766 (
            .O(N__12119),
            .I(N__12096));
    InMux I__1765 (
            .O(N__12118),
            .I(N__12096));
    InMux I__1764 (
            .O(N__12117),
            .I(N__12096));
    InMux I__1763 (
            .O(N__12116),
            .I(N__12096));
    InMux I__1762 (
            .O(N__12115),
            .I(N__12096));
    InMux I__1761 (
            .O(N__12114),
            .I(N__12096));
    InMux I__1760 (
            .O(N__12113),
            .I(N__12096));
    LocalMux I__1759 (
            .O(N__12096),
            .I(\uart.un1_state_2_0 ));
    InMux I__1758 (
            .O(N__12093),
            .I(N__12090));
    LocalMux I__1757 (
            .O(N__12090),
            .I(\uart.N_151 ));
    InMux I__1756 (
            .O(N__12087),
            .I(N__12081));
    InMux I__1755 (
            .O(N__12086),
            .I(N__12078));
    InMux I__1754 (
            .O(N__12085),
            .I(N__12075));
    InMux I__1753 (
            .O(N__12084),
            .I(N__12072));
    LocalMux I__1752 (
            .O(N__12081),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__1751 (
            .O(N__12078),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__1750 (
            .O(N__12075),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__1749 (
            .O(N__12072),
            .I(\uart.stateZ0Z_2 ));
    InMux I__1748 (
            .O(N__12063),
            .I(N__12060));
    LocalMux I__1747 (
            .O(N__12060),
            .I(\uart.N_159 ));
    CascadeMux I__1746 (
            .O(N__12057),
            .I(\uart.timer_Count_0_sqmuxa_1_cascade_ ));
    InMux I__1745 (
            .O(N__12054),
            .I(N__12048));
    InMux I__1744 (
            .O(N__12053),
            .I(N__12048));
    LocalMux I__1743 (
            .O(N__12048),
            .I(\uart.N_180 ));
    CascadeMux I__1742 (
            .O(N__12045),
            .I(\uart.N_180_cascade_ ));
    InMux I__1741 (
            .O(N__12042),
            .I(N__12033));
    InMux I__1740 (
            .O(N__12041),
            .I(N__12033));
    InMux I__1739 (
            .O(N__12040),
            .I(N__12033));
    LocalMux I__1738 (
            .O(N__12033),
            .I(N__12029));
    InMux I__1737 (
            .O(N__12032),
            .I(N__12026));
    Odrv4 I__1736 (
            .O(N__12029),
            .I(\uart.un1_state_5_0 ));
    LocalMux I__1735 (
            .O(N__12026),
            .I(\uart.un1_state_5_0 ));
    InMux I__1734 (
            .O(N__12021),
            .I(N__12017));
    InMux I__1733 (
            .O(N__12020),
            .I(N__12014));
    LocalMux I__1732 (
            .O(N__12017),
            .I(\uart.N_143_0 ));
    LocalMux I__1731 (
            .O(N__12014),
            .I(\uart.N_143_0 ));
    CascadeMux I__1730 (
            .O(N__12009),
            .I(N__12006));
    InMux I__1729 (
            .O(N__12006),
            .I(N__12000));
    InMux I__1728 (
            .O(N__12005),
            .I(N__12000));
    LocalMux I__1727 (
            .O(N__12000),
            .I(\scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ));
    InMux I__1726 (
            .O(N__11997),
            .I(\scaler_1.un2_source_data_0_cry_7 ));
    InMux I__1725 (
            .O(N__11994),
            .I(N__11990));
    InMux I__1724 (
            .O(N__11993),
            .I(N__11987));
    LocalMux I__1723 (
            .O(N__11990),
            .I(\scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ));
    LocalMux I__1722 (
            .O(N__11987),
            .I(\scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ));
    CascadeMux I__1721 (
            .O(N__11982),
            .I(N__11979));
    InMux I__1720 (
            .O(N__11979),
            .I(N__11976));
    LocalMux I__1719 (
            .O(N__11976),
            .I(\scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ));
    InMux I__1718 (
            .O(N__11973),
            .I(bfn_3_29_0_));
    InMux I__1717 (
            .O(N__11970),
            .I(\scaler_1.un2_source_data_0_cry_9 ));
    CEMux I__1716 (
            .O(N__11967),
            .I(N__11940));
    CEMux I__1715 (
            .O(N__11966),
            .I(N__11940));
    CEMux I__1714 (
            .O(N__11965),
            .I(N__11940));
    CEMux I__1713 (
            .O(N__11964),
            .I(N__11940));
    CEMux I__1712 (
            .O(N__11963),
            .I(N__11940));
    CEMux I__1711 (
            .O(N__11962),
            .I(N__11940));
    CEMux I__1710 (
            .O(N__11961),
            .I(N__11940));
    CEMux I__1709 (
            .O(N__11960),
            .I(N__11940));
    CEMux I__1708 (
            .O(N__11959),
            .I(N__11940));
    GlobalMux I__1707 (
            .O(N__11940),
            .I(N__11937));
    gio2CtrlBuf I__1706 (
            .O(N__11937),
            .I(frame_decoder_dv_c_0_g));
    CascadeMux I__1705 (
            .O(N__11934),
            .I(N__11931));
    InMux I__1704 (
            .O(N__11931),
            .I(N__11928));
    LocalMux I__1703 (
            .O(N__11928),
            .I(N__11925));
    Span4Mux_s3_h I__1702 (
            .O(N__11925),
            .I(N__11922));
    Span4Mux_v I__1701 (
            .O(N__11922),
            .I(N__11919));
    Odrv4 I__1700 (
            .O(N__11919),
            .I(frame_decoder_OFF3data_1));
    CEMux I__1699 (
            .O(N__11916),
            .I(N__11913));
    LocalMux I__1698 (
            .O(N__11913),
            .I(N__11909));
    CEMux I__1697 (
            .O(N__11912),
            .I(N__11906));
    Span4Mux_v I__1696 (
            .O(N__11909),
            .I(N__11903));
    LocalMux I__1695 (
            .O(N__11906),
            .I(N__11900));
    Odrv4 I__1694 (
            .O(N__11903),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    Odrv4 I__1693 (
            .O(N__11900),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    InMux I__1692 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__1691 (
            .O(N__11892),
            .I(\uart_sync.aux_2__0_Z0Z_0 ));
    InMux I__1690 (
            .O(N__11889),
            .I(N__11886));
    LocalMux I__1689 (
            .O(N__11886),
            .I(N__11883));
    Odrv12 I__1688 (
            .O(N__11883),
            .I(\uart_sync.aux_3__0_Z0Z_0 ));
    InMux I__1687 (
            .O(N__11880),
            .I(N__11877));
    LocalMux I__1686 (
            .O(N__11877),
            .I(N__11874));
    Odrv4 I__1685 (
            .O(N__11874),
            .I(scaler_4_data_14));
    InMux I__1684 (
            .O(N__11871),
            .I(bfn_3_27_0_));
    CascadeMux I__1683 (
            .O(N__11868),
            .I(N__11865));
    InMux I__1682 (
            .O(N__11865),
            .I(N__11862));
    LocalMux I__1681 (
            .O(N__11862),
            .I(\scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__1680 (
            .O(N__11859),
            .I(N__11854));
    CascadeMux I__1679 (
            .O(N__11858),
            .I(N__11851));
    InMux I__1678 (
            .O(N__11857),
            .I(N__11847));
    LocalMux I__1677 (
            .O(N__11854),
            .I(N__11844));
    InMux I__1676 (
            .O(N__11851),
            .I(N__11839));
    InMux I__1675 (
            .O(N__11850),
            .I(N__11839));
    LocalMux I__1674 (
            .O(N__11847),
            .I(\scaler_1.un2_source_data_0 ));
    Odrv4 I__1673 (
            .O(N__11844),
            .I(\scaler_1.un2_source_data_0 ));
    LocalMux I__1672 (
            .O(N__11839),
            .I(\scaler_1.un2_source_data_0 ));
    InMux I__1671 (
            .O(N__11832),
            .I(\scaler_1.un2_source_data_0_cry_1 ));
    CascadeMux I__1670 (
            .O(N__11829),
            .I(N__11826));
    InMux I__1669 (
            .O(N__11826),
            .I(N__11820));
    InMux I__1668 (
            .O(N__11825),
            .I(N__11820));
    LocalMux I__1667 (
            .O(N__11820),
            .I(\scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ));
    InMux I__1666 (
            .O(N__11817),
            .I(\scaler_1.un2_source_data_0_cry_2 ));
    CascadeMux I__1665 (
            .O(N__11814),
            .I(N__11811));
    InMux I__1664 (
            .O(N__11811),
            .I(N__11805));
    InMux I__1663 (
            .O(N__11810),
            .I(N__11805));
    LocalMux I__1662 (
            .O(N__11805),
            .I(\scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ));
    InMux I__1661 (
            .O(N__11802),
            .I(\scaler_1.un2_source_data_0_cry_3 ));
    CascadeMux I__1660 (
            .O(N__11799),
            .I(N__11796));
    InMux I__1659 (
            .O(N__11796),
            .I(N__11790));
    InMux I__1658 (
            .O(N__11795),
            .I(N__11790));
    LocalMux I__1657 (
            .O(N__11790),
            .I(\scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ));
    InMux I__1656 (
            .O(N__11787),
            .I(\scaler_1.un2_source_data_0_cry_4 ));
    CascadeMux I__1655 (
            .O(N__11784),
            .I(N__11781));
    InMux I__1654 (
            .O(N__11781),
            .I(N__11775));
    InMux I__1653 (
            .O(N__11780),
            .I(N__11775));
    LocalMux I__1652 (
            .O(N__11775),
            .I(\scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ));
    InMux I__1651 (
            .O(N__11772),
            .I(\scaler_1.un2_source_data_0_cry_5 ));
    CascadeMux I__1650 (
            .O(N__11769),
            .I(N__11766));
    InMux I__1649 (
            .O(N__11766),
            .I(N__11760));
    InMux I__1648 (
            .O(N__11765),
            .I(N__11760));
    LocalMux I__1647 (
            .O(N__11760),
            .I(\scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ));
    InMux I__1646 (
            .O(N__11757),
            .I(\scaler_1.un2_source_data_0_cry_6 ));
    InMux I__1645 (
            .O(N__11754),
            .I(N__11751));
    LocalMux I__1644 (
            .O(N__11751),
            .I(N__11747));
    InMux I__1643 (
            .O(N__11750),
            .I(N__11744));
    Odrv4 I__1642 (
            .O(N__11747),
            .I(frame_decoder_OFF1data_7));
    LocalMux I__1641 (
            .O(N__11744),
            .I(frame_decoder_OFF1data_7));
    InMux I__1640 (
            .O(N__11739),
            .I(N__11736));
    LocalMux I__1639 (
            .O(N__11736),
            .I(N__11732));
    InMux I__1638 (
            .O(N__11735),
            .I(N__11729));
    Odrv4 I__1637 (
            .O(N__11732),
            .I(frame_decoder_CH1data_7));
    LocalMux I__1636 (
            .O(N__11729),
            .I(frame_decoder_CH1data_7));
    CascadeMux I__1635 (
            .O(N__11724),
            .I(N__11721));
    InMux I__1634 (
            .O(N__11721),
            .I(N__11718));
    LocalMux I__1633 (
            .O(N__11718),
            .I(N__11715));
    Odrv4 I__1632 (
            .O(N__11715),
            .I(\scaler_1.un3_source_data_0_axb_7 ));
    InMux I__1631 (
            .O(N__11712),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__1630 (
            .O(N__11709),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__1629 (
            .O(N__11706),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__1628 (
            .O(N__11703),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__1627 (
            .O(N__11700),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__1626 (
            .O(N__11697),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__1625 (
            .O(N__11694),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__1624 (
            .O(N__11691),
            .I(N__11687));
    CascadeMux I__1623 (
            .O(N__11690),
            .I(N__11684));
    LocalMux I__1622 (
            .O(N__11687),
            .I(N__11679));
    InMux I__1621 (
            .O(N__11684),
            .I(N__11674));
    InMux I__1620 (
            .O(N__11683),
            .I(N__11674));
    InMux I__1619 (
            .O(N__11682),
            .I(N__11671));
    Span4Mux_v I__1618 (
            .O(N__11679),
            .I(N__11668));
    LocalMux I__1617 (
            .O(N__11674),
            .I(N__11665));
    LocalMux I__1616 (
            .O(N__11671),
            .I(\scaler_3.un2_source_data_0 ));
    Odrv4 I__1615 (
            .O(N__11668),
            .I(\scaler_3.un2_source_data_0 ));
    Odrv4 I__1614 (
            .O(N__11665),
            .I(\scaler_3.un2_source_data_0 ));
    InMux I__1613 (
            .O(N__11658),
            .I(N__11655));
    LocalMux I__1612 (
            .O(N__11655),
            .I(N__11651));
    InMux I__1611 (
            .O(N__11654),
            .I(N__11648));
    Span4Mux_h I__1610 (
            .O(N__11651),
            .I(N__11643));
    LocalMux I__1609 (
            .O(N__11648),
            .I(N__11643));
    Span4Mux_v I__1608 (
            .O(N__11643),
            .I(N__11640));
    Odrv4 I__1607 (
            .O(N__11640),
            .I(\uart_frame_decoder.source_offset2data_1_sqmuxa ));
    CascadeMux I__1606 (
            .O(N__11637),
            .I(N__11633));
    InMux I__1605 (
            .O(N__11636),
            .I(N__11630));
    InMux I__1604 (
            .O(N__11633),
            .I(N__11627));
    LocalMux I__1603 (
            .O(N__11630),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    LocalMux I__1602 (
            .O(N__11627),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    InMux I__1601 (
            .O(N__11622),
            .I(N__11619));
    LocalMux I__1600 (
            .O(N__11619),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa ));
    CascadeMux I__1599 (
            .O(N__11616),
            .I(N__11613));
    InMux I__1598 (
            .O(N__11613),
            .I(N__11607));
    InMux I__1597 (
            .O(N__11612),
            .I(N__11607));
    LocalMux I__1596 (
            .O(N__11607),
            .I(\uart_frame_decoder.state_1Z0Z_9 ));
    InMux I__1595 (
            .O(N__11604),
            .I(N__11600));
    InMux I__1594 (
            .O(N__11603),
            .I(N__11597));
    LocalMux I__1593 (
            .O(N__11600),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    LocalMux I__1592 (
            .O(N__11597),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    InMux I__1591 (
            .O(N__11592),
            .I(N__11589));
    LocalMux I__1590 (
            .O(N__11589),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__1589 (
            .O(N__11586),
            .I(N__11577));
    InMux I__1588 (
            .O(N__11585),
            .I(N__11574));
    InMux I__1587 (
            .O(N__11584),
            .I(N__11571));
    InMux I__1586 (
            .O(N__11583),
            .I(N__11567));
    InMux I__1585 (
            .O(N__11582),
            .I(N__11564));
    InMux I__1584 (
            .O(N__11581),
            .I(N__11561));
    InMux I__1583 (
            .O(N__11580),
            .I(N__11558));
    LocalMux I__1582 (
            .O(N__11577),
            .I(N__11555));
    LocalMux I__1581 (
            .O(N__11574),
            .I(N__11548));
    LocalMux I__1580 (
            .O(N__11571),
            .I(N__11548));
    CascadeMux I__1579 (
            .O(N__11570),
            .I(N__11545));
    LocalMux I__1578 (
            .O(N__11567),
            .I(N__11533));
    LocalMux I__1577 (
            .O(N__11564),
            .I(N__11533));
    LocalMux I__1576 (
            .O(N__11561),
            .I(N__11533));
    LocalMux I__1575 (
            .O(N__11558),
            .I(N__11533));
    Span4Mux_s3_h I__1574 (
            .O(N__11555),
            .I(N__11533));
    InMux I__1573 (
            .O(N__11554),
            .I(N__11530));
    InMux I__1572 (
            .O(N__11553),
            .I(N__11527));
    Span4Mux_v I__1571 (
            .O(N__11548),
            .I(N__11524));
    InMux I__1570 (
            .O(N__11545),
            .I(N__11519));
    InMux I__1569 (
            .O(N__11544),
            .I(N__11519));
    Span4Mux_v I__1568 (
            .O(N__11533),
            .I(N__11514));
    LocalMux I__1567 (
            .O(N__11530),
            .I(N__11514));
    LocalMux I__1566 (
            .O(N__11527),
            .I(uart_data_7));
    Odrv4 I__1565 (
            .O(N__11524),
            .I(uart_data_7));
    LocalMux I__1564 (
            .O(N__11519),
            .I(uart_data_7));
    Odrv4 I__1563 (
            .O(N__11514),
            .I(uart_data_7));
    InMux I__1562 (
            .O(N__11505),
            .I(N__11502));
    LocalMux I__1561 (
            .O(N__11502),
            .I(N__11499));
    Span4Mux_s2_v I__1560 (
            .O(N__11499),
            .I(N__11495));
    InMux I__1559 (
            .O(N__11498),
            .I(N__11492));
    Span4Mux_v I__1558 (
            .O(N__11495),
            .I(N__11487));
    LocalMux I__1557 (
            .O(N__11492),
            .I(N__11487));
    Odrv4 I__1556 (
            .O(N__11487),
            .I(frame_decoder_CH4data_7));
    CEMux I__1555 (
            .O(N__11484),
            .I(N__11481));
    LocalMux I__1554 (
            .O(N__11481),
            .I(N__11478));
    Span4Mux_s3_v I__1553 (
            .O(N__11478),
            .I(N__11474));
    CEMux I__1552 (
            .O(N__11477),
            .I(N__11471));
    Span4Mux_v I__1551 (
            .O(N__11474),
            .I(N__11468));
    LocalMux I__1550 (
            .O(N__11471),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    Odrv4 I__1549 (
            .O(N__11468),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__1548 (
            .O(N__11463),
            .I(N__11460));
    LocalMux I__1547 (
            .O(N__11460),
            .I(N__11456));
    InMux I__1546 (
            .O(N__11459),
            .I(N__11453));
    Span4Mux_v I__1545 (
            .O(N__11456),
            .I(N__11448));
    LocalMux I__1544 (
            .O(N__11453),
            .I(N__11448));
    Odrv4 I__1543 (
            .O(N__11448),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa ));
    CEMux I__1542 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__1541 (
            .O(N__11442),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__1540 (
            .O(N__11439),
            .I(N__11436));
    LocalMux I__1539 (
            .O(N__11436),
            .I(N__11431));
    InMux I__1538 (
            .O(N__11435),
            .I(N__11427));
    CascadeMux I__1537 (
            .O(N__11434),
            .I(N__11424));
    Span4Mux_v I__1536 (
            .O(N__11431),
            .I(N__11421));
    InMux I__1535 (
            .O(N__11430),
            .I(N__11418));
    LocalMux I__1534 (
            .O(N__11427),
            .I(N__11415));
    InMux I__1533 (
            .O(N__11424),
            .I(N__11412));
    Odrv4 I__1532 (
            .O(N__11421),
            .I(frame_decoder_OFF1data_0));
    LocalMux I__1531 (
            .O(N__11418),
            .I(frame_decoder_OFF1data_0));
    Odrv4 I__1530 (
            .O(N__11415),
            .I(frame_decoder_OFF1data_0));
    LocalMux I__1529 (
            .O(N__11412),
            .I(frame_decoder_OFF1data_0));
    InMux I__1528 (
            .O(N__11403),
            .I(N__11399));
    InMux I__1527 (
            .O(N__11402),
            .I(N__11396));
    LocalMux I__1526 (
            .O(N__11399),
            .I(N__11391));
    LocalMux I__1525 (
            .O(N__11396),
            .I(N__11388));
    InMux I__1524 (
            .O(N__11395),
            .I(N__11385));
    InMux I__1523 (
            .O(N__11394),
            .I(N__11382));
    Span4Mux_v I__1522 (
            .O(N__11391),
            .I(N__11375));
    Span4Mux_s3_v I__1521 (
            .O(N__11388),
            .I(N__11375));
    LocalMux I__1520 (
            .O(N__11385),
            .I(N__11375));
    LocalMux I__1519 (
            .O(N__11382),
            .I(frame_decoder_CH1data_0));
    Odrv4 I__1518 (
            .O(N__11375),
            .I(frame_decoder_CH1data_0));
    CascadeMux I__1517 (
            .O(N__11370),
            .I(N__11367));
    InMux I__1516 (
            .O(N__11367),
            .I(N__11361));
    InMux I__1515 (
            .O(N__11366),
            .I(N__11361));
    LocalMux I__1514 (
            .O(N__11361),
            .I(\scaler_2.un3_source_data_0_cry_1_c_RNILSPH ));
    InMux I__1513 (
            .O(N__11358),
            .I(\scaler_2.un2_source_data_0_cry_2 ));
    CascadeMux I__1512 (
            .O(N__11355),
            .I(N__11352));
    InMux I__1511 (
            .O(N__11352),
            .I(N__11346));
    InMux I__1510 (
            .O(N__11351),
            .I(N__11346));
    LocalMux I__1509 (
            .O(N__11346),
            .I(\scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ));
    InMux I__1508 (
            .O(N__11343),
            .I(\scaler_2.un2_source_data_0_cry_3 ));
    CascadeMux I__1507 (
            .O(N__11340),
            .I(N__11337));
    InMux I__1506 (
            .O(N__11337),
            .I(N__11331));
    InMux I__1505 (
            .O(N__11336),
            .I(N__11331));
    LocalMux I__1504 (
            .O(N__11331),
            .I(\scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ));
    InMux I__1503 (
            .O(N__11328),
            .I(\scaler_2.un2_source_data_0_cry_4 ));
    CascadeMux I__1502 (
            .O(N__11325),
            .I(N__11322));
    InMux I__1501 (
            .O(N__11322),
            .I(N__11316));
    InMux I__1500 (
            .O(N__11321),
            .I(N__11316));
    LocalMux I__1499 (
            .O(N__11316),
            .I(\scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ));
    InMux I__1498 (
            .O(N__11313),
            .I(\scaler_2.un2_source_data_0_cry_5 ));
    CascadeMux I__1497 (
            .O(N__11310),
            .I(N__11307));
    InMux I__1496 (
            .O(N__11307),
            .I(N__11301));
    InMux I__1495 (
            .O(N__11306),
            .I(N__11301));
    LocalMux I__1494 (
            .O(N__11301),
            .I(\scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ));
    InMux I__1493 (
            .O(N__11298),
            .I(\scaler_2.un2_source_data_0_cry_6 ));
    CascadeMux I__1492 (
            .O(N__11295),
            .I(N__11292));
    InMux I__1491 (
            .O(N__11292),
            .I(N__11286));
    InMux I__1490 (
            .O(N__11291),
            .I(N__11286));
    LocalMux I__1489 (
            .O(N__11286),
            .I(\scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ));
    InMux I__1488 (
            .O(N__11283),
            .I(\scaler_2.un2_source_data_0_cry_7 ));
    InMux I__1487 (
            .O(N__11280),
            .I(N__11276));
    InMux I__1486 (
            .O(N__11279),
            .I(N__11273));
    LocalMux I__1485 (
            .O(N__11276),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ));
    LocalMux I__1484 (
            .O(N__11273),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ));
    CascadeMux I__1483 (
            .O(N__11268),
            .I(N__11265));
    InMux I__1482 (
            .O(N__11265),
            .I(N__11262));
    LocalMux I__1481 (
            .O(N__11262),
            .I(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ));
    InMux I__1480 (
            .O(N__11259),
            .I(bfn_3_22_0_));
    InMux I__1479 (
            .O(N__11256),
            .I(\scaler_2.un2_source_data_0_cry_9 ));
    InMux I__1478 (
            .O(N__11253),
            .I(N__11249));
    InMux I__1477 (
            .O(N__11252),
            .I(N__11246));
    LocalMux I__1476 (
            .O(N__11249),
            .I(N__11236));
    LocalMux I__1475 (
            .O(N__11246),
            .I(N__11236));
    InMux I__1474 (
            .O(N__11245),
            .I(N__11233));
    InMux I__1473 (
            .O(N__11244),
            .I(N__11230));
    InMux I__1472 (
            .O(N__11243),
            .I(N__11227));
    InMux I__1471 (
            .O(N__11242),
            .I(N__11224));
    InMux I__1470 (
            .O(N__11241),
            .I(N__11221));
    Span4Mux_v I__1469 (
            .O(N__11236),
            .I(N__11217));
    LocalMux I__1468 (
            .O(N__11233),
            .I(N__11214));
    LocalMux I__1467 (
            .O(N__11230),
            .I(N__11204));
    LocalMux I__1466 (
            .O(N__11227),
            .I(N__11204));
    LocalMux I__1465 (
            .O(N__11224),
            .I(N__11204));
    LocalMux I__1464 (
            .O(N__11221),
            .I(N__11201));
    InMux I__1463 (
            .O(N__11220),
            .I(N__11198));
    Span4Mux_v I__1462 (
            .O(N__11217),
            .I(N__11195));
    Span4Mux_s3_h I__1461 (
            .O(N__11214),
            .I(N__11192));
    InMux I__1460 (
            .O(N__11213),
            .I(N__11189));
    InMux I__1459 (
            .O(N__11212),
            .I(N__11184));
    InMux I__1458 (
            .O(N__11211),
            .I(N__11184));
    Span4Mux_v I__1457 (
            .O(N__11204),
            .I(N__11177));
    Span4Mux_s3_h I__1456 (
            .O(N__11201),
            .I(N__11177));
    LocalMux I__1455 (
            .O(N__11198),
            .I(N__11177));
    Odrv4 I__1454 (
            .O(N__11195),
            .I(uart_data_0));
    Odrv4 I__1453 (
            .O(N__11192),
            .I(uart_data_0));
    LocalMux I__1452 (
            .O(N__11189),
            .I(uart_data_0));
    LocalMux I__1451 (
            .O(N__11184),
            .I(uart_data_0));
    Odrv4 I__1450 (
            .O(N__11177),
            .I(uart_data_0));
    InMux I__1449 (
            .O(N__11166),
            .I(N__11162));
    CascadeMux I__1448 (
            .O(N__11165),
            .I(N__11158));
    LocalMux I__1447 (
            .O(N__11162),
            .I(N__11155));
    CascadeMux I__1446 (
            .O(N__11161),
            .I(N__11152));
    InMux I__1445 (
            .O(N__11158),
            .I(N__11147));
    Span4Mux_h I__1444 (
            .O(N__11155),
            .I(N__11144));
    InMux I__1443 (
            .O(N__11152),
            .I(N__11137));
    InMux I__1442 (
            .O(N__11151),
            .I(N__11137));
    InMux I__1441 (
            .O(N__11150),
            .I(N__11137));
    LocalMux I__1440 (
            .O(N__11147),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    Odrv4 I__1439 (
            .O(N__11144),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__1438 (
            .O(N__11137),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    CascadeMux I__1437 (
            .O(N__11130),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ));
    InMux I__1436 (
            .O(N__11127),
            .I(N__11124));
    LocalMux I__1435 (
            .O(N__11124),
            .I(N__11120));
    InMux I__1434 (
            .O(N__11123),
            .I(N__11117));
    Odrv4 I__1433 (
            .O(N__11120),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ));
    LocalMux I__1432 (
            .O(N__11117),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ));
    InMux I__1431 (
            .O(N__11112),
            .I(N__11108));
    CascadeMux I__1430 (
            .O(N__11111),
            .I(N__11105));
    LocalMux I__1429 (
            .O(N__11108),
            .I(N__11102));
    InMux I__1428 (
            .O(N__11105),
            .I(N__11099));
    Odrv4 I__1427 (
            .O(N__11102),
            .I(\uart.data_AuxZ0Z_5 ));
    LocalMux I__1426 (
            .O(N__11099),
            .I(\uart.data_AuxZ0Z_5 ));
    InMux I__1425 (
            .O(N__11094),
            .I(N__11090));
    InMux I__1424 (
            .O(N__11093),
            .I(N__11087));
    LocalMux I__1423 (
            .O(N__11090),
            .I(N__11076));
    LocalMux I__1422 (
            .O(N__11087),
            .I(N__11076));
    InMux I__1421 (
            .O(N__11086),
            .I(N__11073));
    InMux I__1420 (
            .O(N__11085),
            .I(N__11070));
    InMux I__1419 (
            .O(N__11084),
            .I(N__11067));
    InMux I__1418 (
            .O(N__11083),
            .I(N__11064));
    InMux I__1417 (
            .O(N__11082),
            .I(N__11061));
    CascadeMux I__1416 (
            .O(N__11081),
            .I(N__11058));
    Span4Mux_v I__1415 (
            .O(N__11076),
            .I(N__11051));
    LocalMux I__1414 (
            .O(N__11073),
            .I(N__11051));
    LocalMux I__1413 (
            .O(N__11070),
            .I(N__11051));
    LocalMux I__1412 (
            .O(N__11067),
            .I(N__11048));
    LocalMux I__1411 (
            .O(N__11064),
            .I(N__11040));
    LocalMux I__1410 (
            .O(N__11061),
            .I(N__11040));
    InMux I__1409 (
            .O(N__11058),
            .I(N__11037));
    Span4Mux_v I__1408 (
            .O(N__11051),
            .I(N__11034));
    Span4Mux_s3_h I__1407 (
            .O(N__11048),
            .I(N__11031));
    InMux I__1406 (
            .O(N__11047),
            .I(N__11028));
    InMux I__1405 (
            .O(N__11046),
            .I(N__11023));
    InMux I__1404 (
            .O(N__11045),
            .I(N__11023));
    Span4Mux_v I__1403 (
            .O(N__11040),
            .I(N__11018));
    LocalMux I__1402 (
            .O(N__11037),
            .I(N__11018));
    Odrv4 I__1401 (
            .O(N__11034),
            .I(uart_data_5));
    Odrv4 I__1400 (
            .O(N__11031),
            .I(uart_data_5));
    LocalMux I__1399 (
            .O(N__11028),
            .I(uart_data_5));
    LocalMux I__1398 (
            .O(N__11023),
            .I(uart_data_5));
    Odrv4 I__1397 (
            .O(N__11018),
            .I(uart_data_5));
    InMux I__1396 (
            .O(N__11007),
            .I(N__11004));
    LocalMux I__1395 (
            .O(N__11004),
            .I(N__11000));
    CascadeMux I__1394 (
            .O(N__11003),
            .I(N__10997));
    Span4Mux_v I__1393 (
            .O(N__11000),
            .I(N__10994));
    InMux I__1392 (
            .O(N__10997),
            .I(N__10991));
    Odrv4 I__1391 (
            .O(N__10994),
            .I(\uart.data_AuxZ1Z_2 ));
    LocalMux I__1390 (
            .O(N__10991),
            .I(\uart.data_AuxZ1Z_2 ));
    InMux I__1389 (
            .O(N__10986),
            .I(N__10982));
    InMux I__1388 (
            .O(N__10985),
            .I(N__10979));
    LocalMux I__1387 (
            .O(N__10982),
            .I(N__10969));
    LocalMux I__1386 (
            .O(N__10979),
            .I(N__10969));
    InMux I__1385 (
            .O(N__10978),
            .I(N__10966));
    InMux I__1384 (
            .O(N__10977),
            .I(N__10963));
    InMux I__1383 (
            .O(N__10976),
            .I(N__10960));
    InMux I__1382 (
            .O(N__10975),
            .I(N__10957));
    InMux I__1381 (
            .O(N__10974),
            .I(N__10954));
    Span4Mux_v I__1380 (
            .O(N__10969),
            .I(N__10946));
    LocalMux I__1379 (
            .O(N__10966),
            .I(N__10946));
    LocalMux I__1378 (
            .O(N__10963),
            .I(N__10946));
    LocalMux I__1377 (
            .O(N__10960),
            .I(N__10936));
    LocalMux I__1376 (
            .O(N__10957),
            .I(N__10936));
    LocalMux I__1375 (
            .O(N__10954),
            .I(N__10936));
    InMux I__1374 (
            .O(N__10953),
            .I(N__10933));
    Span4Mux_v I__1373 (
            .O(N__10946),
            .I(N__10930));
    InMux I__1372 (
            .O(N__10945),
            .I(N__10927));
    InMux I__1371 (
            .O(N__10944),
            .I(N__10922));
    InMux I__1370 (
            .O(N__10943),
            .I(N__10922));
    Span4Mux_v I__1369 (
            .O(N__10936),
            .I(N__10917));
    LocalMux I__1368 (
            .O(N__10933),
            .I(N__10917));
    Odrv4 I__1367 (
            .O(N__10930),
            .I(uart_data_2));
    LocalMux I__1366 (
            .O(N__10927),
            .I(uart_data_2));
    LocalMux I__1365 (
            .O(N__10922),
            .I(uart_data_2));
    Odrv4 I__1364 (
            .O(N__10917),
            .I(uart_data_2));
    InMux I__1363 (
            .O(N__10908),
            .I(N__10905));
    LocalMux I__1362 (
            .O(N__10905),
            .I(N__10901));
    InMux I__1361 (
            .O(N__10904),
            .I(N__10898));
    Odrv4 I__1360 (
            .O(N__10901),
            .I(\uart.data_AuxZ0Z_7 ));
    LocalMux I__1359 (
            .O(N__10898),
            .I(\uart.data_AuxZ0Z_7 ));
    InMux I__1358 (
            .O(N__10893),
            .I(N__10890));
    LocalMux I__1357 (
            .O(N__10890),
            .I(N__10886));
    InMux I__1356 (
            .O(N__10889),
            .I(N__10883));
    Odrv12 I__1355 (
            .O(N__10886),
            .I(\uart.data_AuxZ1Z_1 ));
    LocalMux I__1354 (
            .O(N__10883),
            .I(\uart.data_AuxZ1Z_1 ));
    InMux I__1353 (
            .O(N__10878),
            .I(\scaler_2.un2_source_data_0_cry_1 ));
    CascadeMux I__1352 (
            .O(N__10875),
            .I(N__10872));
    InMux I__1351 (
            .O(N__10872),
            .I(N__10869));
    LocalMux I__1350 (
            .O(N__10869),
            .I(N__10866));
    Odrv12 I__1349 (
            .O(N__10866),
            .I(\uart.N_177 ));
    CascadeMux I__1348 (
            .O(N__10863),
            .I(\uart.state_srsts_0_0_0_cascade_ ));
    InMux I__1347 (
            .O(N__10860),
            .I(N__10857));
    LocalMux I__1346 (
            .O(N__10857),
            .I(N__10853));
    InMux I__1345 (
            .O(N__10856),
            .I(N__10850));
    Odrv4 I__1344 (
            .O(N__10853),
            .I(\uart_frame_decoder.state_1_RNI592GZ0Z_10 ));
    LocalMux I__1343 (
            .O(N__10850),
            .I(\uart_frame_decoder.state_1_RNI592GZ0Z_10 ));
    InMux I__1342 (
            .O(N__10845),
            .I(N__10842));
    LocalMux I__1341 (
            .O(N__10842),
            .I(\uart_frame_decoder.state_1_RNO_3Z0Z_0 ));
    InMux I__1340 (
            .O(N__10839),
            .I(N__10836));
    LocalMux I__1339 (
            .O(N__10836),
            .I(\uart_frame_decoder.N_168_i_1 ));
    CascadeMux I__1338 (
            .O(N__10833),
            .I(N__10830));
    InMux I__1337 (
            .O(N__10830),
            .I(N__10827));
    LocalMux I__1336 (
            .O(N__10827),
            .I(\uart_frame_decoder.state_1_RNO_2Z0Z_0 ));
    InMux I__1335 (
            .O(N__10824),
            .I(N__10820));
    InMux I__1334 (
            .O(N__10823),
            .I(N__10817));
    LocalMux I__1333 (
            .O(N__10820),
            .I(N__10814));
    LocalMux I__1332 (
            .O(N__10817),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    Odrv4 I__1331 (
            .O(N__10814),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    InMux I__1330 (
            .O(N__10809),
            .I(N__10800));
    InMux I__1329 (
            .O(N__10808),
            .I(N__10800));
    InMux I__1328 (
            .O(N__10807),
            .I(N__10800));
    LocalMux I__1327 (
            .O(N__10800),
            .I(N__10797));
    Odrv4 I__1326 (
            .O(N__10797),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    InMux I__1325 (
            .O(N__10794),
            .I(N__10788));
    InMux I__1324 (
            .O(N__10793),
            .I(N__10788));
    LocalMux I__1323 (
            .O(N__10788),
            .I(N__10785));
    Span4Mux_v I__1322 (
            .O(N__10785),
            .I(N__10782));
    Odrv4 I__1321 (
            .O(N__10782),
            .I(\uart_frame_decoder.N_79_4 ));
    InMux I__1320 (
            .O(N__10779),
            .I(N__10776));
    LocalMux I__1319 (
            .O(N__10776),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ));
    InMux I__1318 (
            .O(N__10773),
            .I(N__10769));
    CascadeMux I__1317 (
            .O(N__10772),
            .I(N__10766));
    LocalMux I__1316 (
            .O(N__10769),
            .I(N__10763));
    InMux I__1315 (
            .O(N__10766),
            .I(N__10760));
    Odrv4 I__1314 (
            .O(N__10763),
            .I(\uart.data_AuxZ1Z_0 ));
    LocalMux I__1313 (
            .O(N__10760),
            .I(\uart.data_AuxZ1Z_0 ));
    InMux I__1312 (
            .O(N__10755),
            .I(N__10752));
    LocalMux I__1311 (
            .O(N__10752),
            .I(N__10749));
    Odrv4 I__1310 (
            .O(N__10749),
            .I(\uart.data_Auxce_0_0_0 ));
    CascadeMux I__1309 (
            .O(N__10746),
            .I(N__10743));
    InMux I__1308 (
            .O(N__10743),
            .I(N__10740));
    LocalMux I__1307 (
            .O(N__10740),
            .I(N__10737));
    Odrv4 I__1306 (
            .O(N__10737),
            .I(\uart.data_Auxce_0_1 ));
    InMux I__1305 (
            .O(N__10734),
            .I(N__10731));
    LocalMux I__1304 (
            .O(N__10731),
            .I(N__10728));
    Odrv4 I__1303 (
            .O(N__10728),
            .I(\uart.data_Auxce_0_3 ));
    InMux I__1302 (
            .O(N__10725),
            .I(N__10722));
    LocalMux I__1301 (
            .O(N__10722),
            .I(N__10719));
    Odrv4 I__1300 (
            .O(N__10719),
            .I(\uart.data_Auxce_0_5 ));
    InMux I__1299 (
            .O(N__10716),
            .I(N__10713));
    LocalMux I__1298 (
            .O(N__10713),
            .I(N__10710));
    Odrv4 I__1297 (
            .O(N__10710),
            .I(\uart.data_Auxce_0_6 ));
    InMux I__1296 (
            .O(N__10707),
            .I(N__10704));
    LocalMux I__1295 (
            .O(N__10704),
            .I(\uart.CO1 ));
    CascadeMux I__1294 (
            .O(N__10701),
            .I(N__10697));
    CascadeMux I__1293 (
            .O(N__10700),
            .I(N__10694));
    InMux I__1292 (
            .O(N__10697),
            .I(N__10686));
    InMux I__1291 (
            .O(N__10694),
            .I(N__10686));
    InMux I__1290 (
            .O(N__10693),
            .I(N__10686));
    LocalMux I__1289 (
            .O(N__10686),
            .I(\uart.N_133_0 ));
    CascadeMux I__1288 (
            .O(N__10683),
            .I(\uart.N_177_cascade_ ));
    InMux I__1287 (
            .O(N__10680),
            .I(N__10677));
    LocalMux I__1286 (
            .O(N__10677),
            .I(\uart.state_srsts_i_0_3 ));
    CascadeMux I__1285 (
            .O(N__10674),
            .I(\uart.N_168_1_cascade_ ));
    InMux I__1284 (
            .O(N__10671),
            .I(N__10668));
    LocalMux I__1283 (
            .O(N__10668),
            .I(\uart.N_154_0 ));
    CascadeMux I__1282 (
            .O(N__10665),
            .I(N__10662));
    InMux I__1281 (
            .O(N__10662),
            .I(N__10656));
    InMux I__1280 (
            .O(N__10661),
            .I(N__10656));
    LocalMux I__1279 (
            .O(N__10656),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ));
    InMux I__1278 (
            .O(N__10653),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    CascadeMux I__1277 (
            .O(N__10650),
            .I(N__10647));
    InMux I__1276 (
            .O(N__10647),
            .I(N__10641));
    InMux I__1275 (
            .O(N__10646),
            .I(N__10641));
    LocalMux I__1274 (
            .O(N__10641),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ));
    InMux I__1273 (
            .O(N__10638),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    CascadeMux I__1272 (
            .O(N__10635),
            .I(N__10632));
    InMux I__1271 (
            .O(N__10632),
            .I(N__10626));
    InMux I__1270 (
            .O(N__10631),
            .I(N__10626));
    LocalMux I__1269 (
            .O(N__10626),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNI15MI ));
    InMux I__1268 (
            .O(N__10623),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__1267 (
            .O(N__10620),
            .I(N__10617));
    InMux I__1266 (
            .O(N__10617),
            .I(N__10611));
    InMux I__1265 (
            .O(N__10616),
            .I(N__10611));
    LocalMux I__1264 (
            .O(N__10611),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNI49NI ));
    InMux I__1263 (
            .O(N__10608),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__1262 (
            .O(N__10605),
            .I(N__10602));
    InMux I__1261 (
            .O(N__10602),
            .I(N__10596));
    InMux I__1260 (
            .O(N__10601),
            .I(N__10596));
    LocalMux I__1259 (
            .O(N__10596),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ));
    InMux I__1258 (
            .O(N__10593),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__1257 (
            .O(N__10590),
            .I(N__10587));
    InMux I__1256 (
            .O(N__10587),
            .I(N__10581));
    InMux I__1255 (
            .O(N__10586),
            .I(N__10581));
    LocalMux I__1254 (
            .O(N__10581),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ));
    InMux I__1253 (
            .O(N__10578),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__1252 (
            .O(N__10575),
            .I(N__10571));
    InMux I__1251 (
            .O(N__10574),
            .I(N__10568));
    LocalMux I__1250 (
            .O(N__10571),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ));
    LocalMux I__1249 (
            .O(N__10568),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ));
    CascadeMux I__1248 (
            .O(N__10563),
            .I(N__10560));
    InMux I__1247 (
            .O(N__10560),
            .I(N__10557));
    LocalMux I__1246 (
            .O(N__10557),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__1245 (
            .O(N__10554),
            .I(bfn_2_30_0_));
    InMux I__1244 (
            .O(N__10551),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__1243 (
            .O(N__10548),
            .I(N__10545));
    LocalMux I__1242 (
            .O(N__10545),
            .I(frame_decoder_OFF1data_6));
    CascadeMux I__1241 (
            .O(N__10542),
            .I(N__10539));
    InMux I__1240 (
            .O(N__10539),
            .I(N__10536));
    LocalMux I__1239 (
            .O(N__10536),
            .I(N__10533));
    Odrv4 I__1238 (
            .O(N__10533),
            .I(frame_decoder_CH1data_6));
    InMux I__1237 (
            .O(N__10530),
            .I(\scaler_1.un3_source_data_0_cry_5 ));
    InMux I__1236 (
            .O(N__10527),
            .I(\scaler_1.un3_source_data_0_cry_6 ));
    InMux I__1235 (
            .O(N__10524),
            .I(bfn_2_28_0_));
    InMux I__1234 (
            .O(N__10521),
            .I(\scaler_1.un3_source_data_0_cry_8 ));
    InMux I__1233 (
            .O(N__10518),
            .I(N__10515));
    LocalMux I__1232 (
            .O(N__10515),
            .I(\scaler_1.N_771_i_l_ofxZ0 ));
    InMux I__1231 (
            .O(N__10512),
            .I(N__10508));
    InMux I__1230 (
            .O(N__10511),
            .I(N__10505));
    LocalMux I__1229 (
            .O(N__10508),
            .I(N__10500));
    LocalMux I__1228 (
            .O(N__10505),
            .I(N__10497));
    InMux I__1227 (
            .O(N__10504),
            .I(N__10494));
    InMux I__1226 (
            .O(N__10503),
            .I(N__10491));
    Odrv4 I__1225 (
            .O(N__10500),
            .I(frame_decoder_CH4data_0));
    Odrv12 I__1224 (
            .O(N__10497),
            .I(frame_decoder_CH4data_0));
    LocalMux I__1223 (
            .O(N__10494),
            .I(frame_decoder_CH4data_0));
    LocalMux I__1222 (
            .O(N__10491),
            .I(frame_decoder_CH4data_0));
    CascadeMux I__1221 (
            .O(N__10482),
            .I(N__10478));
    InMux I__1220 (
            .O(N__10481),
            .I(N__10475));
    InMux I__1219 (
            .O(N__10478),
            .I(N__10470));
    LocalMux I__1218 (
            .O(N__10475),
            .I(N__10467));
    InMux I__1217 (
            .O(N__10474),
            .I(N__10464));
    InMux I__1216 (
            .O(N__10473),
            .I(N__10461));
    LocalMux I__1215 (
            .O(N__10470),
            .I(N__10458));
    Odrv12 I__1214 (
            .O(N__10467),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__1213 (
            .O(N__10464),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__1212 (
            .O(N__10461),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__1211 (
            .O(N__10458),
            .I(frame_decoder_OFF4data_0));
    CascadeMux I__1210 (
            .O(N__10449),
            .I(N__10446));
    InMux I__1209 (
            .O(N__10446),
            .I(N__10443));
    LocalMux I__1208 (
            .O(N__10443),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNO_2 ));
    InMux I__1207 (
            .O(N__10440),
            .I(N__10435));
    CascadeMux I__1206 (
            .O(N__10439),
            .I(N__10432));
    InMux I__1205 (
            .O(N__10438),
            .I(N__10428));
    LocalMux I__1204 (
            .O(N__10435),
            .I(N__10425));
    InMux I__1203 (
            .O(N__10432),
            .I(N__10420));
    InMux I__1202 (
            .O(N__10431),
            .I(N__10420));
    LocalMux I__1201 (
            .O(N__10428),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__1200 (
            .O(N__10425),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__1199 (
            .O(N__10420),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__1198 (
            .O(N__10413),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    InMux I__1197 (
            .O(N__10410),
            .I(N__10407));
    LocalMux I__1196 (
            .O(N__10407),
            .I(N__10404));
    Odrv4 I__1195 (
            .O(N__10404),
            .I(frame_decoder_CH1data_1));
    CascadeMux I__1194 (
            .O(N__10401),
            .I(N__10398));
    InMux I__1193 (
            .O(N__10398),
            .I(N__10395));
    LocalMux I__1192 (
            .O(N__10395),
            .I(frame_decoder_OFF1data_1));
    InMux I__1191 (
            .O(N__10392),
            .I(\scaler_1.un3_source_data_0_cry_0 ));
    InMux I__1190 (
            .O(N__10389),
            .I(N__10386));
    LocalMux I__1189 (
            .O(N__10386),
            .I(N__10383));
    Odrv4 I__1188 (
            .O(N__10383),
            .I(frame_decoder_CH1data_2));
    CascadeMux I__1187 (
            .O(N__10380),
            .I(N__10377));
    InMux I__1186 (
            .O(N__10377),
            .I(N__10374));
    LocalMux I__1185 (
            .O(N__10374),
            .I(frame_decoder_OFF1data_2));
    InMux I__1184 (
            .O(N__10371),
            .I(\scaler_1.un3_source_data_0_cry_1 ));
    InMux I__1183 (
            .O(N__10368),
            .I(N__10365));
    LocalMux I__1182 (
            .O(N__10365),
            .I(N__10362));
    Odrv4 I__1181 (
            .O(N__10362),
            .I(frame_decoder_CH1data_3));
    CascadeMux I__1180 (
            .O(N__10359),
            .I(N__10356));
    InMux I__1179 (
            .O(N__10356),
            .I(N__10353));
    LocalMux I__1178 (
            .O(N__10353),
            .I(frame_decoder_OFF1data_3));
    InMux I__1177 (
            .O(N__10350),
            .I(\scaler_1.un3_source_data_0_cry_2 ));
    CascadeMux I__1176 (
            .O(N__10347),
            .I(N__10344));
    InMux I__1175 (
            .O(N__10344),
            .I(N__10341));
    LocalMux I__1174 (
            .O(N__10341),
            .I(frame_decoder_OFF1data_4));
    InMux I__1173 (
            .O(N__10338),
            .I(\scaler_1.un3_source_data_0_cry_3 ));
    InMux I__1172 (
            .O(N__10335),
            .I(N__10332));
    LocalMux I__1171 (
            .O(N__10332),
            .I(N__10329));
    Odrv4 I__1170 (
            .O(N__10329),
            .I(frame_decoder_CH1data_5));
    CascadeMux I__1169 (
            .O(N__10326),
            .I(N__10323));
    InMux I__1168 (
            .O(N__10323),
            .I(N__10320));
    LocalMux I__1167 (
            .O(N__10320),
            .I(frame_decoder_OFF1data_5));
    InMux I__1166 (
            .O(N__10317),
            .I(\scaler_1.un3_source_data_0_cry_4 ));
    InMux I__1165 (
            .O(N__10314),
            .I(N__10311));
    LocalMux I__1164 (
            .O(N__10311),
            .I(frame_decoder_CH3data_1));
    InMux I__1163 (
            .O(N__10308),
            .I(N__10305));
    LocalMux I__1162 (
            .O(N__10305),
            .I(frame_decoder_CH3data_2));
    InMux I__1161 (
            .O(N__10302),
            .I(N__10299));
    LocalMux I__1160 (
            .O(N__10299),
            .I(frame_decoder_CH3data_3));
    InMux I__1159 (
            .O(N__10296),
            .I(N__10293));
    LocalMux I__1158 (
            .O(N__10293),
            .I(frame_decoder_CH3data_4));
    InMux I__1157 (
            .O(N__10290),
            .I(N__10287));
    LocalMux I__1156 (
            .O(N__10287),
            .I(frame_decoder_CH3data_5));
    InMux I__1155 (
            .O(N__10284),
            .I(N__10281));
    LocalMux I__1154 (
            .O(N__10281),
            .I(frame_decoder_CH3data_6));
    InMux I__1153 (
            .O(N__10278),
            .I(N__10274));
    InMux I__1152 (
            .O(N__10277),
            .I(N__10271));
    LocalMux I__1151 (
            .O(N__10274),
            .I(frame_decoder_CH3data_7));
    LocalMux I__1150 (
            .O(N__10271),
            .I(frame_decoder_CH3data_7));
    InMux I__1149 (
            .O(N__10266),
            .I(N__10260));
    InMux I__1148 (
            .O(N__10265),
            .I(N__10260));
    LocalMux I__1147 (
            .O(N__10260),
            .I(frame_decoder_CH2data_7));
    CascadeMux I__1146 (
            .O(N__10257),
            .I(N__10254));
    InMux I__1145 (
            .O(N__10254),
            .I(N__10248));
    InMux I__1144 (
            .O(N__10253),
            .I(N__10248));
    LocalMux I__1143 (
            .O(N__10248),
            .I(N__10245));
    Odrv4 I__1142 (
            .O(N__10245),
            .I(frame_decoder_OFF2data_7));
    InMux I__1141 (
            .O(N__10242),
            .I(N__10239));
    LocalMux I__1140 (
            .O(N__10239),
            .I(\scaler_2.N_783_i_l_ofxZ0 ));
    InMux I__1139 (
            .O(N__10236),
            .I(N__10232));
    InMux I__1138 (
            .O(N__10235),
            .I(N__10229));
    LocalMux I__1137 (
            .O(N__10232),
            .I(N__10226));
    LocalMux I__1136 (
            .O(N__10229),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa ));
    Odrv12 I__1135 (
            .O(N__10226),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa ));
    CEMux I__1134 (
            .O(N__10221),
            .I(N__10218));
    LocalMux I__1133 (
            .O(N__10218),
            .I(N__10215));
    Span4Mux_s3_h I__1132 (
            .O(N__10215),
            .I(N__10212));
    Odrv4 I__1131 (
            .O(N__10212),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    CascadeMux I__1130 (
            .O(N__10209),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    InMux I__1129 (
            .O(N__10206),
            .I(N__10203));
    LocalMux I__1128 (
            .O(N__10203),
            .I(N__10199));
    InMux I__1127 (
            .O(N__10202),
            .I(N__10196));
    Odrv4 I__1126 (
            .O(N__10199),
            .I(frame_decoder_OFF3data_7));
    LocalMux I__1125 (
            .O(N__10196),
            .I(frame_decoder_OFF3data_7));
    InMux I__1124 (
            .O(N__10191),
            .I(N__10188));
    LocalMux I__1123 (
            .O(N__10188),
            .I(\scaler_3.un3_source_data_0_axb_7 ));
    CascadeMux I__1122 (
            .O(N__10185),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ));
    CascadeMux I__1121 (
            .O(N__10182),
            .I(N__10179));
    InMux I__1120 (
            .O(N__10179),
            .I(N__10176));
    LocalMux I__1119 (
            .O(N__10176),
            .I(frame_decoder_OFF2data_4));
    InMux I__1118 (
            .O(N__10173),
            .I(\scaler_2.un3_source_data_0_cry_3 ));
    InMux I__1117 (
            .O(N__10170),
            .I(N__10167));
    LocalMux I__1116 (
            .O(N__10167),
            .I(frame_decoder_CH2data_5));
    CascadeMux I__1115 (
            .O(N__10164),
            .I(N__10161));
    InMux I__1114 (
            .O(N__10161),
            .I(N__10158));
    LocalMux I__1113 (
            .O(N__10158),
            .I(frame_decoder_OFF2data_5));
    InMux I__1112 (
            .O(N__10155),
            .I(\scaler_2.un3_source_data_0_cry_4 ));
    InMux I__1111 (
            .O(N__10152),
            .I(N__10149));
    LocalMux I__1110 (
            .O(N__10149),
            .I(frame_decoder_CH2data_6));
    CascadeMux I__1109 (
            .O(N__10146),
            .I(N__10143));
    InMux I__1108 (
            .O(N__10143),
            .I(N__10140));
    LocalMux I__1107 (
            .O(N__10140),
            .I(frame_decoder_OFF2data_6));
    InMux I__1106 (
            .O(N__10137),
            .I(\scaler_2.un3_source_data_0_cry_5 ));
    InMux I__1105 (
            .O(N__10134),
            .I(\scaler_2.un3_source_data_0_cry_6 ));
    InMux I__1104 (
            .O(N__10131),
            .I(bfn_2_22_0_));
    InMux I__1103 (
            .O(N__10128),
            .I(\scaler_2.un3_source_data_0_cry_8 ));
    InMux I__1102 (
            .O(N__10125),
            .I(N__10122));
    LocalMux I__1101 (
            .O(N__10122),
            .I(\scaler_2.un3_source_data_0_axb_7 ));
    InMux I__1100 (
            .O(N__10119),
            .I(N__10115));
    InMux I__1099 (
            .O(N__10118),
            .I(N__10112));
    LocalMux I__1098 (
            .O(N__10115),
            .I(N__10109));
    LocalMux I__1097 (
            .O(N__10112),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa ));
    Odrv12 I__1096 (
            .O(N__10109),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa ));
    CEMux I__1095 (
            .O(N__10104),
            .I(N__10101));
    LocalMux I__1094 (
            .O(N__10101),
            .I(N__10098));
    Odrv4 I__1093 (
            .O(N__10098),
            .I(\uart_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    InMux I__1092 (
            .O(N__10095),
            .I(N__10092));
    LocalMux I__1091 (
            .O(N__10092),
            .I(frame_decoder_CH2data_1));
    CascadeMux I__1090 (
            .O(N__10089),
            .I(N__10086));
    InMux I__1089 (
            .O(N__10086),
            .I(N__10083));
    LocalMux I__1088 (
            .O(N__10083),
            .I(frame_decoder_OFF2data_1));
    InMux I__1087 (
            .O(N__10080),
            .I(\scaler_2.un3_source_data_0_cry_0 ));
    InMux I__1086 (
            .O(N__10077),
            .I(N__10074));
    LocalMux I__1085 (
            .O(N__10074),
            .I(frame_decoder_CH2data_2));
    CascadeMux I__1084 (
            .O(N__10071),
            .I(N__10068));
    InMux I__1083 (
            .O(N__10068),
            .I(N__10065));
    LocalMux I__1082 (
            .O(N__10065),
            .I(N__10062));
    Odrv4 I__1081 (
            .O(N__10062),
            .I(frame_decoder_OFF2data_2));
    InMux I__1080 (
            .O(N__10059),
            .I(\scaler_2.un3_source_data_0_cry_1 ));
    InMux I__1079 (
            .O(N__10056),
            .I(N__10053));
    LocalMux I__1078 (
            .O(N__10053),
            .I(frame_decoder_CH2data_3));
    CascadeMux I__1077 (
            .O(N__10050),
            .I(N__10047));
    InMux I__1076 (
            .O(N__10047),
            .I(N__10044));
    LocalMux I__1075 (
            .O(N__10044),
            .I(frame_decoder_OFF2data_3));
    InMux I__1074 (
            .O(N__10041),
            .I(\scaler_2.un3_source_data_0_cry_2 ));
    InMux I__1073 (
            .O(N__10038),
            .I(N__10035));
    LocalMux I__1072 (
            .O(N__10035),
            .I(frame_decoder_CH2data_4));
    InMux I__1071 (
            .O(N__10032),
            .I(N__10028));
    InMux I__1070 (
            .O(N__10031),
            .I(N__10025));
    LocalMux I__1069 (
            .O(N__10028),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    LocalMux I__1068 (
            .O(N__10025),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    InMux I__1067 (
            .O(N__10020),
            .I(N__10017));
    LocalMux I__1066 (
            .O(N__10017),
            .I(N__10013));
    InMux I__1065 (
            .O(N__10016),
            .I(N__10010));
    Span4Mux_v I__1064 (
            .O(N__10013),
            .I(N__10007));
    LocalMux I__1063 (
            .O(N__10010),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    Odrv4 I__1062 (
            .O(N__10007),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    CascadeMux I__1061 (
            .O(N__10002),
            .I(N__9998));
    InMux I__1060 (
            .O(N__10001),
            .I(N__9994));
    InMux I__1059 (
            .O(N__9998),
            .I(N__9989));
    InMux I__1058 (
            .O(N__9997),
            .I(N__9989));
    LocalMux I__1057 (
            .O(N__9994),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    LocalMux I__1056 (
            .O(N__9989),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    InMux I__1055 (
            .O(N__9984),
            .I(N__9978));
    InMux I__1054 (
            .O(N__9983),
            .I(N__9971));
    InMux I__1053 (
            .O(N__9982),
            .I(N__9971));
    InMux I__1052 (
            .O(N__9981),
            .I(N__9971));
    LocalMux I__1051 (
            .O(N__9978),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    LocalMux I__1050 (
            .O(N__9971),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    CascadeMux I__1049 (
            .O(N__9966),
            .I(N__9962));
    InMux I__1048 (
            .O(N__9965),
            .I(N__9957));
    InMux I__1047 (
            .O(N__9962),
            .I(N__9954));
    InMux I__1046 (
            .O(N__9961),
            .I(N__9949));
    InMux I__1045 (
            .O(N__9960),
            .I(N__9949));
    LocalMux I__1044 (
            .O(N__9957),
            .I(\uart_frame_decoder.count8_0 ));
    LocalMux I__1043 (
            .O(N__9954),
            .I(\uart_frame_decoder.count8_0 ));
    LocalMux I__1042 (
            .O(N__9949),
            .I(\uart_frame_decoder.count8_0 ));
    CascadeMux I__1041 (
            .O(N__9942),
            .I(\uart_frame_decoder.state_1_ns_i_i_0_0_cascade_ ));
    InMux I__1040 (
            .O(N__9939),
            .I(N__9934));
    InMux I__1039 (
            .O(N__9938),
            .I(N__9929));
    InMux I__1038 (
            .O(N__9937),
            .I(N__9929));
    LocalMux I__1037 (
            .O(N__9934),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__1036 (
            .O(N__9929),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    InMux I__1035 (
            .O(N__9924),
            .I(N__9920));
    InMux I__1034 (
            .O(N__9923),
            .I(N__9917));
    LocalMux I__1033 (
            .O(N__9920),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__1032 (
            .O(N__9917),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    CascadeMux I__1031 (
            .O(N__9912),
            .I(N__9908));
    InMux I__1030 (
            .O(N__9911),
            .I(N__9905));
    InMux I__1029 (
            .O(N__9908),
            .I(N__9902));
    LocalMux I__1028 (
            .O(N__9905),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__1027 (
            .O(N__9902),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    InMux I__1026 (
            .O(N__9897),
            .I(N__9892));
    InMux I__1025 (
            .O(N__9896),
            .I(N__9887));
    InMux I__1024 (
            .O(N__9895),
            .I(N__9887));
    LocalMux I__1023 (
            .O(N__9892),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__1022 (
            .O(N__9887),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    InMux I__1021 (
            .O(N__9882),
            .I(N__9878));
    InMux I__1020 (
            .O(N__9881),
            .I(N__9875));
    LocalMux I__1019 (
            .O(N__9878),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__1018 (
            .O(N__9875),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    CascadeMux I__1017 (
            .O(N__9870),
            .I(\uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ));
    InMux I__1016 (
            .O(N__9867),
            .I(N__9864));
    LocalMux I__1015 (
            .O(N__9864),
            .I(\uart_frame_decoder.WDT8lto13_1 ));
    CascadeMux I__1014 (
            .O(N__9861),
            .I(\uart_frame_decoder.WDT8lt14_0_cascade_ ));
    CascadeMux I__1013 (
            .O(N__9858),
            .I(N__9854));
    InMux I__1012 (
            .O(N__9857),
            .I(N__9851));
    InMux I__1011 (
            .O(N__9854),
            .I(N__9848));
    LocalMux I__1010 (
            .O(N__9851),
            .I(\uart_frame_decoder.WDT8_0_i ));
    LocalMux I__1009 (
            .O(N__9848),
            .I(\uart_frame_decoder.WDT8_0_i ));
    InMux I__1008 (
            .O(N__9843),
            .I(N__9839));
    InMux I__1007 (
            .O(N__9842),
            .I(N__9836));
    LocalMux I__1006 (
            .O(N__9839),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__1005 (
            .O(N__9836),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    InMux I__1004 (
            .O(N__9831),
            .I(N__9827));
    InMux I__1003 (
            .O(N__9830),
            .I(N__9824));
    LocalMux I__1002 (
            .O(N__9827),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__1001 (
            .O(N__9824),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    CascadeMux I__1000 (
            .O(N__9819),
            .I(N__9815));
    InMux I__999 (
            .O(N__9818),
            .I(N__9812));
    InMux I__998 (
            .O(N__9815),
            .I(N__9809));
    LocalMux I__997 (
            .O(N__9812),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__996 (
            .O(N__9809),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    InMux I__995 (
            .O(N__9804),
            .I(N__9800));
    InMux I__994 (
            .O(N__9803),
            .I(N__9797));
    LocalMux I__993 (
            .O(N__9800),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__992 (
            .O(N__9797),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    InMux I__991 (
            .O(N__9792),
            .I(N__9789));
    LocalMux I__990 (
            .O(N__9789),
            .I(\uart_frame_decoder.WDT_RNIM6B11Z0Z_4 ));
    InMux I__989 (
            .O(N__9786),
            .I(N__9781));
    InMux I__988 (
            .O(N__9785),
            .I(N__9778));
    InMux I__987 (
            .O(N__9784),
            .I(N__9775));
    LocalMux I__986 (
            .O(N__9781),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__985 (
            .O(N__9778),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__984 (
            .O(N__9775),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    CascadeMux I__983 (
            .O(N__9768),
            .I(N__9764));
    InMux I__982 (
            .O(N__9767),
            .I(N__9760));
    InMux I__981 (
            .O(N__9764),
            .I(N__9757));
    InMux I__980 (
            .O(N__9763),
            .I(N__9754));
    LocalMux I__979 (
            .O(N__9760),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__978 (
            .O(N__9757),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__977 (
            .O(N__9754),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    InMux I__976 (
            .O(N__9747),
            .I(N__9744));
    LocalMux I__975 (
            .O(N__9744),
            .I(\uart_frame_decoder.WDT8lt14_0 ));
    CascadeMux I__974 (
            .O(N__9741),
            .I(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_ ));
    InMux I__973 (
            .O(N__9738),
            .I(N__9732));
    InMux I__972 (
            .O(N__9737),
            .I(N__9732));
    LocalMux I__971 (
            .O(N__9732),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    InMux I__970 (
            .O(N__9729),
            .I(N__9726));
    LocalMux I__969 (
            .O(N__9726),
            .I(N__9723));
    Span4Mux_s3_v I__968 (
            .O(N__9723),
            .I(N__9720));
    Odrv4 I__967 (
            .O(N__9720),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__966 (
            .O(N__9717),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__965 (
            .O(N__9714),
            .I(bfn_1_30_0_));
    InMux I__964 (
            .O(N__9711),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    InMux I__963 (
            .O(N__9708),
            .I(N__9704));
    InMux I__962 (
            .O(N__9707),
            .I(N__9701));
    LocalMux I__961 (
            .O(N__9704),
            .I(N__9696));
    LocalMux I__960 (
            .O(N__9701),
            .I(N__9696));
    Odrv12 I__959 (
            .O(N__9696),
            .I(frame_decoder_OFF4data_7));
    InMux I__958 (
            .O(N__9693),
            .I(N__9690));
    LocalMux I__957 (
            .O(N__9690),
            .I(\scaler_4.N_807_i_l_ofxZ0 ));
    InMux I__956 (
            .O(N__9687),
            .I(N__9683));
    InMux I__955 (
            .O(N__9686),
            .I(N__9680));
    LocalMux I__954 (
            .O(N__9683),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__953 (
            .O(N__9680),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    InMux I__952 (
            .O(N__9675),
            .I(N__9672));
    LocalMux I__951 (
            .O(N__9672),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__950 (
            .O(N__9669),
            .I(N__9666));
    InMux I__949 (
            .O(N__9666),
            .I(N__9663));
    LocalMux I__948 (
            .O(N__9663),
            .I(N__9660));
    Odrv4 I__947 (
            .O(N__9660),
            .I(frame_decoder_OFF4data_1));
    InMux I__946 (
            .O(N__9657),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__945 (
            .O(N__9654),
            .I(N__9651));
    LocalMux I__944 (
            .O(N__9651),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__943 (
            .O(N__9648),
            .I(N__9645));
    InMux I__942 (
            .O(N__9645),
            .I(N__9642));
    LocalMux I__941 (
            .O(N__9642),
            .I(N__9639));
    Odrv4 I__940 (
            .O(N__9639),
            .I(frame_decoder_OFF4data_2));
    InMux I__939 (
            .O(N__9636),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__938 (
            .O(N__9633),
            .I(N__9630));
    LocalMux I__937 (
            .O(N__9630),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__936 (
            .O(N__9627),
            .I(N__9624));
    InMux I__935 (
            .O(N__9624),
            .I(N__9621));
    LocalMux I__934 (
            .O(N__9621),
            .I(N__9618));
    Odrv4 I__933 (
            .O(N__9618),
            .I(frame_decoder_OFF4data_3));
    InMux I__932 (
            .O(N__9615),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__931 (
            .O(N__9612),
            .I(N__9609));
    LocalMux I__930 (
            .O(N__9609),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__929 (
            .O(N__9606),
            .I(N__9603));
    InMux I__928 (
            .O(N__9603),
            .I(N__9600));
    LocalMux I__927 (
            .O(N__9600),
            .I(N__9597));
    Odrv4 I__926 (
            .O(N__9597),
            .I(frame_decoder_OFF4data_4));
    InMux I__925 (
            .O(N__9594),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__924 (
            .O(N__9591),
            .I(N__9588));
    LocalMux I__923 (
            .O(N__9588),
            .I(N__9585));
    Odrv4 I__922 (
            .O(N__9585),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__921 (
            .O(N__9582),
            .I(N__9579));
    InMux I__920 (
            .O(N__9579),
            .I(N__9576));
    LocalMux I__919 (
            .O(N__9576),
            .I(frame_decoder_CH4data_5));
    InMux I__918 (
            .O(N__9573),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__917 (
            .O(N__9570),
            .I(N__9567));
    LocalMux I__916 (
            .O(N__9567),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__915 (
            .O(N__9564),
            .I(N__9561));
    InMux I__914 (
            .O(N__9561),
            .I(N__9558));
    LocalMux I__913 (
            .O(N__9558),
            .I(N__9555));
    Odrv4 I__912 (
            .O(N__9555),
            .I(frame_decoder_OFF4data_6));
    InMux I__911 (
            .O(N__9552),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    CEMux I__910 (
            .O(N__9549),
            .I(N__9546));
    LocalMux I__909 (
            .O(N__9546),
            .I(N__9543));
    Span4Mux_v I__908 (
            .O(N__9543),
            .I(N__9540));
    Odrv4 I__907 (
            .O(N__9540),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    CascadeMux I__906 (
            .O(N__9537),
            .I(N__9534));
    InMux I__905 (
            .O(N__9534),
            .I(N__9528));
    InMux I__904 (
            .O(N__9533),
            .I(N__9528));
    LocalMux I__903 (
            .O(N__9528),
            .I(N__9525));
    Odrv4 I__902 (
            .O(N__9525),
            .I(\scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ));
    InMux I__901 (
            .O(N__9522),
            .I(\scaler_3.un2_source_data_0_cry_6 ));
    CascadeMux I__900 (
            .O(N__9519),
            .I(N__9516));
    InMux I__899 (
            .O(N__9516),
            .I(N__9510));
    InMux I__898 (
            .O(N__9515),
            .I(N__9510));
    LocalMux I__897 (
            .O(N__9510),
            .I(N__9507));
    Odrv4 I__896 (
            .O(N__9507),
            .I(\scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ));
    InMux I__895 (
            .O(N__9504),
            .I(\scaler_3.un2_source_data_0_cry_7 ));
    InMux I__894 (
            .O(N__9501),
            .I(N__9498));
    LocalMux I__893 (
            .O(N__9498),
            .I(N__9494));
    InMux I__892 (
            .O(N__9497),
            .I(N__9491));
    Odrv4 I__891 (
            .O(N__9494),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ));
    LocalMux I__890 (
            .O(N__9491),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ));
    CascadeMux I__889 (
            .O(N__9486),
            .I(N__9483));
    InMux I__888 (
            .O(N__9483),
            .I(N__9480));
    LocalMux I__887 (
            .O(N__9480),
            .I(N__9477));
    Odrv4 I__886 (
            .O(N__9477),
            .I(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ));
    InMux I__885 (
            .O(N__9474),
            .I(bfn_1_26_0_));
    InMux I__884 (
            .O(N__9471),
            .I(\scaler_3.un2_source_data_0_cry_9 ));
    InMux I__883 (
            .O(N__9468),
            .I(N__9465));
    LocalMux I__882 (
            .O(N__9465),
            .I(\scaler_3.N_795_i_l_ofxZ0 ));
    CascadeMux I__881 (
            .O(N__9462),
            .I(N__9459));
    InMux I__880 (
            .O(N__9459),
            .I(N__9456));
    LocalMux I__879 (
            .O(N__9456),
            .I(\scaler_3.un2_source_data_0_cry_1_c_RNO_1 ));
    InMux I__878 (
            .O(N__9453),
            .I(\scaler_3.un2_source_data_0_cry_1 ));
    CascadeMux I__877 (
            .O(N__9450),
            .I(N__9447));
    InMux I__876 (
            .O(N__9447),
            .I(N__9441));
    InMux I__875 (
            .O(N__9446),
            .I(N__9441));
    LocalMux I__874 (
            .O(N__9441),
            .I(N__9438));
    Odrv12 I__873 (
            .O(N__9438),
            .I(\scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ));
    InMux I__872 (
            .O(N__9435),
            .I(\scaler_3.un2_source_data_0_cry_2 ));
    CascadeMux I__871 (
            .O(N__9432),
            .I(N__9429));
    InMux I__870 (
            .O(N__9429),
            .I(N__9423));
    InMux I__869 (
            .O(N__9428),
            .I(N__9423));
    LocalMux I__868 (
            .O(N__9423),
            .I(N__9420));
    Odrv4 I__867 (
            .O(N__9420),
            .I(\scaler_3.un3_source_data_0_cry_2_c_RNIR08I ));
    InMux I__866 (
            .O(N__9417),
            .I(\scaler_3.un2_source_data_0_cry_3 ));
    CascadeMux I__865 (
            .O(N__9414),
            .I(N__9411));
    InMux I__864 (
            .O(N__9411),
            .I(N__9405));
    InMux I__863 (
            .O(N__9410),
            .I(N__9405));
    LocalMux I__862 (
            .O(N__9405),
            .I(N__9402));
    Odrv4 I__861 (
            .O(N__9402),
            .I(\scaler_3.un3_source_data_0_cry_3_c_RNIU49I ));
    InMux I__860 (
            .O(N__9399),
            .I(\scaler_3.un2_source_data_0_cry_4 ));
    CascadeMux I__859 (
            .O(N__9396),
            .I(N__9393));
    InMux I__858 (
            .O(N__9393),
            .I(N__9387));
    InMux I__857 (
            .O(N__9392),
            .I(N__9387));
    LocalMux I__856 (
            .O(N__9387),
            .I(N__9384));
    Odrv4 I__855 (
            .O(N__9384),
            .I(\scaler_3.un3_source_data_0_cry_4_c_RNI19AI ));
    InMux I__854 (
            .O(N__9381),
            .I(\scaler_3.un2_source_data_0_cry_5 ));
    CascadeMux I__853 (
            .O(N__9378),
            .I(N__9375));
    InMux I__852 (
            .O(N__9375),
            .I(N__9372));
    LocalMux I__851 (
            .O(N__9372),
            .I(frame_decoder_OFF3data_3));
    InMux I__850 (
            .O(N__9369),
            .I(\scaler_3.un3_source_data_0_cry_2 ));
    CascadeMux I__849 (
            .O(N__9366),
            .I(N__9363));
    InMux I__848 (
            .O(N__9363),
            .I(N__9360));
    LocalMux I__847 (
            .O(N__9360),
            .I(frame_decoder_OFF3data_4));
    InMux I__846 (
            .O(N__9357),
            .I(\scaler_3.un3_source_data_0_cry_3 ));
    CascadeMux I__845 (
            .O(N__9354),
            .I(N__9351));
    InMux I__844 (
            .O(N__9351),
            .I(N__9348));
    LocalMux I__843 (
            .O(N__9348),
            .I(frame_decoder_OFF3data_5));
    InMux I__842 (
            .O(N__9345),
            .I(\scaler_3.un3_source_data_0_cry_4 ));
    CascadeMux I__841 (
            .O(N__9342),
            .I(N__9339));
    InMux I__840 (
            .O(N__9339),
            .I(N__9336));
    LocalMux I__839 (
            .O(N__9336),
            .I(frame_decoder_OFF3data_6));
    InMux I__838 (
            .O(N__9333),
            .I(\scaler_3.un3_source_data_0_cry_5 ));
    InMux I__837 (
            .O(N__9330),
            .I(\scaler_3.un3_source_data_0_cry_6 ));
    InMux I__836 (
            .O(N__9327),
            .I(bfn_1_24_0_));
    InMux I__835 (
            .O(N__9324),
            .I(\scaler_3.un3_source_data_0_cry_8 ));
    InMux I__834 (
            .O(N__9321),
            .I(\scaler_3.un3_source_data_0_cry_0 ));
    CascadeMux I__833 (
            .O(N__9318),
            .I(N__9315));
    InMux I__832 (
            .O(N__9315),
            .I(N__9312));
    LocalMux I__831 (
            .O(N__9312),
            .I(frame_decoder_OFF3data_2));
    InMux I__830 (
            .O(N__9309),
            .I(\scaler_3.un3_source_data_0_cry_1 ));
    InMux I__829 (
            .O(N__9306),
            .I(N__9302));
    InMux I__828 (
            .O(N__9305),
            .I(N__9299));
    LocalMux I__827 (
            .O(N__9302),
            .I(\uart_frame_decoder.count8_0_i ));
    LocalMux I__826 (
            .O(N__9299),
            .I(\uart_frame_decoder.count8_0_i ));
    InMux I__825 (
            .O(N__9294),
            .I(N__9291));
    LocalMux I__824 (
            .O(N__9291),
            .I(\uart_frame_decoder.count_i_2 ));
    InMux I__823 (
            .O(N__9288),
            .I(\uart_frame_decoder.count8 ));
    InMux I__822 (
            .O(N__9285),
            .I(N__9279));
    InMux I__821 (
            .O(N__9284),
            .I(N__9279));
    LocalMux I__820 (
            .O(N__9279),
            .I(\uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21 ));
    CascadeMux I__819 (
            .O(N__9276),
            .I(\uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_ ));
    CascadeMux I__818 (
            .O(N__9273),
            .I(N__9269));
    InMux I__817 (
            .O(N__9272),
            .I(N__9264));
    InMux I__816 (
            .O(N__9269),
            .I(N__9264));
    LocalMux I__815 (
            .O(N__9264),
            .I(\uart_frame_decoder.count_RNIV5MSZ0Z_0 ));
    SRMux I__814 (
            .O(N__9261),
            .I(N__9258));
    LocalMux I__813 (
            .O(N__9258),
            .I(N__9254));
    SRMux I__812 (
            .O(N__9257),
            .I(N__9251));
    Span4Mux_v I__811 (
            .O(N__9254),
            .I(N__9246));
    LocalMux I__810 (
            .O(N__9251),
            .I(N__9246));
    Odrv4 I__809 (
            .O(N__9246),
            .I(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__808 (
            .O(N__9243),
            .I(\uart_frame_decoder.un1_WDT_cry_8 ));
    InMux I__807 (
            .O(N__9240),
            .I(\uart_frame_decoder.un1_WDT_cry_9 ));
    InMux I__806 (
            .O(N__9237),
            .I(\uart_frame_decoder.un1_WDT_cry_10 ));
    InMux I__805 (
            .O(N__9234),
            .I(\uart_frame_decoder.un1_WDT_cry_11 ));
    InMux I__804 (
            .O(N__9231),
            .I(\uart_frame_decoder.un1_WDT_cry_12 ));
    InMux I__803 (
            .O(N__9228),
            .I(\uart_frame_decoder.un1_WDT_cry_13 ));
    InMux I__802 (
            .O(N__9225),
            .I(\uart_frame_decoder.un1_WDT_cry_14 ));
    InMux I__801 (
            .O(N__9222),
            .I(N__9219));
    LocalMux I__800 (
            .O(N__9219),
            .I(\uart_frame_decoder.count8_axb_1 ));
    InMux I__799 (
            .O(N__9216),
            .I(N__9213));
    LocalMux I__798 (
            .O(N__9213),
            .I(\uart_frame_decoder.WDTZ0Z_1 ));
    InMux I__797 (
            .O(N__9210),
            .I(\uart_frame_decoder.un1_WDT_cry_0 ));
    InMux I__796 (
            .O(N__9207),
            .I(N__9204));
    LocalMux I__795 (
            .O(N__9204),
            .I(\uart_frame_decoder.WDTZ0Z_2 ));
    InMux I__794 (
            .O(N__9201),
            .I(\uart_frame_decoder.un1_WDT_cry_1 ));
    InMux I__793 (
            .O(N__9198),
            .I(N__9195));
    LocalMux I__792 (
            .O(N__9195),
            .I(\uart_frame_decoder.WDTZ0Z_3 ));
    InMux I__791 (
            .O(N__9192),
            .I(\uart_frame_decoder.un1_WDT_cry_2 ));
    InMux I__790 (
            .O(N__9189),
            .I(\uart_frame_decoder.un1_WDT_cry_3 ));
    InMux I__789 (
            .O(N__9186),
            .I(\uart_frame_decoder.un1_WDT_cry_4 ));
    InMux I__788 (
            .O(N__9183),
            .I(\uart_frame_decoder.un1_WDT_cry_5 ));
    InMux I__787 (
            .O(N__9180),
            .I(\uart_frame_decoder.un1_WDT_cry_6 ));
    InMux I__786 (
            .O(N__9177),
            .I(bfn_1_18_0_));
    InMux I__785 (
            .O(N__9174),
            .I(N__9171));
    LocalMux I__784 (
            .O(N__9171),
            .I(\uart_frame_decoder.WDTZ0Z_0 ));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(\scaler_3.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(\scaler_3.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(\scaler_2.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_3_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_22_0_ (
            .carryinitin(\scaler_2.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_3_22_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_27_0_));
    defparam IN_MUX_bfv_2_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_28_0_ (
            .carryinitin(\scaler_1.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_2_28_0_));
    defparam IN_MUX_bfv_3_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(\scaler_1.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_4_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_29_0_));
    defparam IN_MUX_bfv_4_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_13 ),
            .carryinitout(bfn_4_30_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_3_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_3_27_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_4_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_28_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_13 ),
            .carryinitout(bfn_4_28_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_4_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_13 ),
            .carryinitout(bfn_4_25_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\uart_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_11_26_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__24524),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB frame_decoder_dv_c_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__14886),
            .GLOBALBUFFEROUTPUT(frame_decoder_dv_c_0_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__20943),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_238_i_0_g ));
    GND GND (
            .Y(GNDG0));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24360),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_512_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uart_frame_decoder.WDT_0_LC_1_17_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_0_LC_1_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_0_LC_1_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_0_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__9174),
            .in2(N__9858),
            .in3(N__9857),
            .lcout(\uart_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_1_LC_1_17_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_1_LC_1_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_1_LC_1_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_1_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__9216),
            .in2(_gnd_net_),
            .in3(N__9210),
            .lcout(\uart_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_2_LC_1_17_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_2_LC_1_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_2_LC_1_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_2_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__9207),
            .in2(_gnd_net_),
            .in3(N__9201),
            .lcout(\uart_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_3_LC_1_17_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_3_LC_1_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_3_LC_1_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_3_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__9198),
            .in2(_gnd_net_),
            .in3(N__9192),
            .lcout(\uart_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_4_LC_1_17_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_4_LC_1_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_4_LC_1_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_4_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__9804),
            .in2(_gnd_net_),
            .in3(N__9189),
            .lcout(\uart_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_5_LC_1_17_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_5_LC_1_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_5_LC_1_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_5_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__9831),
            .in2(_gnd_net_),
            .in3(N__9186),
            .lcout(\uart_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_6_LC_1_17_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_6_LC_1_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_6_LC_1_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_6_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__9843),
            .in2(_gnd_net_),
            .in3(N__9183),
            .lcout(\uart_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_7_LC_1_17_7 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_7_LC_1_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_7_LC_1_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_7_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__9818),
            .in2(_gnd_net_),
            .in3(N__9180),
            .lcout(\uart_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__23875),
            .ce(),
            .sr(N__9261));
    defparam \uart_frame_decoder.WDT_8_LC_1_18_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_8_LC_1_18_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_8_LC_1_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_8_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__9687),
            .in2(_gnd_net_),
            .in3(N__9177),
            .lcout(\uart_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_9_LC_1_18_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_9_LC_1_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_9_LC_1_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_9_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__9882),
            .in2(_gnd_net_),
            .in3(N__9243),
            .lcout(\uart_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_10_LC_1_18_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_10_LC_1_18_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_10_LC_1_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_10_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__9924),
            .in2(_gnd_net_),
            .in3(N__9240),
            .lcout(\uart_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_11_LC_1_18_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_11_LC_1_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_11_LC_1_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_11_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__9939),
            .in2(_gnd_net_),
            .in3(N__9237),
            .lcout(\uart_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_12_LC_1_18_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_12_LC_1_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_12_LC_1_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_12_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__9897),
            .in2(_gnd_net_),
            .in3(N__9234),
            .lcout(\uart_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_13_LC_1_18_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_13_LC_1_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_13_LC_1_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_13_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__9911),
            .in2(_gnd_net_),
            .in3(N__9231),
            .lcout(\uart_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_14_LC_1_18_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_14_LC_1_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_14_LC_1_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_14_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__9767),
            .in2(_gnd_net_),
            .in3(N__9228),
            .lcout(\uart_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.WDT_15_LC_1_18_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_15_LC_1_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_15_LC_1_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_frame_decoder.WDT_15_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__9786),
            .in2(_gnd_net_),
            .in3(N__9225),
            .lcout(\uart_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23871),
            .ce(),
            .sr(N__9257));
    defparam \uart_frame_decoder.count8_cry_0_c_LC_1_19_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_1_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__9305),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\uart_frame_decoder.count8_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_1_19_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_1_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_1_c_inv_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__9222),
            .in2(_gnd_net_),
            .in3(N__9981),
            .lcout(\uart_frame_decoder.count8_axb_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_0 ),
            .carryout(\uart_frame_decoder.count8_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_1_19_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_1_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_inv_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__9294),
            .in2(N__24690),
            .in3(N__9997),
            .lcout(\uart_frame_decoder.count_i_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_1 ),
            .carryout(\uart_frame_decoder.count8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_1_19_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_1_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.count8_THRU_LUT4_0_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9288),
            .lcout(\uart_frame_decoder.count8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_1_LC_1_19_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_1_LC_1_19_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_1_LC_1_19_4 .LUT_INIT=16'b0000000010100101;
    LogicCell40 \uart_frame_decoder.count_1_LC_1_19_4  (
            .in0(N__9982),
            .in1(_gnd_net_),
            .in2(N__9273),
            .in3(N__9284),
            .lcout(\uart_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23866),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_2_LC_1_19_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_2_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_2_LC_1_19_5 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \uart_frame_decoder.count_2_LC_1_19_5  (
            .in0(N__9285),
            .in1(N__9272),
            .in2(N__10002),
            .in3(N__9983),
            .lcout(\uart_frame_decoder.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23866),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_1_19_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_1_19_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_1_19_6  (
            .in0(N__13116),
            .in1(N__24507),
            .in2(N__13173),
            .in3(N__13004),
            .lcout(\uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21 ),
            .ltout(\uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_0_LC_1_19_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_0_LC_1_19_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_0_LC_1_19_7 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \uart_frame_decoder.count_0_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__10860),
            .in2(N__9276),
            .in3(N__9965),
            .lcout(\uart_frame_decoder.count8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23866),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.source_data_1_4_LC_1_20_0 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_4_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_4_LC_1_20_0 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \scaler_1.source_data_1_4_LC_1_20_0  (
            .in0(N__11403),
            .in1(N__14946),
            .in2(N__16067),
            .in3(N__11439),
            .lcout(scaler_1_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23862),
            .ce(),
            .sr(N__23358));
    defparam \scaler_4.source_data_1_4_LC_1_20_3 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_1_20_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_1_20_3  (
            .in0(N__14947),
            .in1(N__10481),
            .in2(N__16091),
            .in3(N__10511),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23862),
            .ce(),
            .sr(N__23358));
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_1_20_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_1_20_5 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \uart_frame_decoder.count_RNIV5MS_0_LC_1_20_5  (
            .in0(N__13172),
            .in1(_gnd_net_),
            .in2(N__13119),
            .in3(N__9961),
            .lcout(\uart_frame_decoder.count_RNIV5MSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_1_20_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_1_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__13112),
            .in2(_gnd_net_),
            .in3(N__23496),
            .lcout(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_1_20_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_1_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_inv_LC_1_20_7  (
            .in0(N__9306),
            .in1(N__24716),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(\uart_frame_decoder.count8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_1_21_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_1_21_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_1_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_0_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11245),
            .lcout(frame_decoder_CH2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_1_21_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_1_21_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_1_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_1_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12777),
            .lcout(frame_decoder_CH2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_1_21_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_1_21_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_1_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_2_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10977),
            .lcout(frame_decoder_CH2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_1_21_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_1_21_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_1_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_3_LC_1_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12528),
            .lcout(frame_decoder_CH2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_1_21_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_1_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_4_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15093),
            .lcout(frame_decoder_CH2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_1_21_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_1_21_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_1_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_5_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11084),
            .lcout(frame_decoder_CH2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_1_21_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_1_21_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_1_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_6_LC_1_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12438),
            .lcout(frame_decoder_CH2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_1_21_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_1_21_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_1_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_7_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11584),
            .lcout(frame_decoder_CH2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23857),
            .ce(N__10221),
            .sr(N__23362));
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_1_22_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_1_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_0_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11241),
            .lcout(frame_decoder_OFF3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_1_22_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_1_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_2_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10978),
            .lcout(frame_decoder_OFF3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_1_22_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_1_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_3_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12529),
            .lcout(frame_decoder_OFF3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_1_22_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_4_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15094),
            .lcout(frame_decoder_OFF3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_1_22_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_5_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11085),
            .lcout(frame_decoder_OFF3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_1_22_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_1_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_6_LC_1_22_6  (
            .in0(N__12439),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_1_22_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_7_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11585),
            .lcout(frame_decoder_OFF3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23853),
            .ce(N__11912),
            .sr(N__23367));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_1_23_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_1_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(N__13459),
            .in2(N__13503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_1_23_1 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_1_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(N__10314),
            .in2(N__11934),
            .in3(N__9321),
            .lcout(\scaler_3.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_0 ),
            .carryout(\scaler_3.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_1_23_2 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_1_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__10308),
            .in2(N__9318),
            .in3(N__9309),
            .lcout(\scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_1 ),
            .carryout(\scaler_3.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_1_23_3 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_1_23_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_1_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(N__10302),
            .in2(N__9378),
            .in3(N__9369),
            .lcout(\scaler_3.un3_source_data_0_cry_2_c_RNIR08I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_2 ),
            .carryout(\scaler_3.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_1_23_4 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_1_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(N__10296),
            .in2(N__9366),
            .in3(N__9357),
            .lcout(\scaler_3.un3_source_data_0_cry_3_c_RNIU49I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_3 ),
            .carryout(\scaler_3.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_1_23_5 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_1_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(N__10290),
            .in2(N__9354),
            .in3(N__9345),
            .lcout(\scaler_3.un3_source_data_0_cry_4_c_RNI19AI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_4 ),
            .carryout(\scaler_3.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_1_23_6 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_1_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(N__10284),
            .in2(N__9342),
            .in3(N__9333),
            .lcout(\scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_5 ),
            .carryout(\scaler_3.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_1_23_7 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_1_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(N__10191),
            .in2(_gnd_net_),
            .in3(N__9330),
            .lcout(\scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_6 ),
            .carryout(\scaler_3.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_1_24_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_1_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_1_24_0  (
            .in0(_gnd_net_),
            .in1(N__9468),
            .in2(N__24750),
            .in3(N__9327),
            .lcout(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_1_24_1 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_1_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_1_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9324),
            .lcout(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIQ6GQ_9_LC_1_24_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIQ6GQ_9_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIQ6GQ_9_LC_1_24_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNIQ6GQ_9_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(N__13289),
            .in2(_gnd_net_),
            .in3(N__23501),
            .lcout(\uart_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIOK9H_4_LC_1_24_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIOK9H_4_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIOK9H_4_LC_1_24_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIOK9H_4_LC_1_24_3  (
            .in0(N__10020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13118),
            .lcout(\uart_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_1_24_4 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_1_24_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(N__9707),
            .in2(_gnd_net_),
            .in3(N__11498),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_1_24_5 .C_ON=1'b0;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_1_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_1_24_5  (
            .in0(N__11682),
            .in1(N__13504),
            .in2(_gnd_net_),
            .in3(N__13460),
            .lcout(\scaler_3.un2_source_data_0_cry_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.N_795_i_l_ofx_LC_1_24_7 .C_ON=1'b0;
    defparam \scaler_3.N_795_i_l_ofx_LC_1_24_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.N_795_i_l_ofx_LC_1_24_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_3.N_795_i_l_ofx_LC_1_24_7  (
            .in0(_gnd_net_),
            .in1(N__10206),
            .in2(_gnd_net_),
            .in3(N__10278),
            .lcout(\scaler_3.N_795_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_1_25_0 .C_ON=1'b1;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_1_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_LC_1_25_0  (
            .in0(_gnd_net_),
            .in1(N__11683),
            .in2(N__9462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.source_data_1_esr_6_LC_1_25_1 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_6_LC_1_25_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_6_LC_1_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_6_LC_1_25_1  (
            .in0(_gnd_net_),
            .in1(N__9446),
            .in2(N__11690),
            .in3(N__9453),
            .lcout(scaler_3_data_6),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_1 ),
            .carryout(\scaler_3.un2_source_data_0_cry_2 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_7_LC_1_25_2 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_7_LC_1_25_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_7_LC_1_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_7_LC_1_25_2  (
            .in0(_gnd_net_),
            .in1(N__9428),
            .in2(N__9450),
            .in3(N__9435),
            .lcout(scaler_3_data_7),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_2 ),
            .carryout(\scaler_3.un2_source_data_0_cry_3 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_8_LC_1_25_3 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_8_LC_1_25_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_8_LC_1_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_8_LC_1_25_3  (
            .in0(_gnd_net_),
            .in1(N__9410),
            .in2(N__9432),
            .in3(N__9417),
            .lcout(scaler_3_data_8),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_3 ),
            .carryout(\scaler_3.un2_source_data_0_cry_4 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_9_LC_1_25_4 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_9_LC_1_25_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_9_LC_1_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_9_LC_1_25_4  (
            .in0(_gnd_net_),
            .in1(N__9392),
            .in2(N__9414),
            .in3(N__9399),
            .lcout(scaler_3_data_9),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_4 ),
            .carryout(\scaler_3.un2_source_data_0_cry_5 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_10_LC_1_25_5 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_10_LC_1_25_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_10_LC_1_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_10_LC_1_25_5  (
            .in0(_gnd_net_),
            .in1(N__9533),
            .in2(N__9396),
            .in3(N__9381),
            .lcout(scaler_3_data_10),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_5 ),
            .carryout(\scaler_3.un2_source_data_0_cry_6 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_11_LC_1_25_6 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_11_LC_1_25_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_11_LC_1_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_11_LC_1_25_6  (
            .in0(_gnd_net_),
            .in1(N__9515),
            .in2(N__9537),
            .in3(N__9522),
            .lcout(scaler_3_data_11),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_6 ),
            .carryout(\scaler_3.un2_source_data_0_cry_7 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_12_LC_1_25_7 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_12_LC_1_25_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_12_LC_1_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_12_LC_1_25_7  (
            .in0(_gnd_net_),
            .in1(N__9497),
            .in2(N__9519),
            .in3(N__9504),
            .lcout(scaler_3_data_12),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_7 ),
            .carryout(\scaler_3.un2_source_data_0_cry_8 ),
            .clk(N__23843),
            .ce(N__11965),
            .sr(N__23388));
    defparam \scaler_3.source_data_1_esr_13_LC_1_26_0 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_13_LC_1_26_0 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_13_LC_1_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_13_LC_1_26_0  (
            .in0(_gnd_net_),
            .in1(N__9501),
            .in2(N__9486),
            .in3(N__9474),
            .lcout(scaler_3_data_13),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_9 ),
            .clk(N__23837),
            .ce(N__11964),
            .sr(N__23394));
    defparam \scaler_3.source_data_1_esr_14_LC_1_26_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_14_LC_1_26_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_14_LC_1_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_3.source_data_1_esr_14_LC_1_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9471),
            .lcout(scaler_3_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23837),
            .ce(N__11964),
            .sr(N__23394));
    defparam \scaler_4.source_data_1_esr_5_LC_1_26_5 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_1_26_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_1_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_1_26_5  (
            .in0(N__10440),
            .in1(N__10474),
            .in2(_gnd_net_),
            .in3(N__10512),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23837),
            .ce(N__11964),
            .sr(N__23394));
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_1_27_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_1_27_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_1_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_0_LC_1_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11252),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_1_27_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_1_27_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_1_27_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_1_LC_1_27_1  (
            .in0(N__12786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_1_27_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_1_27_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_1_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_2_LC_1_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10985),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_1_27_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_1_27_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_1_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_3_LC_1_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12545),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_1_27_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_1_27_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_1_27_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_4_LC_1_27_4  (
            .in0(N__15107),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_1_27_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_1_27_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_1_27_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_5_LC_1_27_5  (
            .in0(N__11093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_1_27_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_1_27_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_1_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_6_LC_1_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12456),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_1_27_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_1_27_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_1_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_7_LC_1_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11586),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23832),
            .ce(N__9549),
            .sr(N__23398));
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_1_28_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_1_28_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_1_28_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_0_LC_1_28_0  (
            .in0(N__11253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_1_28_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_1_28_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_1_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_2_LC_1_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10986),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_1_28_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_1_28_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_1_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_3_LC_1_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12546),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_1_28_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_1_28_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_1_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_4_LC_1_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15108),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_1_28_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_1_28_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_1_28_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_5_LC_1_28_4  (
            .in0(N__11094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_1_28_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_1_28_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_1_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_6_LC_1_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12457),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_1_28_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_1_28_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_1_28_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_1_LC_1_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12787),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23828),
            .ce(N__11484),
            .sr(N__23402));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_1_29_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_1_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_1_29_0  (
            .in0(_gnd_net_),
            .in1(N__10503),
            .in2(N__10482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_1_29_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_1_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_1_29_1  (
            .in0(_gnd_net_),
            .in1(N__9675),
            .in2(N__9669),
            .in3(N__9657),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_1_29_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_1_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_1_29_2  (
            .in0(_gnd_net_),
            .in1(N__9654),
            .in2(N__9648),
            .in3(N__9636),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_1_29_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_1_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_1_29_3  (
            .in0(_gnd_net_),
            .in1(N__9633),
            .in2(N__9627),
            .in3(N__9615),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_1_29_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_1_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_1_29_4  (
            .in0(_gnd_net_),
            .in1(N__9612),
            .in2(N__9606),
            .in3(N__9594),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNI15MI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_1_29_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_1_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_1_29_5  (
            .in0(_gnd_net_),
            .in1(N__9591),
            .in2(N__9582),
            .in3(N__9573),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNI49NI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_1_29_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_1_29_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_1_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_1_29_6  (
            .in0(_gnd_net_),
            .in1(N__9570),
            .in2(N__9564),
            .in3(N__9552),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_1_29_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_1_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_1_29_7  (
            .in0(_gnd_net_),
            .in1(N__9729),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_1_30_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_1_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(N__9693),
            .in2(N__24768),
            .in3(N__9714),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_1_30_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_1_30_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_1_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9711),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_807_i_l_ofx_LC_1_30_7 .C_ON=1'b0;
    defparam \scaler_4.N_807_i_l_ofx_LC_1_30_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_807_i_l_ofx_LC_1_30_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \scaler_4.N_807_i_l_ofx_LC_1_30_7  (
            .in0(N__9708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11505),
            .lcout(\scaler_4.N_807_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_0_LC_2_15_0 .C_ON=1'b0;
    defparam \uart.bit_Count_0_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_0_LC_2_15_0 .LUT_INIT=16'b0010001011001100;
    LogicCell40 \uart.bit_Count_0_LC_2_15_0  (
            .in0(N__10693),
            .in1(N__12876),
            .in2(_gnd_net_),
            .in3(N__12040),
            .lcout(\uart.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23878),
            .ce(),
            .sr(N__23341));
    defparam \uart.bit_Count_2_LC_2_15_2 .C_ON=1'b0;
    defparam \uart.bit_Count_2_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_2_LC_2_15_2 .LUT_INIT=16'b0101000110100010;
    LogicCell40 \uart.bit_Count_2_LC_2_15_2  (
            .in0(N__12985),
            .in1(N__12042),
            .in2(N__10701),
            .in3(N__10707),
            .lcout(\uart.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23878),
            .ce(),
            .sr(N__23341));
    defparam \uart.bit_Count_1_LC_2_15_4 .C_ON=1'b0;
    defparam \uart.bit_Count_1_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_1_LC_2_15_4 .LUT_INIT=16'b0110000010101010;
    LogicCell40 \uart.bit_Count_1_LC_2_15_4  (
            .in0(N__12929),
            .in1(N__12877),
            .in2(N__10700),
            .in3(N__12041),
            .lcout(\uart.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23878),
            .ce(),
            .sr(N__23341));
    defparam \uart.state_RNO_1_3_LC_2_16_0 .C_ON=1'b0;
    defparam \uart.state_RNO_1_3_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_3_LC_2_16_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uart.state_RNO_1_3_LC_2_16_0  (
            .in0(N__10671),
            .in1(N__12277),
            .in2(_gnd_net_),
            .in3(N__24486),
            .lcout(\uart.state_srsts_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_1_LC_2_16_6 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_1_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_1_LC_2_16_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart.data_Aux_RNO_0_1_LC_2_16_6  (
            .in0(N__12981),
            .in1(N__12923),
            .in2(_gnd_net_),
            .in3(N__12862),
            .lcout(\uart.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIDK7E_8_LC_2_17_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIDK7E_8_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIDK7E_8_LC_2_17_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_frame_decoder.WDT_RNIDK7E_8_LC_2_17_0  (
            .in0(N__9895),
            .in1(N__9937),
            .in2(_gnd_net_),
            .in3(N__9686),
            .lcout(\uart_frame_decoder.WDT8lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_2_17_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_2_17_1 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \uart_frame_decoder.WDT_RNIAGPB_10_LC_2_17_1  (
            .in0(N__9938),
            .in1(N__9923),
            .in2(N__9912),
            .in3(N__9896),
            .lcout(),
            .ltout(\uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIM8N32_9_LC_2_17_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIM8N32_9_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIM8N32_9_LC_2_17_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \uart_frame_decoder.WDT_RNIM8N32_9_LC_2_17_2  (
            .in0(N__9881),
            .in1(N__9792),
            .in2(N__9870),
            .in3(N__9867),
            .lcout(\uart_frame_decoder.WDT8lt14_0 ),
            .ltout(\uart_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_2_17_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_2_17_3 .LUT_INIT=16'b0011001100111111;
    LogicCell40 \uart_frame_decoder.WDT_RNI17K92_15_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__9784),
            .in2(N__9861),
            .in3(N__9763),
            .lcout(\uart_frame_decoder.WDT8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIM6B11_4_LC_2_17_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIM6B11_4_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIM6B11_4_LC_2_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_frame_decoder.WDT_RNIM6B11_4_LC_2_17_4  (
            .in0(N__9842),
            .in1(N__9830),
            .in2(N__9819),
            .in3(N__9803),
            .lcout(\uart_frame_decoder.WDT_RNIM6B11Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIJUEI2_15_LC_2_17_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIJUEI2_15_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIJUEI2_15_LC_2_17_5 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \uart_frame_decoder.WDT_RNIJUEI2_15_LC_2_17_5  (
            .in0(N__9785),
            .in1(N__13062),
            .in2(N__9768),
            .in3(N__9747),
            .lcout(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15 ),
            .ltout(\uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_3_LC_2_17_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_3_LC_2_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_3_LC_2_17_6 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \uart_frame_decoder.state_1_3_LC_2_17_6  (
            .in0(N__10118),
            .in1(_gnd_net_),
            .in2(N__9741),
            .in3(N__9738),
            .lcout(\uart_frame_decoder.state_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23872),
            .ce(),
            .sr(N__23343));
    defparam \uart_frame_decoder.state_1_RNINJ9H_3_LC_2_17_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNINJ9H_3_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNINJ9H_3_LC_2_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNINJ9H_3_LC_2_17_7  (
            .in0(N__9737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13061),
            .lcout(\uart_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_1_LC_2_18_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_1_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_1_LC_2_18_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_1_LC_2_18_1  (
            .in0(N__10779),
            .in1(N__12704),
            .in2(N__11165),
            .in3(N__13234),
            .lcout(\uart_frame_decoder.state_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23867),
            .ce(),
            .sr(N__23345));
    defparam \uart_frame_decoder.state_1_2_LC_2_18_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_2_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_2_LC_2_18_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_2_LC_2_18_4  (
            .in0(N__13235),
            .in1(N__10032),
            .in2(N__12708),
            .in3(N__11127),
            .lcout(\uart_frame_decoder.state_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23867),
            .ce(),
            .sr(N__23345));
    defparam \uart_frame_decoder.state_1_RNIMI9H_2_LC_2_18_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIMI9H_2_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIMI9H_2_LC_2_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIMI9H_2_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__10031),
            .in2(_gnd_net_),
            .in3(N__13089),
            .lcout(\uart_frame_decoder.source_CH1data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_4_LC_2_18_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_4_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_4_LC_2_18_7 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uart_frame_decoder.state_1_4_LC_2_18_7  (
            .in0(N__10235),
            .in1(N__10016),
            .in2(_gnd_net_),
            .in3(N__13236),
            .lcout(\uart_frame_decoder.state_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23867),
            .ce(),
            .sr(N__23345));
    defparam \uart_frame_decoder.count_RNIM2UL1_2_LC_2_19_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNIM2UL1_2_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNIM2UL1_2_LC_2_19_0 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \uart_frame_decoder.count_RNIM2UL1_2_LC_2_19_0  (
            .in0(N__10001),
            .in1(N__9984),
            .in2(N__9966),
            .in3(N__10856),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_o2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_2_19_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_2_19_4 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_1_0_LC_2_19_4  (
            .in0(N__11123),
            .in1(N__12698),
            .in2(N__10833),
            .in3(N__10845),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_i_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_0_LC_2_19_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_0_LC_2_19_5 .SEQ_MODE=4'b1001;
    defparam \uart_frame_decoder.state_1_0_LC_2_19_5 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \uart_frame_decoder.state_1_0_LC_2_19_5  (
            .in0(N__10839),
            .in1(N__13301),
            .in2(N__9942),
            .in3(N__13246),
            .lcout(\uart_frame_decoder.state_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23863),
            .ce(),
            .sr(N__23348));
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_2_20_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_2_20_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_2_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_0_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11213),
            .lcout(frame_decoder_OFF2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_2_20_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_2_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_1_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12741),
            .lcout(frame_decoder_OFF2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_2_20_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_2_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_2_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10945),
            .lcout(frame_decoder_OFF2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_2_20_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_2_20_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_3_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__12509),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_2_20_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_2_20_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_2_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_4_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15073),
            .lcout(frame_decoder_OFF2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_2_20_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_2_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_5_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11047),
            .lcout(frame_decoder_OFF2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_2_20_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_2_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_6_LC_2_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12417),
            .lcout(frame_decoder_OFF2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_2_20_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_2_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_7_LC_2_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11553),
            .lcout(frame_decoder_OFF2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23858),
            .ce(N__10104),
            .sr(N__23352));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_21_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(N__15174),
            .in2(N__15222),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_2_21_1 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_2_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(N__10095),
            .in2(N__10089),
            .in3(N__10080),
            .lcout(\scaler_2.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_0 ),
            .carryout(\scaler_2.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_2_21_2 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_2_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(N__10077),
            .in2(N__10071),
            .in3(N__10059),
            .lcout(\scaler_2.un3_source_data_0_cry_1_c_RNILSPH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_1 ),
            .carryout(\scaler_2.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_2_21_3 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_2_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(N__10056),
            .in2(N__10050),
            .in3(N__10041),
            .lcout(\scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_2 ),
            .carryout(\scaler_2.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_2_21_4 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_2_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_2_21_4  (
            .in0(_gnd_net_),
            .in1(N__10038),
            .in2(N__10182),
            .in3(N__10173),
            .lcout(\scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_3 ),
            .carryout(\scaler_2.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_2_21_5 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_2_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(N__10170),
            .in2(N__10164),
            .in3(N__10155),
            .lcout(\scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_4 ),
            .carryout(\scaler_2.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_2_21_6 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_2_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__10152),
            .in2(N__10146),
            .in3(N__10137),
            .lcout(\scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_5 ),
            .carryout(\scaler_2.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_2_21_7 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_2_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(N__10125),
            .in2(_gnd_net_),
            .in3(N__10134),
            .lcout(\scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_6 ),
            .carryout(\scaler_2.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_2_22_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_2_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__10242),
            .in2(N__24749),
            .in3(N__10131),
            .lcout(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_22_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10128),
            .lcout(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_2_22_2 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_2_22_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(N__10253),
            .in2(_gnd_net_),
            .in3(N__10265),
            .lcout(\scaler_2.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIJVFQ_2_LC_2_22_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIJVFQ_2_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIJVFQ_2_LC_2_22_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_RNIJVFQ_2_LC_2_22_4  (
            .in0(N__10119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23498),
            .lcout(\uart_frame_decoder.source_CH1data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIO4GQ_7_LC_2_22_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIO4GQ_7_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIO4GQ_7_LC_2_22_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_RNIO4GQ_7_LC_2_22_5  (
            .in0(N__23499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11654),
            .lcout(\uart_frame_decoder.source_offset2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_2_22_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_2_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_2_22_6  (
            .in0(N__11220),
            .in1(N__11554),
            .in2(N__11081),
            .in3(N__10953),
            .lcout(\uart_frame_decoder.N_79_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.N_783_i_l_ofx_LC_2_22_7 .C_ON=1'b0;
    defparam \scaler_2.N_783_i_l_ofx_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.N_783_i_l_ofx_LC_2_22_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \scaler_2.N_783_i_l_ofx_LC_2_22_7  (
            .in0(N__10266),
            .in1(_gnd_net_),
            .in2(N__10257),
            .in3(_gnd_net_),
            .lcout(\scaler_2.N_783_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIK0GQ_3_LC_2_23_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIK0GQ_3_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIK0GQ_3_LC_2_23_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNIK0GQ_3_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__10236),
            .in2(_gnd_net_),
            .in3(N__23495),
            .lcout(\uart_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIPL9H_5_LC_2_23_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIPL9H_5_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIPL9H_5_LC_2_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIPL9H_5_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__11603),
            .in2(_gnd_net_),
            .in3(N__13110),
            .lcout(\uart_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIM2GQ_5_LC_2_23_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIM2GQ_5_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIM2GQ_5_LC_2_23_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_frame_decoder.state_1_RNIM2GQ_5_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10209),
            .in3(N__23493),
            .lcout(\uart_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_2_23_4 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_2_23_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(N__10202),
            .in2(_gnd_net_),
            .in3(N__10277),
            .lcout(\scaler_3.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNISO9H_8_LC_2_23_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNISO9H_8_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNISO9H_8_LC_2_23_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uart_frame_decoder.state_1_RNISO9H_8_LC_2_23_6  (
            .in0(N__13111),
            .in1(_gnd_net_),
            .in2(N__11637),
            .in3(_gnd_net_),
            .lcout(\uart_frame_decoder.source_offset3data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIP5GQ_8_LC_2_23_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIP5GQ_8_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIP5GQ_8_LC_2_23_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_frame_decoder.state_1_RNIP5GQ_8_LC_2_23_7  (
            .in0(N__23494),
            .in1(_gnd_net_),
            .in2(N__10185),
            .in3(_gnd_net_),
            .lcout(\uart_frame_decoder.source_offset3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_2_24_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_2_24_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_2_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_0_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11242),
            .lcout(frame_decoder_CH3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_2_24_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_2_24_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_2_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_1_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12778),
            .lcout(frame_decoder_CH3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_2_24_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_2_24_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_2_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_2_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10974),
            .lcout(frame_decoder_CH3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_2_24_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_2_24_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_2_24_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_3_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__12530),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_2_24_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_2_24_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_2_24_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_4_LC_2_24_4  (
            .in0(N__15095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_2_24_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_2_24_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_2_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_5_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11086),
            .lcout(frame_decoder_CH3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_2_24_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_2_24_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_2_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_6_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12455),
            .lcout(frame_decoder_CH3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_2_24_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_2_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_7_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11580),
            .lcout(frame_decoder_CH3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23844),
            .ce(N__11445),
            .sr(N__23374));
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_2_25_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_2_25_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_2_25_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_0_LC_2_25_0  (
            .in0(N__11243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH1data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_2_25_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_2_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_2_LC_2_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10975),
            .lcout(frame_decoder_CH1data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_2_25_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_2_25_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_2_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_3_LC_2_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12543),
            .lcout(frame_decoder_CH1data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_2_25_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_2_25_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_2_25_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_1_LC_2_25_4  (
            .in0(N__12779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH1data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_2_25_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_2_25_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_2_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_5_LC_2_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11082),
            .lcout(frame_decoder_CH1data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_2_25_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_2_25_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_2_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_6_LC_2_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12458),
            .lcout(frame_decoder_CH1data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_2_25_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_2_25_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_2_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_7_LC_2_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11581),
            .lcout(frame_decoder_CH1data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23838),
            .ce(N__15017),
            .sr(N__23382));
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_2_26_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_2_26_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_2_26_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_0_LC_2_26_0  (
            .in0(N__11244),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF1data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_2_26_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_2_26_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_2_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_1_LC_2_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12788),
            .lcout(frame_decoder_OFF1data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_2_26_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_2_26_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_2_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_2_LC_2_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10976),
            .lcout(frame_decoder_OFF1data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_2_26_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_2_26_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_2_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_3_LC_2_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12544),
            .lcout(frame_decoder_OFF1data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_2_26_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_2_26_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_2_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_4_LC_2_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15106),
            .lcout(frame_decoder_OFF1data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_2_26_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_2_26_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_2_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_5_LC_2_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11083),
            .lcout(frame_decoder_OFF1data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_2_26_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_2_26_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_2_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_6_LC_2_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12459),
            .lcout(frame_decoder_OFF1data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_2_26_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_2_26_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_2_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_7_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11582),
            .lcout(frame_decoder_OFF1data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23833),
            .ce(N__13401),
            .sr(N__23389));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_2_27_0 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_2_27_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_2_27_0  (
            .in0(_gnd_net_),
            .in1(N__11395),
            .in2(N__11434),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(\scaler_1.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_2_27_1 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_2_27_1 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_2_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_2_27_1  (
            .in0(_gnd_net_),
            .in1(N__10410),
            .in2(N__10401),
            .in3(N__10392),
            .lcout(\scaler_1.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_0 ),
            .carryout(\scaler_1.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_2_27_2 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_2_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_2_27_2  (
            .in0(_gnd_net_),
            .in1(N__10389),
            .in2(N__10380),
            .in3(N__10371),
            .lcout(\scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_1 ),
            .carryout(\scaler_1.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_2_27_3 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_2_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_2_27_3  (
            .in0(_gnd_net_),
            .in1(N__10368),
            .in2(N__10359),
            .in3(N__10350),
            .lcout(\scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_2 ),
            .carryout(\scaler_1.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_2_27_4 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_2_27_4 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_2_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_2_27_4  (
            .in0(_gnd_net_),
            .in1(N__15033),
            .in2(N__10347),
            .in3(N__10338),
            .lcout(\scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_3 ),
            .carryout(\scaler_1.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_2_27_5 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_2_27_5 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_2_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_2_27_5  (
            .in0(_gnd_net_),
            .in1(N__10335),
            .in2(N__10326),
            .in3(N__10317),
            .lcout(\scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_4 ),
            .carryout(\scaler_1.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_2_27_6 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_2_27_6 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_2_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_2_27_6  (
            .in0(_gnd_net_),
            .in1(N__10548),
            .in2(N__10542),
            .in3(N__10530),
            .lcout(\scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_5 ),
            .carryout(\scaler_1.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_2_27_7 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_2_27_7 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_2_27_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_2_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11724),
            .in3(N__10527),
            .lcout(\scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_6 ),
            .carryout(\scaler_1.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_2_28_0 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_2_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_2_28_0  (
            .in0(_gnd_net_),
            .in1(N__10518),
            .in2(N__24767),
            .in3(N__10524),
            .lcout(\scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ),
            .ltout(),
            .carryin(bfn_2_28_0_),
            .carryout(\scaler_1.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_2_28_1 .C_ON=1'b0;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_2_28_1 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_2_28_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_2_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10521),
            .lcout(\scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.N_771_i_l_ofx_LC_2_28_3 .C_ON=1'b0;
    defparam \scaler_1.N_771_i_l_ofx_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \scaler_1.N_771_i_l_ofx_LC_2_28_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_1.N_771_i_l_ofx_LC_2_28_3  (
            .in0(_gnd_net_),
            .in1(N__11754),
            .in2(_gnd_net_),
            .in3(N__11739),
            .lcout(\scaler_1.N_771_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_2_28_5 .C_ON=1'b0;
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_2_28_5 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_2_28_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_2_28_5  (
            .in0(N__11435),
            .in1(N__11857),
            .in2(_gnd_net_),
            .in3(N__11402),
            .lcout(\scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_2_28_7 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_2_28_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_2_28_7  (
            .in0(N__10438),
            .in1(N__10504),
            .in2(_gnd_net_),
            .in3(N__10473),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_2_29_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_2_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_2_29_0  (
            .in0(_gnd_net_),
            .in1(N__10431),
            .in2(N__10449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_2_29_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_2_29_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_2_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_2_29_1  (
            .in0(_gnd_net_),
            .in1(N__10661),
            .in2(N__10439),
            .in3(N__10413),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_7_LC_2_29_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_2_29_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_2_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_2_29_2  (
            .in0(_gnd_net_),
            .in1(N__10646),
            .in2(N__10665),
            .in3(N__10653),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_8_LC_2_29_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_2_29_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_2_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_2_29_3  (
            .in0(_gnd_net_),
            .in1(N__10631),
            .in2(N__10650),
            .in3(N__10638),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_9_LC_2_29_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_2_29_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_2_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_2_29_4  (
            .in0(_gnd_net_),
            .in1(N__10616),
            .in2(N__10635),
            .in3(N__10623),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_10_LC_2_29_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_2_29_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_2_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__10601),
            .in2(N__10620),
            .in3(N__10608),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_11_LC_2_29_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_2_29_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_2_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_2_29_6  (
            .in0(_gnd_net_),
            .in1(N__10586),
            .in2(N__10605),
            .in3(N__10593),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_12_LC_2_29_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_2_29_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_2_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_2_29_7  (
            .in0(_gnd_net_),
            .in1(N__10574),
            .in2(N__10590),
            .in3(N__10578),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__23818),
            .ce(N__11961),
            .sr(N__23403));
    defparam \scaler_4.source_data_1_esr_13_LC_2_30_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_2_30_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_2_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_2_30_0  (
            .in0(_gnd_net_),
            .in1(N__10575),
            .in2(N__10563),
            .in3(N__10554),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__23812),
            .ce(N__11959),
            .sr(N__23405));
    defparam \scaler_4.source_data_1_esr_14_LC_2_30_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_2_30_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_2_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_2_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10551),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23812),
            .ce(N__11959),
            .sr(N__23405));
    defparam \uart.bit_Count_RNO_0_2_LC_3_15_1 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_2_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_2_LC_3_15_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.bit_Count_RNO_0_2_LC_3_15_1  (
            .in0(N__12921),
            .in1(N__12860),
            .in2(_gnd_net_),
            .in3(N__12032),
            .lcout(\uart.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNI4ENK_3_LC_3_15_5 .C_ON=1'b0;
    defparam \uart.state_RNI4ENK_3_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNI4ENK_3_LC_3_15_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \uart.state_RNI4ENK_3_LC_3_15_5  (
            .in0(N__12922),
            .in1(N__12861),
            .in2(N__12986),
            .in3(N__12275),
            .lcout(\uart.N_133_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNIETHE_2_LC_3_16_0 .C_ON=1'b0;
    defparam \uart.bit_Count_RNIETHE_2_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNIETHE_2_LC_3_16_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.bit_Count_RNIETHE_2_LC_3_16_0  (
            .in0(N__12973),
            .in1(N__12918),
            .in2(_gnd_net_),
            .in3(N__12855),
            .lcout(\uart.N_177 ),
            .ltout(\uart.N_177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIBAKE2_6_LC_3_16_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIBAKE2_6_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIBAKE2_6_LC_3_16_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uart.timer_Count_RNIBAKE2_6_LC_3_16_1  (
            .in0(N__14248),
            .in1(N__14298),
            .in2(N__10683),
            .in3(N__12021),
            .lcout(\uart.N_168_1 ),
            .ltout(\uart.N_168_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_3_LC_3_16_2 .C_ON=1'b0;
    defparam \uart.state_3_LC_3_16_2 .SEQ_MODE=4'b1000;
    defparam \uart.state_3_LC_3_16_2 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \uart.state_3_LC_3_16_2  (
            .in0(N__12087),
            .in1(N__10680),
            .in2(N__10674),
            .in3(N__12147),
            .lcout(\uart.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23873),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_5_LC_3_16_3 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_5_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_5_LC_3_16_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart.data_Aux_RNO_0_5_LC_3_16_3  (
            .in0(N__12858),
            .in1(N__12976),
            .in2(_gnd_net_),
            .in3(N__12925),
            .lcout(\uart.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_6_LC_3_16_4 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_6_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_6_LC_3_16_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart.data_Aux_RNO_0_6_LC_3_16_4  (
            .in0(N__12977),
            .in1(N__12920),
            .in2(_gnd_net_),
            .in3(N__12859),
            .lcout(\uart.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_0_LC_3_16_5 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_0_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_0_LC_3_16_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart.data_Aux_RNO_0_0_LC_3_16_5  (
            .in0(N__12856),
            .in1(N__12974),
            .in2(_gnd_net_),
            .in3(N__12924),
            .lcout(\uart.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_3_LC_3_16_6 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_3_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_3_LC_3_16_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart.data_Aux_RNO_0_3_LC_3_16_6  (
            .in0(N__12975),
            .in1(N__12919),
            .in2(_gnd_net_),
            .in3(N__12857),
            .lcout(\uart.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_3_3_LC_3_16_7 .C_ON=1'b0;
    defparam \uart.state_RNO_3_3_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_3_3_LC_3_16_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.state_RNO_3_3_LC_3_16_7  (
            .in0(N__12084),
            .in1(N__14247),
            .in2(_gnd_net_),
            .in3(N__14297),
            .lcout(\uart.N_154_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_7_LC_3_17_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_7_LC_3_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_7_LC_3_17_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uart_frame_decoder.state_1_7_LC_3_17_2  (
            .in0(N__13416),
            .in1(N__10823),
            .in2(_gnd_net_),
            .in3(N__13237),
            .lcout(\uart_frame_decoder.state_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23868),
            .ce(),
            .sr(N__23342));
    defparam \uart.data_rdy_LC_3_17_5 .C_ON=1'b0;
    defparam \uart.data_rdy_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_rdy_LC_3_17_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uart.data_rdy_LC_3_17_5  (
            .in0(N__12207),
            .in1(N__14250),
            .in2(N__12638),
            .in3(N__12310),
            .lcout(uart_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23868),
            .ce(),
            .sr(N__23342));
    defparam \uart.data_Aux_0_LC_3_18_0 .C_ON=1'b0;
    defparam \uart.data_Aux_0_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_0_LC_3_18_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart.data_Aux_0_LC_3_18_0  (
            .in0(N__12627),
            .in1(N__10755),
            .in2(N__10772),
            .in3(N__12113),
            .lcout(\uart.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_1_LC_3_18_1 .C_ON=1'b0;
    defparam \uart.data_Aux_1_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_1_LC_3_18_1 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uart.data_Aux_1_LC_3_18_1  (
            .in0(N__12114),
            .in1(N__12630),
            .in2(N__10746),
            .in3(N__10889),
            .lcout(\uart.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_2_LC_3_18_2 .C_ON=1'b0;
    defparam \uart.data_Aux_2_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_2_LC_3_18_2 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart.data_Aux_2_LC_3_18_2  (
            .in0(N__12628),
            .in1(N__12822),
            .in2(N__11003),
            .in3(N__12115),
            .lcout(\uart.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_3_LC_3_18_3 .C_ON=1'b0;
    defparam \uart.data_Aux_3_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_3_LC_3_18_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart.data_Aux_3_LC_3_18_3  (
            .in0(N__12116),
            .in1(N__12631),
            .in2(N__12563),
            .in3(N__10734),
            .lcout(\uart.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_4_LC_3_18_4 .C_ON=1'b0;
    defparam \uart.data_Aux_4_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_4_LC_3_18_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart.data_Aux_4_LC_3_18_4  (
            .in0(N__12629),
            .in1(N__12348),
            .in2(N__13346),
            .in3(N__12117),
            .lcout(\uart.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_5_LC_3_18_5 .C_ON=1'b0;
    defparam \uart.data_Aux_5_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_5_LC_3_18_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart.data_Aux_5_LC_3_18_5  (
            .in0(N__12118),
            .in1(N__12632),
            .in2(N__11111),
            .in3(N__10725),
            .lcout(\uart.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_6_LC_3_18_6 .C_ON=1'b0;
    defparam \uart.data_Aux_6_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_6_LC_3_18_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart.data_Aux_6_LC_3_18_6  (
            .in0(N__10716),
            .in1(N__12470),
            .in2(N__12639),
            .in3(N__12119),
            .lcout(\uart.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.data_Aux_7_LC_3_18_7 .C_ON=1'b0;
    defparam \uart.data_Aux_7_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_7_LC_3_18_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uart.data_Aux_7_LC_3_18_7  (
            .in0(N__12120),
            .in1(N__12633),
            .in2(N__10875),
            .in3(N__10904),
            .lcout(\uart.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23864),
            .ce(),
            .sr(N__12321));
    defparam \uart.state_RNO_0_0_LC_3_19_0 .C_ON=1'b0;
    defparam \uart.state_RNO_0_0_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_0_LC_3_19_0 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart.state_RNO_0_0_LC_3_19_0  (
            .in0(N__12681),
            .in1(N__12626),
            .in2(_gnd_net_),
            .in3(N__23503),
            .lcout(),
            .ltout(\uart.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_0_LC_3_19_1 .C_ON=1'b0;
    defparam \uart.state_0_LC_3_19_1 .SEQ_MODE=4'b1000;
    defparam \uart.state_0_LC_3_19_1 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart.state_0_LC_3_19_1  (
            .in0(N__12208),
            .in1(N__14249),
            .in2(N__10863),
            .in3(N__12312),
            .lcout(\uart.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23859),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI592G_10_LC_3_19_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI592G_10_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI592G_10_LC_3_19_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uart_frame_decoder.state_1_RNI592G_10_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__13156),
            .in2(_gnd_net_),
            .in3(N__13090),
            .lcout(\uart_frame_decoder.state_1_RNI592GZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_3_19_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_3_19_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_3_0_LC_3_19_3  (
            .in0(N__13157),
            .in1(N__11151),
            .in2(_gnd_net_),
            .in3(N__10793),
            .lcout(\uart_frame_decoder.state_1_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_3_19_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_3_19_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_0_LC_3_19_4  (
            .in0(N__10808),
            .in1(_gnd_net_),
            .in2(N__11161),
            .in3(N__13161),
            .lcout(\uart_frame_decoder.N_168_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_3_19_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_3_19_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_2_0_LC_3_19_5  (
            .in0(N__13092),
            .in1(N__11150),
            .in2(N__13168),
            .in3(N__10807),
            .lcout(\uart_frame_decoder.state_1_RNO_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIRN9H_7_LC_3_19_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIRN9H_7_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIRN9H_7_LC_3_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIRN9H_7_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__10824),
            .in2(_gnd_net_),
            .in3(N__13091),
            .lcout(\uart_frame_decoder.source_offset2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_3_19_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_3_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_1_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__10809),
            .in2(_gnd_net_),
            .in3(N__10794),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_0_LC_3_20_0 .C_ON=1'b0;
    defparam \uart.data_0_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_0_LC_3_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart.data_0_LC_3_20_0  (
            .in0(N__11212),
            .in1(N__10773),
            .in2(_gnd_net_),
            .in3(N__13382),
            .lcout(uart_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23854),
            .ce(),
            .sr(N__13329));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_3_20_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_3_20_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__11045),
            .in2(_gnd_net_),
            .in3(N__11211),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI12LB1_1_LC_3_20_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI12LB1_1_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI12LB1_1_LC_3_20_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_frame_decoder.state_1_RNI12LB1_1_LC_3_20_2  (
            .in0(N__11166),
            .in1(N__11544),
            .in2(N__11130),
            .in3(N__10943),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_5_LC_3_20_3 .C_ON=1'b0;
    defparam \uart.data_5_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_5_LC_3_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.data_5_LC_3_20_3  (
            .in0(N__13385),
            .in1(N__11112),
            .in2(_gnd_net_),
            .in3(N__11046),
            .lcout(uart_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23854),
            .ce(),
            .sr(N__13329));
    defparam \uart.data_2_LC_3_20_4 .C_ON=1'b0;
    defparam \uart.data_2_LC_3_20_4 .SEQ_MODE=4'b1000;
    defparam \uart.data_2_LC_3_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart.data_2_LC_3_20_4  (
            .in0(N__11007),
            .in1(N__10944),
            .in2(_gnd_net_),
            .in3(N__13384),
            .lcout(uart_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23854),
            .ce(),
            .sr(N__13329));
    defparam \uart.data_7_LC_3_20_5 .C_ON=1'b0;
    defparam \uart.data_7_LC_3_20_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_7_LC_3_20_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uart.data_7_LC_3_20_5  (
            .in0(N__13386),
            .in1(_gnd_net_),
            .in2(N__11570),
            .in3(N__10908),
            .lcout(uart_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23854),
            .ce(),
            .sr(N__13329));
    defparam \uart.data_1_LC_3_20_6 .C_ON=1'b0;
    defparam \uart.data_1_LC_3_20_6 .SEQ_MODE=4'b1000;
    defparam \uart.data_1_LC_3_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart.data_1_LC_3_20_6  (
            .in0(N__10893),
            .in1(N__12740),
            .in2(_gnd_net_),
            .in3(N__13383),
            .lcout(uart_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23854),
            .ce(),
            .sr(N__13329));
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_3_21_0 .C_ON=1'b1;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_3_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__14598),
            .in2(N__14580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_6_LC_3_21_1 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_6_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_6_LC_3_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_6_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__11366),
            .in2(N__14606),
            .in3(N__10878),
            .lcout(scaler_2_data_6),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_1 ),
            .carryout(\scaler_2.un2_source_data_0_cry_2 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_7_LC_3_21_2 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_7_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_7_LC_3_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_7_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__11351),
            .in2(N__11370),
            .in3(N__11358),
            .lcout(scaler_2_data_7),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_2 ),
            .carryout(\scaler_2.un2_source_data_0_cry_3 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_8_LC_3_21_3 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_8_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_8_LC_3_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_8_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__11336),
            .in2(N__11355),
            .in3(N__11343),
            .lcout(scaler_2_data_8),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_3 ),
            .carryout(\scaler_2.un2_source_data_0_cry_4 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_9_LC_3_21_4 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_9_LC_3_21_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_9_LC_3_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_9_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__11321),
            .in2(N__11340),
            .in3(N__11328),
            .lcout(scaler_2_data_9),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_4 ),
            .carryout(\scaler_2.un2_source_data_0_cry_5 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_10_LC_3_21_5 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_10_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_10_LC_3_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_10_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(N__11306),
            .in2(N__11325),
            .in3(N__11313),
            .lcout(scaler_2_data_10),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_5 ),
            .carryout(\scaler_2.un2_source_data_0_cry_6 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_11_LC_3_21_6 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_11_LC_3_21_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_11_LC_3_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_11_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__11291),
            .in2(N__11310),
            .in3(N__11298),
            .lcout(scaler_2_data_11),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_6 ),
            .carryout(\scaler_2.un2_source_data_0_cry_7 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_12_LC_3_21_7 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_12_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_12_LC_3_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_12_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__11279),
            .in2(N__11295),
            .in3(N__11283),
            .lcout(scaler_2_data_12),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_7 ),
            .carryout(\scaler_2.un2_source_data_0_cry_8 ),
            .clk(N__23850),
            .ce(N__11967),
            .sr(N__23353));
    defparam \scaler_2.source_data_1_esr_13_LC_3_22_0 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_13_LC_3_22_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_13_LC_3_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_13_LC_3_22_0  (
            .in0(_gnd_net_),
            .in1(N__11280),
            .in2(N__11268),
            .in3(N__11259),
            .lcout(scaler_2_data_13),
            .ltout(),
            .carryin(bfn_3_22_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_9 ),
            .clk(N__23848),
            .ce(N__11966),
            .sr(N__23359));
    defparam \scaler_2.source_data_1_esr_14_LC_3_22_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_14_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_14_LC_3_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_2.source_data_1_esr_14_LC_3_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11256),
            .lcout(scaler_2_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23848),
            .ce(N__11966),
            .sr(N__23359));
    defparam \scaler_2.source_data_1_esr_5_LC_3_22_5 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_5_LC_3_22_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_5_LC_3_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.source_data_1_esr_5_LC_3_22_5  (
            .in0(N__15229),
            .in1(N__14602),
            .in2(_gnd_net_),
            .in3(N__15194),
            .lcout(scaler_2_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23848),
            .ce(N__11966),
            .sr(N__23359));
    defparam \scaler_3.source_data_1_esr_5_LC_3_22_7 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_5_LC_3_22_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_5_LC_3_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.source_data_1_esr_5_LC_3_22_7  (
            .in0(N__13505),
            .in1(N__11691),
            .in2(_gnd_net_),
            .in3(N__13473),
            .lcout(scaler_3_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23848),
            .ce(N__11966),
            .sr(N__23359));
    defparam \uart_frame_decoder.state_1_8_LC_3_23_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_8_LC_3_23_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_8_LC_3_23_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uart_frame_decoder.state_1_8_LC_3_23_2  (
            .in0(N__11636),
            .in1(N__11658),
            .in2(_gnd_net_),
            .in3(N__13265),
            .lcout(\uart_frame_decoder.state_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23845),
            .ce(),
            .sr(N__23363));
    defparam \uart_frame_decoder.state_1_9_LC_3_23_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_9_LC_3_23_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_9_LC_3_23_3 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \uart_frame_decoder.state_1_9_LC_3_23_3  (
            .in0(N__13266),
            .in1(_gnd_net_),
            .in2(N__11616),
            .in3(N__11622),
            .lcout(\uart_frame_decoder.state_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23845),
            .ce(),
            .sr(N__23363));
    defparam \uart_frame_decoder.state_1_RNITP9H_9_LC_3_23_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNITP9H_9_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNITP9H_9_LC_3_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNITP9H_9_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(N__11612),
            .in2(_gnd_net_),
            .in3(N__13106),
            .lcout(\uart_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_5_LC_3_23_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_5_LC_3_23_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_5_LC_3_23_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uart_frame_decoder.state_1_5_LC_3_23_6  (
            .in0(N__11604),
            .in1(N__11463),
            .in2(_gnd_net_),
            .in3(N__13263),
            .lcout(\uart_frame_decoder.state_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23845),
            .ce(),
            .sr(N__23363));
    defparam \uart_frame_decoder.state_1_6_LC_3_23_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_6_LC_3_23_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_6_LC_3_23_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uart_frame_decoder.state_1_6_LC_3_23_7  (
            .in0(N__13264),
            .in1(N__11592),
            .in2(_gnd_net_),
            .in3(N__13430),
            .lcout(\uart_frame_decoder.state_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23845),
            .ce(),
            .sr(N__23363));
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_3_24_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_3_24_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_3_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_7_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11583),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23839),
            .ce(N__11477),
            .sr(N__23368));
    defparam \uart_frame_decoder.state_1_RNIL1GQ_4_LC_3_24_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIL1GQ_4_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIL1GQ_4_LC_3_24_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNIL1GQ_4_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__11459),
            .in2(_gnd_net_),
            .in3(N__23502),
            .lcout(\uart_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.source_data_1_esr_5_LC_3_25_0 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_5_LC_3_25_0 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_5_LC_3_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_1.source_data_1_esr_5_LC_3_25_0  (
            .in0(N__11859),
            .in1(N__11430),
            .in2(_gnd_net_),
            .in3(N__11394),
            .lcout(scaler_1_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23834),
            .ce(N__11963),
            .sr(N__23375));
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_3_25_7 .C_ON=1'b0;
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_3_25_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(N__11750),
            .in2(_gnd_net_),
            .in3(N__11735),
            .lcout(\scaler_1.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_3_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_3_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__13526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_3_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_3_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__16613),
            .in2(_gnd_net_),
            .in3(N__11712),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_3_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_3_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__16688),
            .in2(_gnd_net_),
            .in3(N__11709),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_3_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_3_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__15284),
            .in2(_gnd_net_),
            .in3(N__11706),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_3_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_3_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13616),
            .in3(N__11703),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_3_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_3_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_3_26_5  (
            .in0(_gnd_net_),
            .in1(N__13208),
            .in2(_gnd_net_),
            .in3(N__11700),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_3_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_3_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_3_26_6  (
            .in0(_gnd_net_),
            .in1(N__15134),
            .in2(_gnd_net_),
            .in3(N__11697),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_3_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_3_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_3_26_7  (
            .in0(_gnd_net_),
            .in1(N__13559),
            .in2(N__24771),
            .in3(N__11694),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_3_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_3_27_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__11880),
            .in2(_gnd_net_),
            .in3(N__11871),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23823),
            .ce(N__16261),
            .sr(N__23390));
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_3_28_0 .C_ON=1'b1;
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_3_28_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_3_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_1.un2_source_data_0_cry_1_c_LC_3_28_0  (
            .in0(_gnd_net_),
            .in1(N__11850),
            .in2(N__11868),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_28_0_),
            .carryout(\scaler_1.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.source_data_1_esr_6_LC_3_28_1 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_6_LC_3_28_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_6_LC_3_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_6_LC_3_28_1  (
            .in0(_gnd_net_),
            .in1(N__11825),
            .in2(N__11858),
            .in3(N__11832),
            .lcout(scaler_1_data_6),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_1 ),
            .carryout(\scaler_1.un2_source_data_0_cry_2 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_7_LC_3_28_2 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_7_LC_3_28_2 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_7_LC_3_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_7_LC_3_28_2  (
            .in0(_gnd_net_),
            .in1(N__11810),
            .in2(N__11829),
            .in3(N__11817),
            .lcout(scaler_1_data_7),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_2 ),
            .carryout(\scaler_1.un2_source_data_0_cry_3 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_8_LC_3_28_3 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_8_LC_3_28_3 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_8_LC_3_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_8_LC_3_28_3  (
            .in0(_gnd_net_),
            .in1(N__11795),
            .in2(N__11814),
            .in3(N__11802),
            .lcout(scaler_1_data_8),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_3 ),
            .carryout(\scaler_1.un2_source_data_0_cry_4 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_9_LC_3_28_4 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_9_LC_3_28_4 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_9_LC_3_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_9_LC_3_28_4  (
            .in0(_gnd_net_),
            .in1(N__11780),
            .in2(N__11799),
            .in3(N__11787),
            .lcout(scaler_1_data_9),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_4 ),
            .carryout(\scaler_1.un2_source_data_0_cry_5 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_10_LC_3_28_5 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_10_LC_3_28_5 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_10_LC_3_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_10_LC_3_28_5  (
            .in0(_gnd_net_),
            .in1(N__11765),
            .in2(N__11784),
            .in3(N__11772),
            .lcout(scaler_1_data_10),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_5 ),
            .carryout(\scaler_1.un2_source_data_0_cry_6 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_11_LC_3_28_6 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_11_LC_3_28_6 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_11_LC_3_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_11_LC_3_28_6  (
            .in0(_gnd_net_),
            .in1(N__12005),
            .in2(N__11769),
            .in3(N__11757),
            .lcout(scaler_1_data_11),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_6 ),
            .carryout(\scaler_1.un2_source_data_0_cry_7 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_12_LC_3_28_7 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_12_LC_3_28_7 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_12_LC_3_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_12_LC_3_28_7  (
            .in0(_gnd_net_),
            .in1(N__11993),
            .in2(N__12009),
            .in3(N__11997),
            .lcout(scaler_1_data_12),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_7 ),
            .carryout(\scaler_1.un2_source_data_0_cry_8 ),
            .clk(N__23819),
            .ce(N__11962),
            .sr(N__23395));
    defparam \scaler_1.source_data_1_esr_13_LC_3_29_0 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_13_LC_3_29_0 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_13_LC_3_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_13_LC_3_29_0  (
            .in0(_gnd_net_),
            .in1(N__11994),
            .in2(N__11982),
            .in3(N__11973),
            .lcout(scaler_1_data_13),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(\scaler_1.un2_source_data_0_cry_9 ),
            .clk(N__23813),
            .ce(N__11960),
            .sr(N__23399));
    defparam \scaler_1.source_data_1_esr_14_LC_3_29_1 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_14_LC_3_29_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_14_LC_3_29_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_1.source_data_1_esr_14_LC_3_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11970),
            .lcout(scaler_1_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23813),
            .ce(N__11960),
            .sr(N__23399));
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_3_30_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_3_30_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_3_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_1_LC_3_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12792),
            .lcout(frame_decoder_OFF3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23808),
            .ce(N__11916),
            .sr(N__23404));
    defparam \uart_sync.aux_2__0__0_LC_4_9_2 .C_ON=1'b0;
    defparam \uart_sync.aux_2__0__0_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_2__0__0_LC_4_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_2__0__0_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13980),
            .lcout(\uart_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23881),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.aux_3__0__0_LC_4_10_0 .C_ON=1'b0;
    defparam \uart_sync.aux_3__0__0_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_3__0__0_LC_4_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_3__0__0_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11895),
            .lcout(\uart_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23880),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_1_LC_4_13_3 .C_ON=1'b0;
    defparam \uart.timer_Count_1_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_1_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.timer_Count_1_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__14143),
            .in2(_gnd_net_),
            .in3(N__13972),
            .lcout(\uart.timer_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23879),
            .ce(),
            .sr(N__14183));
    defparam \uart.state_RNO_0_2_LC_4_14_3 .C_ON=1'b0;
    defparam \uart.state_RNO_0_2_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_2_LC_4_14_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \uart.state_RNO_0_2_LC_4_14_3  (
            .in0(N__12595),
            .in1(N__12659),
            .in2(_gnd_net_),
            .in3(N__12086),
            .lcout(\uart.N_151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.Q_0__0_LC_4_14_6 .C_ON=1'b0;
    defparam \uart_sync.Q_0__0_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_sync.Q_0__0_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.Q_0__0_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11889),
            .lcout(uart_input_sync),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIB0BC_2_LC_4_15_0 .C_ON=1'b0;
    defparam \uart.state_RNIB0BC_2_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIB0BC_2_LC_4_15_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.state_RNIB0BC_2_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__12085),
            .in2(_gnd_net_),
            .in3(N__12273),
            .lcout(\uart.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_2_LC_4_15_1 .C_ON=1'b0;
    defparam \uart.state_2_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \uart.state_2_LC_4_15_1 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \uart.state_2_LC_4_15_1  (
            .in0(N__12093),
            .in1(N__12054),
            .in2(N__12666),
            .in3(N__24463),
            .lcout(\uart.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23874),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIGITG2_0_4_LC_4_15_2 .C_ON=1'b0;
    defparam \uart.state_RNIGITG2_0_4_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIGITG2_0_4_LC_4_15_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uart.state_RNIGITG2_0_4_LC_4_15_2  (
            .in0(N__14218),
            .in1(_gnd_net_),
            .in2(N__12216),
            .in3(N__12309),
            .lcout(),
            .ltout(\uart.timer_Count_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNILCH65_2_LC_4_15_3 .C_ON=1'b0;
    defparam \uart.state_RNILCH65_2_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNILCH65_2_LC_4_15_3 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \uart.state_RNILCH65_2_LC_4_15_3  (
            .in0(N__12063),
            .in1(N__12053),
            .in2(N__12057),
            .in3(N__24462),
            .lcout(\uart.timer_Count_1_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNITC202_6_LC_4_15_4 .C_ON=1'b0;
    defparam \uart.timer_Count_RNITC202_6_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNITC202_6_LC_4_15_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart.timer_Count_RNITC202_6_LC_4_15_4  (
            .in0(N__14217),
            .in1(N__14279),
            .in2(_gnd_net_),
            .in3(N__12020),
            .lcout(\uart.N_180 ),
            .ltout(\uart.N_180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIAFDC2_3_LC_4_15_5 .C_ON=1'b0;
    defparam \uart.state_RNIAFDC2_3_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIAFDC2_3_LC_4_15_5 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \uart.state_RNIAFDC2_3_LC_4_15_5  (
            .in0(N__12272),
            .in1(_gnd_net_),
            .in2(N__12045),
            .in3(N__12209),
            .lcout(\uart.un1_state_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNINU001_1_LC_4_15_6 .C_ON=1'b0;
    defparam \uart.timer_Count_RNINU001_1_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNINU001_1_LC_4_15_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart.timer_Count_RNINU001_1_LC_4_15_6  (
            .in0(N__13948),
            .in1(_gnd_net_),
            .in2(N__13926),
            .in3(N__13973),
            .lcout(\uart.N_146_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIQPMA1_2_LC_4_15_7 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIQPMA1_2_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIQPMA1_2_LC_4_15_7 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uart.timer_Count_RNIQPMA1_2_LC_4_15_7  (
            .in0(N__14114),
            .in1(N__13920),
            .in2(N__14328),
            .in3(N__13947),
            .lcout(\uart.N_143_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_4_16_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__14081),
            .in2(_gnd_net_),
            .in3(N__14056),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_4_16_1 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_4_16_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_4_16_1  (
            .in0(N__12365),
            .in1(N__14647),
            .in2(N__12156),
            .in3(N__12342),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23869),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIICSG1_5_LC_4_16_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIICSG1_5_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIICSG1_5_LC_4_16_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uart.timer_Count_RNIICSG1_5_LC_4_16_2  (
            .in0(N__14326),
            .in1(N__12213),
            .in2(N__14291),
            .in3(N__14091),
            .lcout(\uart.un1_state_2_0_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_4_16_3 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_4_16_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_4_16_3  (
            .in0(N__12364),
            .in1(N__14646),
            .in2(_gnd_net_),
            .in3(N__12341),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23869),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIN6202_4_LC_4_16_4 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIN6202_4_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIN6202_4_LC_4_16_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uart.timer_Count_RNIN6202_4_LC_4_16_4  (
            .in0(N__14324),
            .in1(N__12131),
            .in2(N__14290),
            .in3(N__14115),
            .lcout(\uart.N_153_0 ),
            .ltout(\uart.N_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_4_LC_4_16_5 .C_ON=1'b0;
    defparam \uart.state_RNO_0_4_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_4_LC_4_16_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart.state_RNO_0_4_LC_4_16_5  (
            .in0(N__12214),
            .in1(N__24467),
            .in2(N__12153),
            .in3(N__14227),
            .lcout(\uart.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_2_3_LC_4_16_6 .C_ON=1'b0;
    defparam \uart.state_RNO_2_3_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_2_3_LC_4_16_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart.state_RNO_2_3_LC_4_16_6  (
            .in0(N__14325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12274),
            .lcout(),
            .ltout(\uart.state_srsts_i_a3_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_3_LC_4_16_7 .C_ON=1'b0;
    defparam \uart.state_RNO_0_3_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_3_LC_4_16_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \uart.state_RNO_0_3_LC_4_16_7  (
            .in0(N__14116),
            .in1(N__13925),
            .in2(N__12150),
            .in3(N__13950),
            .lcout(\uart.N_170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIMD8T2_3_LC_4_17_0 .C_ON=1'b0;
    defparam \uart.state_RNIMD8T2_3_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIMD8T2_3_LC_4_17_0 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart.state_RNIMD8T2_3_LC_4_17_0  (
            .in0(N__12276),
            .in1(N__12141),
            .in2(N__12215),
            .in3(N__12135),
            .lcout(\uart.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_4_17_1 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_4_17_1 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \reset_module_System.count_2_LC_4_17_1  (
            .in0(N__14022),
            .in1(N__12340),
            .in2(N__14652),
            .in3(N__12366),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23865),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_4_17_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_4_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_4_17_2  (
            .in0(N__14408),
            .in1(N__14423),
            .in2(N__14394),
            .in3(N__14453),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_4_17_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_4_17_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_4_17_3  (
            .in0(N__14012),
            .in1(N__14438),
            .in2(N__14490),
            .in3(N__14033),
            .lcout(),
            .ltout(\reset_module_System.reset6_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_12_LC_4_17_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_4_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_12_LC_4_17_4  (
            .in0(N__14346),
            .in1(N__14080),
            .in2(N__12369),
            .in3(N__12801),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_4_17_5 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_4_17_5 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \reset_module_System.count_0_LC_4_17_5  (
            .in0(N__14648),
            .in1(N__14085),
            .in2(N__12351),
            .in3(N__12339),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23865),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIP8RT_10_LC_4_18_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_4_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_4_18_0  (
            .in0(N__14375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_4_LC_4_18_1 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_4_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_4_LC_4_18_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart.data_Aux_RNO_0_4_LC_4_18_1  (
            .in0(N__12879),
            .in1(_gnd_net_),
            .in2(N__12939),
            .in3(N__12993),
            .lcout(\uart.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_4_18_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_4_18_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_4_18_2  (
            .in0(N__14469),
            .in1(N__14547),
            .in2(N__14514),
            .in3(N__14058),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIAFHL_3_LC_4_18_3 .C_ON=1'b0;
    defparam \uart.state_RNIAFHL_3_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIAFHL_3_LC_4_18_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart.state_RNIAFHL_3_LC_4_18_3  (
            .in0(N__12206),
            .in1(N__12284),
            .in2(_gnd_net_),
            .in3(N__23500),
            .lcout(\uart.state_RNIAFHLZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIGITG2_4_LC_4_18_4 .C_ON=1'b0;
    defparam \uart.state_RNIGITG2_4_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIGITG2_4_LC_4_18_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \uart.state_RNIGITG2_4_LC_4_18_4  (
            .in0(N__12202),
            .in1(N__14240),
            .in2(_gnd_net_),
            .in3(N__12311),
            .lcout(\uart.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_4_LC_4_18_5 .C_ON=1'b0;
    defparam \uart.state_4_LC_4_18_5 .SEQ_MODE=4'b1000;
    defparam \uart.state_4_LC_4_18_5 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \uart.state_4_LC_4_18_5  (
            .in0(N__12285),
            .in1(N__24487),
            .in2(N__12237),
            .in3(N__12225),
            .lcout(\uart.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23860),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_2_LC_4_18_6 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_2_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_2_LC_4_18_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart.data_Aux_RNO_0_2_LC_4_18_6  (
            .in0(N__12992),
            .in1(N__12935),
            .in2(_gnd_net_),
            .in3(N__12878),
            .lcout(\uart.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI53692_14_LC_4_19_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI53692_14_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI53692_14_LC_4_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI53692_14_LC_4_19_0  (
            .in0(N__14564),
            .in1(N__12816),
            .in2(N__14532),
            .in3(N__12807),
            .lcout(\reset_module_System.reset6_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_4_19_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_4_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_4_19_2  (
            .in0(N__12495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12397),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_4_19_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_4_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_4_19_3  (
            .in0(N__15056),
            .in1(N__12739),
            .in2(N__12711),
            .in3(N__13099),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_1_LC_4_19_6 .C_ON=1'b0;
    defparam \uart.state_1_LC_4_19_6 .SEQ_MODE=4'b1000;
    defparam \uart.state_1_LC_4_19_6 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart.state_1_LC_4_19_6  (
            .in0(N__12680),
            .in1(N__12658),
            .in2(N__12637),
            .in3(N__23530),
            .lcout(\uart.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23855),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIQABT2_4_LC_4_19_7 .C_ON=1'b0;
    defparam \uart.state_RNIQABT2_4_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIQABT2_4_LC_4_19_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \uart.state_RNIQABT2_4_LC_4_19_7  (
            .in0(N__12599),
            .in1(N__24500),
            .in2(_gnd_net_),
            .in3(N__13360),
            .lcout(\uart.state_RNIQABT2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_3_LC_4_20_0 .C_ON=1'b0;
    defparam \uart.data_3_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_3_LC_4_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart.data_3_LC_4_20_0  (
            .in0(N__12564),
            .in1(N__12496),
            .in2(_gnd_net_),
            .in3(N__13379),
            .lcout(uart_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23851),
            .ce(),
            .sr(N__13325));
    defparam \uart.data_6_LC_4_20_2 .C_ON=1'b0;
    defparam \uart.data_6_LC_4_20_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_6_LC_4_20_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart.data_6_LC_4_20_2  (
            .in0(N__12477),
            .in1(N__12398),
            .in2(_gnd_net_),
            .in3(N__13381),
            .lcout(uart_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23851),
            .ce(),
            .sr(N__13325));
    defparam \uart_frame_decoder.state_1_RNIQM9H_6_LC_4_20_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIQM9H_6_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIQM9H_6_LC_4_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIQM9H_6_LC_4_20_3  (
            .in0(N__13434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13093),
            .lcout(\uart_frame_decoder.source_offset1data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIN3GQ_6_LC_4_20_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIN3GQ_6_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIN3GQ_6_LC_4_20_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_frame_decoder.state_1_RNIN3GQ_6_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13404),
            .in3(N__23497),
            .lcout(\uart_frame_decoder.source_offset1data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_4_LC_4_20_5 .C_ON=1'b0;
    defparam \uart.data_4_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_4_LC_4_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uart.data_4_LC_4_20_5  (
            .in0(N__13380),
            .in1(N__13347),
            .in2(_gnd_net_),
            .in3(N__15057),
            .lcout(uart_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23851),
            .ce(),
            .sr(N__13325));
    defparam \scaler_1.source_data_valid_LC_4_21_1 .C_ON=1'b0;
    defparam \scaler_1.source_data_valid_LC_4_21_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_valid_LC_4_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \scaler_1.source_data_valid_LC_4_21_1  (
            .in0(N__14916),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(scaler_1_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23849),
            .ce(),
            .sr(N__23349));
    defparam \uart_frame_decoder.state_1_10_LC_4_21_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_10_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_10_LC_4_21_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \uart_frame_decoder.state_1_10_LC_4_21_2  (
            .in0(N__13154),
            .in1(N__13308),
            .in2(N__13290),
            .in3(N__13253),
            .lcout(\uart_frame_decoder.state_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23849),
            .ce(),
            .sr(N__23349));
    defparam \ppm_encoder_1.rudder_11_LC_4_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_4_21_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_4_21_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_4_21_4  (
            .in0(N__13209),
            .in1(N__13185),
            .in2(N__17460),
            .in3(N__18406),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23849),
            .ce(),
            .sr(N__23349));
    defparam \uart_frame_decoder.source_data_valid_LC_4_21_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_data_valid_LC_4_21_7 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \uart_frame_decoder.source_data_valid_LC_4_21_7  (
            .in0(N__13155),
            .in1(N__13117),
            .in2(N__14932),
            .in3(N__13011),
            .lcout(frame_decoder_dv_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23849),
            .ce(),
            .sr(N__23349));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2  (
            .in0(N__15315),
            .in1(N__20256),
            .in2(N__14865),
            .in3(N__20151),
            .lcout(\ppm_encoder_1.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_7_LC_4_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_4_22_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_4_22_6  (
            .in0(N__13749),
            .in1(N__13728),
            .in2(N__17461),
            .in3(N__17147),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23846),
            .ce(),
            .sr(N__23354));
    defparam \ppm_encoder_1.aileron_11_LC_4_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_4_23_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_4_23_0 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_4_23_0  (
            .in0(N__17435),
            .in1(N__13656),
            .in2(N__19405),
            .in3(N__13674),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23840),
            .ce(),
            .sr(N__23360));
    defparam \ppm_encoder_1.throttle_6_LC_4_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_4_23_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_4_23_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_4_23_1  (
            .in0(N__17434),
            .in1(N__13848),
            .in2(_gnd_net_),
            .in3(N__15371),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23840),
            .ce(),
            .sr(N__23360));
    defparam \ppm_encoder_1.rudder_6_LC_4_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_4_23_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_4_23_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_4_23_3  (
            .in0(N__17433),
            .in1(N__13533),
            .in2(_gnd_net_),
            .in3(N__19235),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23840),
            .ce(),
            .sr(N__23360));
    defparam \scaler_3.source_data_1_4_LC_4_23_5 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_4_LC_4_23_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_4_LC_4_23_5 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_3.source_data_1_4_LC_4_23_5  (
            .in0(N__14933),
            .in1(N__13509),
            .in2(N__14624),
            .in3(N__13472),
            .lcout(scaler_3_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23840),
            .ce(),
            .sr(N__23360));
    defparam \ppm_encoder_1.elevator_6_LC_4_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_4_23_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_4_23_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_4_23_7  (
            .in0(N__17432),
            .in1(N__13770),
            .in2(_gnd_net_),
            .in3(N__14735),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23840),
            .ce(),
            .sr(N__23360));
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_4_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_4_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_c_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__14765),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_4_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_4_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__17105),
            .in2(_gnd_net_),
            .in3(N__13443),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_4_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_4_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_4_24_2  (
            .in0(_gnd_net_),
            .in1(N__15929),
            .in2(_gnd_net_),
            .in3(N__13440),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_4_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_4_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_4_24_3  (
            .in0(_gnd_net_),
            .in1(N__14810),
            .in2(_gnd_net_),
            .in3(N__13437),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_4_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_4_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_4_24_4  (
            .in0(_gnd_net_),
            .in1(N__13589),
            .in2(_gnd_net_),
            .in3(N__13677),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_4_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_4_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__13673),
            .in2(_gnd_net_),
            .in3(N__13650),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_4_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_4_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_4_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15992),
            .in3(N__13647),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_4_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_4_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_4_24_7  (
            .in0(_gnd_net_),
            .in1(N__15839),
            .in2(N__24757),
            .in3(N__13644),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_4_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_4_25_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_4_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_4_25_0  (
            .in0(_gnd_net_),
            .in1(N__13641),
            .in2(_gnd_net_),
            .in3(N__13629),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23829),
            .ce(N__16253),
            .sr(N__23369));
    defparam \ppm_encoder_1.throttle_10_LC_4_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_4_26_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_4_26_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_4_26_0  (
            .in0(N__13782),
            .in1(N__13797),
            .in2(N__19958),
            .in3(N__17486),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.rudder_10_LC_4_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_4_26_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_4_26_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_4_26_2  (
            .in0(N__13626),
            .in1(N__13620),
            .in2(N__19931),
            .in3(N__17484),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.aileron_10_LC_4_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_4_26_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_4_26_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_4_26_3  (
            .in0(N__13593),
            .in1(N__13572),
            .in2(N__17529),
            .in3(N__15649),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.rudder_13_LC_4_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_4_26_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_4_26_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_4_26_4  (
            .in0(N__13563),
            .in1(N__13539),
            .in2(N__20663),
            .in3(N__17485),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.elevator_12_LC_4_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_4_26_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_4_26_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_4_26_5  (
            .in0(N__13875),
            .in1(N__13899),
            .in2(N__17530),
            .in3(N__19036),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.elevator_9_LC_4_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_4_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_4_26_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_4_26_6  (
            .in0(N__13692),
            .in1(N__13713),
            .in2(N__14864),
            .in3(N__17483),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.throttle_9_LC_4_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_4_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_4_26_7 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_4_26_7  (
            .in0(N__17476),
            .in1(N__13824),
            .in2(N__19010),
            .in3(N__13809),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23824),
            .ce(),
            .sr(N__23376));
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_4_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_4_27_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_c_LC_4_27_0  (
            .in0(_gnd_net_),
            .in1(N__13769),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_4_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_4_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_4_27_1  (
            .in0(_gnd_net_),
            .in1(N__13748),
            .in2(_gnd_net_),
            .in3(N__13719),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_4_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_4_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_4_27_2  (
            .in0(_gnd_net_),
            .in1(N__16133),
            .in2(_gnd_net_),
            .in3(N__13716),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_4_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_4_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_4_27_3  (
            .in0(_gnd_net_),
            .in1(N__13709),
            .in2(_gnd_net_),
            .in3(N__13686),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_4_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_4_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_4_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_4_27_4  (
            .in0(_gnd_net_),
            .in1(N__15266),
            .in2(_gnd_net_),
            .in3(N__13683),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_4_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_4_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_4_27_5  (
            .in0(_gnd_net_),
            .in1(N__15716),
            .in2(_gnd_net_),
            .in3(N__13680),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_4_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_4_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_4_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_4_27_6  (
            .in0(_gnd_net_),
            .in1(N__13898),
            .in2(_gnd_net_),
            .in3(N__13869),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_4_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_4_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_4_27_7  (
            .in0(_gnd_net_),
            .in1(N__15776),
            .in2(N__24769),
            .in3(N__13866),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_4_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_4_28_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_4_28_0  (
            .in0(_gnd_net_),
            .in1(N__13863),
            .in2(_gnd_net_),
            .in3(N__13851),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23814),
            .ce(N__16266),
            .sr(N__23391));
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_4_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_4_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_c_LC_4_29_0  (
            .in0(_gnd_net_),
            .in1(N__13841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_29_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_29_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_29_1  (
            .in0(_gnd_net_),
            .in1(N__16649),
            .in2(_gnd_net_),
            .in3(N__13830),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_29_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_29_2  (
            .in0(_gnd_net_),
            .in1(N__15878),
            .in2(_gnd_net_),
            .in3(N__13827),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_29_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_29_3  (
            .in0(_gnd_net_),
            .in1(N__13820),
            .in2(_gnd_net_),
            .in3(N__13800),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_29_4  (
            .in0(_gnd_net_),
            .in1(N__13793),
            .in2(_gnd_net_),
            .in3(N__13773),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_29_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_29_5  (
            .in0(_gnd_net_),
            .in1(N__16016),
            .in2(_gnd_net_),
            .in3(N__13998),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_29_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_29_6  (
            .in0(_gnd_net_),
            .in1(N__14990),
            .in2(_gnd_net_),
            .in3(N__13995),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_29_7  (
            .in0(_gnd_net_),
            .in1(N__14972),
            .in2(N__24770),
            .in3(N__13992),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_30_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_30_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_4_30_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_4_30_0  (
            .in0(_gnd_net_),
            .in1(N__13989),
            .in2(_gnd_net_),
            .in3(N__13983),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23802),
            .ce(N__16262),
            .sr(N__23400));
    defparam \uart_sync.aux_1__0__0_LC_5_8_2 .C_ON=1'b0;
    defparam \uart_sync.aux_1__0__0_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_1__0__0_LC_5_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_1__0__0_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15387),
            .lcout(\uart_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23882),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_0_LC_5_13_6 .C_ON=1'b0;
    defparam \uart.timer_Count_0_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_0_LC_5_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart.timer_Count_0_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14142),
            .lcout(\uart.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23877),
            .ce(),
            .sr(N__14184));
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_5_15_0 .C_ON=1'b1;
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart.un4_timer_Count_1_cry_1_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__13974),
            .in2(N__14148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\uart.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_2_LC_5_15_1 .C_ON=1'b1;
    defparam \uart.timer_Count_2_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_2_LC_5_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_2_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__13949),
            .in2(_gnd_net_),
            .in3(N__13929),
            .lcout(\uart.timer_CountZ0Z_2 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_1 ),
            .carryout(\uart.un4_timer_Count_1_cry_2 ),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_3_LC_5_15_2 .C_ON=1'b1;
    defparam \uart.timer_Count_3_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_3_LC_5_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_3_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__13924),
            .in2(_gnd_net_),
            .in3(N__13902),
            .lcout(\uart.timer_CountZ0Z_3 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_2 ),
            .carryout(\uart.un4_timer_Count_1_cry_3 ),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_4_LC_5_15_3 .C_ON=1'b1;
    defparam \uart.timer_Count_4_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_4_LC_5_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_4_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__14118),
            .in2(_gnd_net_),
            .in3(N__14331),
            .lcout(\uart.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_3 ),
            .carryout(\uart.un4_timer_Count_1_cry_4 ),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_5_LC_5_15_4 .C_ON=1'b1;
    defparam \uart.timer_Count_5_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_5_LC_5_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_5_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__14327),
            .in2(_gnd_net_),
            .in3(N__14301),
            .lcout(\uart.timer_CountZ0Z_5 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_4 ),
            .carryout(\uart.un4_timer_Count_1_cry_5 ),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_6_LC_5_15_5 .C_ON=1'b1;
    defparam \uart.timer_Count_6_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_6_LC_5_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_6_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__14289),
            .in2(_gnd_net_),
            .in3(N__14256),
            .lcout(\uart.timer_CountZ0Z_6 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_5 ),
            .carryout(\uart.un4_timer_Count_1_cry_6 ),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_7_LC_5_15_6 .C_ON=1'b0;
    defparam \uart.timer_Count_7_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_7_LC_5_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart.timer_Count_7_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__14233),
            .in2(_gnd_net_),
            .in3(N__14253),
            .lcout(\uart.timer_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23870),
            .ce(),
            .sr(N__14176));
    defparam \uart.timer_Count_RNIQ9BL_0_LC_5_16_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIQ9BL_0_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIQ9BL_0_LC_5_16_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.timer_Count_RNIQ9BL_0_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__14144),
            .in2(_gnd_net_),
            .in3(N__14117),
            .lcout(\uart.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_5_17_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_5_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__14079),
            .in2(N__14057),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_5_17_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_5_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__14034),
            .in2(_gnd_net_),
            .in3(N__14016),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_5_17_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_5_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__14013),
            .in2(_gnd_net_),
            .in3(N__14001),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_5_17_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_5_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__14468),
            .in2(_gnd_net_),
            .in3(N__14457),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_5_17_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_5_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__14454),
            .in2(_gnd_net_),
            .in3(N__14442),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_5_17_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_5_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__14439),
            .in2(_gnd_net_),
            .in3(N__14427),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_5_17_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_5_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__14424),
            .in2(_gnd_net_),
            .in3(N__14412),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_5_17_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_5_17_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_5_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__14409),
            .in2(_gnd_net_),
            .in3(N__14397),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__23861),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_5_18_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_5_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__14393),
            .in2(_gnd_net_),
            .in3(N__14379),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_5_18_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_5_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__14376),
            .in2(_gnd_net_),
            .in3(N__14364),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_5_18_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_5_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__14361),
            .in2(_gnd_net_),
            .in3(N__14349),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_5_18_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_5_18_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_5_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__14345),
            .in2(_gnd_net_),
            .in3(N__14334),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_5_18_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_5_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__14663),
            .in2(_gnd_net_),
            .in3(N__14568),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_5_18_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_5_18_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_5_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__14565),
            .in2(_gnd_net_),
            .in3(N__14553),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_5_18_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_5_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(N__14687),
            .in2(_gnd_net_),
            .in3(N__14550),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_5_18_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_5_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(N__14546),
            .in2(_gnd_net_),
            .in3(N__14535),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__23856),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_5_19_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_5_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__14531),
            .in2(_gnd_net_),
            .in3(N__14517),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__23852),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_5_19_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_5_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__14510),
            .in2(_gnd_net_),
            .in3(N__14496),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__23852),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_5_19_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_5_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__14697),
            .in2(_gnd_net_),
            .in3(N__14493),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__23852),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_5_19_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_5_19_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_5_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(N__14486),
            .in2(_gnd_net_),
            .in3(N__14472),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__23852),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_5_19_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_5_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(N__14675),
            .in2(_gnd_net_),
            .in3(N__14700),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23852),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_5_19_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_5_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_5_19_5  (
            .in0(N__14696),
            .in1(N__14688),
            .in2(N__14676),
            .in3(N__14664),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIJL8F_4_LC_5_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIJL8F_4_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIJL8F_4_LC_5_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIJL8F_4_LC_5_21_0  (
            .in0(N__14792),
            .in1(N__14780),
            .in2(_gnd_net_),
            .in3(N__18826),
            .lcout(\ppm_encoder_1.N_462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_4_LC_5_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_4_LC_5_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_4_LC_5_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_4_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15153),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23847),
            .ce(N__16244),
            .sr(N__23346));
    defparam \ppm_encoder_1.elevator_esr_4_LC_5_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_4_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_4_LC_5_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_4_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14628),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23847),
            .ce(N__16244),
            .sr(N__23346));
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_5_21_4 .C_ON=1'b0;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_5_21_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_5_21_4  (
            .in0(N__15184),
            .in1(N__14607),
            .in2(_gnd_net_),
            .in3(N__15230),
            .lcout(\scaler_2.un2_source_data_0_cry_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_5_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_5_22_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_5_22_0 .LUT_INIT=16'b1110111010101111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_5_22_0  (
            .in0(N__23504),
            .in1(N__18854),
            .in2(N__16374),
            .in3(N__21210),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23841),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_5_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_5_22_2 .LUT_INIT=16'b1100110000111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_5_22_2  (
            .in0(N__17310),
            .in1(N__22132),
            .in2(N__24090),
            .in3(N__21967),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNINGL11_6_LC_5_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNINGL11_6_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNINGL11_6_LC_5_22_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ppm_encoder_1.throttle_RNINGL11_6_LC_5_22_4  (
            .in0(N__15367),
            .in1(N__19230),
            .in2(_gnd_net_),
            .in3(N__19538),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_rn_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_5_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_5_22_5 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_5_22_5  (
            .in0(N__20150),
            .in1(N__14793),
            .in2(N__22134),
            .in3(N__14781),
            .lcout(\ppm_encoder_1.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_22_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_22_6  (
            .in0(N__23505),
            .in1(N__19539),
            .in2(N__18294),
            .in3(N__21209),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23841),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_5_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_5_23_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_5_23_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_5_23_1  (
            .in0(N__14769),
            .in1(N__17487),
            .in2(_gnd_net_),
            .in3(N__14748),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23835),
            .ce(),
            .sr(N__23355));
    defparam \ppm_encoder_1.elevator_RNIDJ141_6_LC_5_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIDJ141_6_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIDJ141_6_LC_5_23_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIDJ141_6_LC_5_23_2  (
            .in0(N__14747),
            .in1(N__17193),
            .in2(N__14739),
            .in3(N__17883),
            .lcout(\ppm_encoder_1.pulses2count_9_0_o2_0_6 ),
            .ltout(\ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI0LED3_6_LC_5_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI0LED3_6_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI0LED3_6_LC_5_23_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.throttle_RNI0LED3_6_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(N__14706),
            .in2(N__14721),
            .in3(N__14718),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNID1DC5_6_LC_5_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID1DC5_6_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID1DC5_6_LC_5_23_4 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID1DC5_6_LC_5_23_4  (
            .in0(N__17718),
            .in1(N__19187),
            .in2(N__14712),
            .in3(N__17051),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI6UPC6_6_LC_5_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI6UPC6_6_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI6UPC6_6_LC_5_23_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI6UPC6_6_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14709),
            .in3(N__17933),
            .lcout(\ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNISGN71_6_LC_5_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNISGN71_6_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNISGN71_6_LC_5_23_7 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \ppm_encoder_1.rudder_RNISGN71_6_LC_5_23_7  (
            .in0(N__18763),
            .in1(N__19231),
            .in2(N__18881),
            .in3(N__19540),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_sn_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI31EQ5_9_LC_5_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI31EQ5_9_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI31EQ5_9_LC_5_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI31EQ5_9_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__17216),
            .in2(_gnd_net_),
            .in3(N__14826),
            .lcout(\ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNICBGI_10_LC_5_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNICBGI_10_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNICBGI_10_LC_5_24_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.throttle_RNICBGI_10_LC_5_24_1  (
            .in0(N__19954),
            .in1(N__18876),
            .in2(_gnd_net_),
            .in3(N__18782),
            .lcout(\ppm_encoder_1.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI55NT_10_LC_5_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI55NT_10_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI55NT_10_LC_5_24_2 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \ppm_encoder_1.elevator_RNI55NT_10_LC_5_24_2  (
            .in0(N__18783),
            .in1(N__15674),
            .in2(N__15650),
            .in3(N__18877),
            .lcout(),
            .ltout(\ppm_encoder_1.N_414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNI5GRA2_10_LC_5_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNI5GRA2_10_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNI5GRA2_10_LC_5_24_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \ppm_encoder_1.rudder_RNI5GRA2_10_LC_5_24_3  (
            .in0(N__19927),
            .in1(N__14880),
            .in2(N__14874),
            .in3(N__19625),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITDM64_10_LC_5_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITDM64_10_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITDM64_10_LC_5_24_4 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITDM64_10_LC_5_24_4  (
            .in0(N__22526),
            .in1(N__17713),
            .in2(N__14871),
            .in3(N__17060),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJ2JB5_10_LC_5_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJ2JB5_10_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJ2JB5_10_LC_5_24_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJ2JB5_10_LC_5_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14868),
            .in3(N__17834),
            .lcout(\ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI4MTK_9_LC_5_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI4MTK_9_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI4MTK_9_LC_5_25_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNI4MTK_9_LC_5_25_0  (
            .in0(N__19000),
            .in1(N__18776),
            .in2(_gnd_net_),
            .in3(N__18897),
            .lcout(\ppm_encoder_1.N_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNILQ941_9_LC_5_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNILQ941_9_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNILQ941_9_LC_5_25_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \ppm_encoder_1.elevator_RNILQ941_9_LC_5_25_1  (
            .in0(N__18898),
            .in1(N__14854),
            .in2(N__18788),
            .in3(N__15310),
            .lcout(),
            .ltout(\ppm_encoder_1.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNI5BFJ2_9_LC_5_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNI5BFJ2_9_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNI5BFJ2_9_LC_5_25_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \ppm_encoder_1.rudder_RNI5BFJ2_9_LC_5_25_2  (
            .in0(N__18955),
            .in1(N__14838),
            .in2(N__14832),
            .in3(N__19624),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILQDI4_9_LC_5_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILQDI4_9_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILQDI4_9_LC_5_25_3 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILQDI4_9_LC_5_25_3  (
            .in0(N__24161),
            .in1(N__17717),
            .in2(N__14829),
            .in3(N__17059),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_9_LC_5_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_5_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_5_25_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_5_25_5  (
            .in0(N__14820),
            .in1(N__14814),
            .in2(N__17540),
            .in3(N__15311),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23825),
            .ce(),
            .sr(N__23364));
    defparam \ppm_encoder_1.rudder_9_LC_5_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_5_26_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_5_26_1  (
            .in0(N__15297),
            .in1(N__15288),
            .in2(N__18965),
            .in3(N__17508),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23820),
            .ce(),
            .sr(N__23370));
    defparam \ppm_encoder_1.elevator_10_LC_5_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_5_26_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_5_26_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_5_26_4  (
            .in0(N__15267),
            .in1(N__15243),
            .in2(N__17541),
            .in3(N__15673),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23820),
            .ce(),
            .sr(N__23370));
    defparam \scaler_2.source_data_1_4_LC_5_26_6 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_4_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_4_LC_5_26_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_2.source_data_1_4_LC_5_26_6  (
            .in0(N__14948),
            .in1(N__15237),
            .in2(N__15152),
            .in3(N__15195),
            .lcout(scaler_2_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23820),
            .ce(),
            .sr(N__23370));
    defparam \ppm_encoder_1.rudder_12_LC_5_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_5_26_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_5_26_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_5_26_7  (
            .in0(N__15135),
            .in1(N__15117),
            .in2(N__18493),
            .in3(N__17507),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23820),
            .ce(),
            .sr(N__23370));
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_5_27_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_5_27_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_5_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_4_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15105),
            .lcout(frame_decoder_CH1data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23815),
            .ce(N__15024),
            .sr(N__23377));
    defparam \ppm_encoder_1.throttle_12_LC_5_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_5_28_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_5_28_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_5_28_6  (
            .in0(N__15000),
            .in1(N__14994),
            .in2(N__17560),
            .in3(N__19360),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23809),
            .ce(),
            .sr(N__23383));
    defparam \ppm_encoder_1.throttle_13_LC_5_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_5_28_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_5_28_7 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_5_28_7  (
            .in0(N__14979),
            .in1(N__14961),
            .in2(N__15867),
            .in3(N__17539),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23809),
            .ce(),
            .sr(N__23383));
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_5_30_5 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_5_30_5 .SEQ_MODE=4'b0000;
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_5_30_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_1.source_data_1_esr_ctle_14_LC_5_30_5  (
            .in0(_gnd_net_),
            .in1(N__14939),
            .in2(_gnd_net_),
            .in3(N__23492),
            .lcout(frame_decoder_dv_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.aux_0__0__0_LC_7_6_2 .C_ON=1'b0;
    defparam \uart_sync.aux_0__0__0_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_0__0__0_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_0__0__0_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15414),
            .lcout(\uart_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23883),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__17462),
            .in2(_gnd_net_),
            .in3(N__23491),
            .lcout(\ppm_encoder_1.scaler_1_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_20_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_20_6  (
            .in0(N__18780),
            .in1(N__15375),
            .in2(N__15351),
            .in3(N__18893),
            .lcout(\ppm_encoder_1.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7JM64_11_LC_7_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7JM64_11_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7JM64_11_LC_7_21_0 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7JM64_11_LC_7_21_0  (
            .in0(N__15333),
            .in1(N__17712),
            .in2(N__20043),
            .in3(N__17050),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIV8JB5_11_LC_7_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIV8JB5_11_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIV8JB5_11_LC_7_21_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIV8JB5_11_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15336),
            .in3(N__19262),
            .lcout(\ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIEKRA2_11_LC_7_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIEKRA2_11_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIEKRA2_11_LC_7_21_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \ppm_encoder_1.rudder_RNIEKRA2_11_LC_7_21_2  (
            .in0(N__20397),
            .in1(N__15729),
            .in2(N__18413),
            .in3(N__15564),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_21_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_21_4  (
            .in0(N__24056),
            .in1(N__21785),
            .in2(N__20931),
            .in3(N__21223),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNII84K_4_LC_7_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNII84K_4_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNII84K_4_LC_7_21_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNII84K_4_LC_7_21_6  (
            .in0(N__17192),
            .in1(N__19877),
            .in2(_gnd_net_),
            .in3(N__20675),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNIGT971_LC_7_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNIGT971_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNIGT971_LC_7_21_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNIGT971_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__20242),
            .in2(N__15327),
            .in3(N__15324),
            .lcout(\ppm_encoder_1.un2_throttle_iv_i_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_7_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_7_22_0 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_7_22_0  (
            .in0(N__19587),
            .in1(N__22632),
            .in2(N__17817),
            .in3(N__21207),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_7_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_7_22_1 .LUT_INIT=16'b1100110010011001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_7_22_1  (
            .in0(N__21208),
            .in1(N__20458),
            .in2(_gnd_net_),
            .in3(N__17737),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_7_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_7_22_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_7_22_2 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_7_22_2  (
            .in0(N__20459),
            .in1(N__16918),
            .in2(N__15429),
            .in3(N__16793),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23830),
            .ce(),
            .sr(N__23350));
    defparam \ppm_encoder_1.init_pulses_4_LC_7_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_7_22_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_7_22_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_7_22_3  (
            .in0(N__16792),
            .in1(N__17973),
            .in2(N__16923),
            .in3(N__15471),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23830),
            .ce(),
            .sr(N__23350));
    defparam \ppm_encoder_1.init_pulses_RNIR7863_4_LC_7_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR7863_4_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR7863_4_LC_7_22_4 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR7863_4_LC_7_22_4  (
            .in0(N__17710),
            .in1(N__15426),
            .in2(N__22640),
            .in3(N__17044),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI398E4_4_LC_7_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI398E4_4_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI398E4_4_LC_7_22_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI398E4_4_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15420),
            .in3(N__16449),
            .lcout(\ppm_encoder_1.init_pulses_RNI398E4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI83R42_0_LC_7_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI83R42_0_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI83R42_0_LC_7_22_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI83R42_0_LC_7_22_6  (
            .in0(N__17735),
            .in1(N__20460),
            .in2(_gnd_net_),
            .in3(N__21205),
            .lcout(\ppm_encoder_1.init_pulses_RNI83R42Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR0RR1_13_LC_7_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0RR1_13_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0RR1_13_LC_7_22_7 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0RR1_13_LC_7_22_7  (
            .in0(N__21206),
            .in1(N__17709),
            .in2(N__21351),
            .in3(N__17736),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_0_LC_7_23_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_0_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_0_LC_7_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIMR0V_0_0_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_7_23_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_7_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__17076),
            .in2(N__17283),
            .in3(N__15417),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_7_23_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_7_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__16323),
            .in2(N__18054),
            .in3(N__15483),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_7_23_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_7_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__16956),
            .in2(N__17265),
            .in3(N__15480),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_7_23_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_7_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__15477),
            .in2(N__16448),
            .in3(N__15465),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_7_23_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_7_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__16308),
            .in2(N__16188),
            .in3(N__15462),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_7_23_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_7_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(N__15459),
            .in2(N__17934),
            .in3(N__15450),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_7_23_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_7_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(N__16380),
            .in2(N__17247),
            .in3(N__15447),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_7_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_7_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__16164),
            .in2(N__18618),
            .in3(N__15444),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_7_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_7_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(N__15441),
            .in2(N__17220),
            .in3(N__15432),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_7_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_7_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(N__15537),
            .in2(N__17838),
            .in3(N__15528),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_7_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_7_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_7_24_3  (
            .in0(_gnd_net_),
            .in1(N__15525),
            .in2(N__19266),
            .in3(N__15516),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_7_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_7_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_7_24_4  (
            .in0(_gnd_net_),
            .in1(N__16389),
            .in2(N__19296),
            .in3(N__15513),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_7_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_7_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__18156),
            .in2(N__15792),
            .in3(N__15510),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_14_LC_7_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_2_14_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_14_LC_7_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_14_LC_7_24_6  (
            .in0(_gnd_net_),
            .in1(N__17583),
            .in2(N__15585),
            .in3(N__15507),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_7_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_7_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_7_24_7  (
            .in0(_gnd_net_),
            .in1(N__16476),
            .in2(N__15576),
            .in3(N__15504),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_7_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_7_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_7_25_0  (
            .in0(_gnd_net_),
            .in1(N__17757),
            .in2(_gnd_net_),
            .in3(N__15501),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_7_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_7_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__15498),
            .in2(_gnd_net_),
            .in3(N__15489),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_7_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_7_25_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_7_25_2  (
            .in0(N__20875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15486),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISRB55_14_LC_7_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISRB55_14_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISRB55_14_LC_7_25_3 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISRB55_14_LC_7_25_3  (
            .in0(N__17715),
            .in1(N__21461),
            .in2(N__21512),
            .in3(N__16317),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINK8A6_14_LC_7_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINK8A6_14_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINK8A6_14_LC_7_25_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINK8A6_14_LC_7_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15588),
            .in3(N__17579),
            .lcout(\ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIN4HJ_12_LC_7_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIN4HJ_12_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIN4HJ_12_LC_7_25_5 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \ppm_encoder_1.elevator_RNIN4HJ_12_LC_7_25_5  (
            .in0(N__20104),
            .in1(N__19043),
            .in2(N__19373),
            .in3(N__20218),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJJM71_15_LC_7_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJJM71_15_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJJM71_15_LC_7_25_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJJM71_15_LC_7_25_6  (
            .in0(N__21813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16472),
            .lcout(\ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNI3HMS_11_LC_7_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNI3HMS_11_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNI3HMS_11_LC_7_25_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.aileron_RNI3HMS_11_LC_7_25_7  (
            .in0(N__20103),
            .in1(N__20217),
            .in2(_gnd_net_),
            .in3(N__19406),
            .lcout(\ppm_encoder_1.N_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_7_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_7_26_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_7_26_0 .LUT_INIT=16'b1110111111001101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_7_26_0  (
            .in0(N__21230),
            .in1(N__23513),
            .in2(N__16363),
            .in3(N__21929),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNIUAMB2_14_LC_7_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNIUAMB2_14_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNIUAMB2_14_LC_7_26_1 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNIUAMB2_14_LC_7_26_1  (
            .in0(N__22121),
            .in1(N__21880),
            .in2(N__15552),
            .in3(N__16404),
            .lcout(\ppm_encoder_1.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIFN3K_2_LC_7_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIFN3K_2_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIFN3K_2_LC_7_26_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIFN3K_2_LC_7_26_2  (
            .in0(N__20235),
            .in1(N__20119),
            .in2(_gnd_net_),
            .in3(N__19830),
            .lcout(\ppm_encoder_1.N_443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_LC_7_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_LC_7_26_3 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_LC_7_26_3  (
            .in0(N__21928),
            .in1(N__20236),
            .in2(N__23532),
            .in3(N__21231),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_i_0_LC_7_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_i_0_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_i_0_LC_7_26_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_i_0_LC_7_26_4  (
            .in0(N__21882),
            .in1(N__19745),
            .in2(_gnd_net_),
            .in3(N__20349),
            .lcout(\ppm_encoder_1.N_114 ),
            .ltout(\ppm_encoder_1.N_114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep2_LC_7_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep2_LC_7_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep2_LC_7_26_5 .LUT_INIT=16'b1110111011001111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep2_LC_7_26_5  (
            .in0(N__20120),
            .in1(N__23523),
            .in2(N__15678),
            .in3(N__21233),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_26_6 .LUT_INIT=16'b0010011100000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_26_6  (
            .in0(N__21881),
            .in1(N__15675),
            .in2(N__15651),
            .in3(N__22122),
            .lcout(\ppm_encoder_1.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_7_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_7_26_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_7_26_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_7_26_7  (
            .in0(N__20350),
            .in1(N__18289),
            .in2(N__23533),
            .in3(N__21232),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIFNBA1_LC_7_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIFNBA1_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIFNBA1_LC_7_27_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIFNBA1_LC_7_27_0  (
            .in0(N__19769),
            .in1(N__24558),
            .in2(N__20815),
            .in3(N__24411),
            .lcout(\ppm_encoder_1.N_348 ),
            .ltout(\ppm_encoder_1.N_348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_7_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_7_27_1 .LUT_INIT=16'b1111100011110010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_7_27_1  (
            .in0(N__16843),
            .in1(N__18321),
            .in2(N__15621),
            .in3(N__18102),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_18_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_7_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_7_27_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_7_27_2 .LUT_INIT=16'b0000110100001100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_7_27_2  (
            .in0(N__15606),
            .in1(N__15618),
            .in2(N__15609),
            .in3(N__17716),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23803),
            .ce(),
            .sr(N__23378));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_3 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_3  (
            .in0(N__21229),
            .in1(N__20348),
            .in2(N__21773),
            .in3(N__21602),
            .lcout(\ppm_encoder_1.init_pulses_18_i_a2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIMOAF1_LC_7_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIMOAF1_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIMOAF1_LC_7_27_6 .LUT_INIT=16'b1111111101100101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIMOAF1_LC_7_27_6  (
            .in0(N__20347),
            .in1(N__19770),
            .in2(N__21620),
            .in3(N__21228),
            .lcout(\ppm_encoder_1.N_241 ),
            .ltout(\ppm_encoder_1.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_7_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_7_27_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_7_27_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_7_27_7  (
            .in0(N__16791),
            .in1(N__15600),
            .in2(N__15591),
            .in3(N__18369),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23803),
            .ce(),
            .sr(N__23378));
    defparam \ppm_encoder_1.elevator_RNIDBNT_13_LC_7_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIDBNT_13_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIDBNT_13_LC_7_28_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \ppm_encoder_1.elevator_RNIDBNT_13_LC_7_28_0  (
            .in0(N__15806),
            .in1(N__20241),
            .in2(N__15741),
            .in3(N__20128),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI06LN1_13_LC_7_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI06LN1_13_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI06LN1_13_LC_7_28_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \ppm_encoder_1.throttle_RNI06LN1_13_LC_7_28_1  (
            .in0(N__15866),
            .in1(N__21907),
            .in2(N__15849),
            .in3(N__22110),
            .lcout(\ppm_encoder_1.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_7_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_7_28_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_7_28_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_7_28_2  (
            .in0(N__15807),
            .in1(N__15846),
            .in2(N__17564),
            .in3(N__15822),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23796),
            .ce(),
            .sr(N__23384));
    defparam \ppm_encoder_1.rudder_RNIAAE02_13_LC_7_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIAAE02_13_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIAAE02_13_LC_7_28_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \ppm_encoder_1.rudder_RNIAAE02_13_LC_7_28_3  (
            .in0(N__20659),
            .in1(N__20362),
            .in2(_gnd_net_),
            .in3(N__17061),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJ94E4_13_LC_7_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJ94E4_13_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJ94E4_13_LC_7_28_4 .LUT_INIT=16'b0101011010101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJ94E4_13_LC_7_28_4  (
            .in0(N__21349),
            .in1(N__21287),
            .in2(N__15798),
            .in3(N__17714),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC11J5_13_LC_7_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC11J5_13_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC11J5_13_LC_7_28_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC11J5_13_LC_7_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15795),
            .in3(N__18145),
            .lcout(\ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_13_LC_7_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_7_28_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_7_28_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_7_28_6  (
            .in0(N__15740),
            .in1(N__15780),
            .in2(N__17565),
            .in3(N__15753),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23796),
            .ce(),
            .sr(N__23384));
    defparam \ppm_encoder_1.elevator_RNIL2HJ_11_LC_7_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIL2HJ_11_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIL2HJ_11_LC_7_29_0 .LUT_INIT=16'b0100010000001100;
    LogicCell40 \ppm_encoder_1.elevator_RNIL2HJ_11_LC_7_29_0  (
            .in0(N__18457),
            .in1(N__20127),
            .in2(N__19988),
            .in3(N__20240),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_11_LC_7_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_7_29_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_7_29_1 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_7_29_1  (
            .in0(N__15720),
            .in1(N__18458),
            .in2(N__15693),
            .in3(N__17534),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23791),
            .ce(),
            .sr(N__23392));
    defparam \ppm_encoder_1.throttle_11_LC_7_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_7_29_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_7_29_2 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_7_29_2  (
            .in0(N__19984),
            .in1(N__16023),
            .in2(N__17559),
            .in3(N__16005),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23791),
            .ce(),
            .sr(N__23392));
    defparam \ppm_encoder_1.aileron_12_LC_8_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_8_19_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_8_19_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_8_19_1  (
            .in0(N__15996),
            .in1(N__15972),
            .in2(N__17552),
            .in3(N__19081),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23842),
            .ce(),
            .sr(N__23344));
    defparam \ppm_encoder_1.throttle_2_LC_8_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_8_19_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_8_19_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__17520),
            .in2(_gnd_net_),
            .in3(N__20614),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23842),
            .ce(),
            .sr(N__23344));
    defparam \ppm_encoder_1.throttle_RNI3LTK_8_LC_8_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI3LTK_8_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI3LTK_8_LC_8_20_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNI3LTK_8_LC_8_20_0  (
            .in0(N__18427),
            .in1(N__18759),
            .in2(_gnd_net_),
            .in3(N__18885),
            .lcout(\ppm_encoder_1.N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIJO941_8_LC_8_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIJO941_8_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIJO941_8_LC_8_20_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIJO941_8_LC_8_20_1  (
            .in0(N__18886),
            .in1(N__18589),
            .in2(N__18781),
            .in3(N__18571),
            .lcout(),
            .ltout(\ppm_encoder_1.N_417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNI17FJ2_8_LC_8_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNI17FJ2_8_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNI17FJ2_8_LC_8_20_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \ppm_encoder_1.rudder_RNI17FJ2_8_LC_8_20_2  (
            .in0(N__18550),
            .in1(N__15957),
            .in2(N__15951),
            .in3(N__19597),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGLDI4_8_LC_8_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGLDI4_8_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGLDI4_8_LC_8_20_3 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGLDI4_8_LC_8_20_3  (
            .in0(N__22692),
            .in1(N__17705),
            .in2(N__15948),
            .in3(N__17049),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_8_LC_8_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_8_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_8_20_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_8_20_5  (
            .in0(N__15945),
            .in1(N__15933),
            .in2(N__17561),
            .in3(N__18572),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23836),
            .ce(),
            .sr(N__23347));
    defparam \ppm_encoder_1.throttle_8_LC_8_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_8_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_8_20_6 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_8_20_6  (
            .in0(N__18428),
            .in1(N__15912),
            .in2(N__15894),
            .in3(N__17548),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23836),
            .ce(),
            .sr(N__23347));
    defparam \ppm_encoder_1.elevator_8_LC_8_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_8_20_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_8_20_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_8_20_7  (
            .in0(N__16155),
            .in1(N__16140),
            .in2(N__17562),
            .in3(N__18590),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23836),
            .ce(),
            .sr(N__23347));
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_21_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_5_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16113),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23831),
            .ce(N__16243),
            .sr(N__23351));
    defparam \ppm_encoder_1.rudder_esr_4_LC_8_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_8_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_8_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16098),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23831),
            .ce(N__16243),
            .sr(N__23351));
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_4_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16074),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23831),
            .ce(N__16243),
            .sr(N__23351));
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_21_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ppm_encoder_1.throttle_esr_5_LC_8_21_3  (
            .in0(N__16050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23831),
            .ce(N__16243),
            .sr(N__23351));
    defparam \ppm_encoder_1.aileron_esr_RNITLTI_5_LC_8_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNITLTI_5_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNITLTI_5_LC_8_22_0 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNITLTI_5_LC_8_22_0  (
            .in0(N__17879),
            .in1(N__16287),
            .in2(N__16038),
            .in3(N__17188),
            .lcout(\ppm_encoder_1.pulses2count_9_i_o2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNI4IR61_5_LC_8_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNI4IR61_5_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNI4IR61_5_LC_8_22_1 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNI4IR61_5_LC_8_22_1  (
            .in0(N__18741),
            .in1(N__19554),
            .in2(N__22310),
            .in3(N__18902),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI8RGL2_5_LC_8_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI8RGL2_5_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI8RGL2_5_LC_8_22_2 .LUT_INIT=16'b0000110011111100;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI8RGL2_5_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__16302),
            .in2(N__16029),
            .in3(N__18920),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIK6FK4_5_LC_8_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIK6FK4_5_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIK6FK4_5_LC_8_22_3 .LUT_INIT=16'b1001100101101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIK6FK4_5_LC_8_22_3  (
            .in0(N__22569),
            .in1(N__17711),
            .in2(N__16026),
            .in3(N__17045),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT8FS5_5_LC_8_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT8FS5_5_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT8FS5_5_LC_8_22_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT8FS5_5_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__16184),
            .in2(N__16311),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI7JNR_5_LC_8_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI7JNR_5_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI7JNR_5_LC_8_22_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI7JNR_5_LC_8_22_5  (
            .in0(N__18932),
            .in1(N__22303),
            .in2(_gnd_net_),
            .in3(N__19553),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_5_LC_8_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_5_LC_8_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_5_LC_8_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_5_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16296),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23826),
            .ce(N__16254),
            .sr(N__23356));
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16281),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23826),
            .ce(N__16254),
            .sr(N__23356));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_8_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_8_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_8_23_0 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_8_23_0  (
            .in0(N__21974),
            .in1(N__18775),
            .in2(N__23534),
            .in3(N__21055),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23821),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI92081_5_LC_8_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI92081_5_LC_8_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI92081_5_LC_8_23_1 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI92081_5_LC_8_23_1  (
            .in0(N__21054),
            .in1(N__17807),
            .in2(N__22576),
            .in3(N__19603),
            .lcout(\ppm_encoder_1.N_252_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITQDQ5_8_LC_8_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITQDQ5_8_LC_8_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITQDQ5_8_LC_8_23_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITQDQ5_8_LC_8_23_2  (
            .in0(_gnd_net_),
            .in1(N__18611),
            .in2(_gnd_net_),
            .in3(N__16173),
            .lcout(\ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_8_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_8_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_8_23_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_8_23_3  (
            .in0(N__17864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17181),
            .lcout(\ppm_encoder_1.N_235 ),
            .ltout(\ppm_encoder_1.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_3_LC_8_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_3_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_3_LC_8_23_4 .LUT_INIT=16'b1111111111101011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_3_LC_8_23_4  (
            .in0(N__19860),
            .in1(N__19815),
            .in2(N__16158),
            .in3(N__21053),
            .lcout(\ppm_encoder_1.N_246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUBDK6_7_LC_8_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUBDK6_7_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUBDK6_7_LC_8_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUBDK6_7_LC_8_23_5  (
            .in0(_gnd_net_),
            .in1(N__17234),
            .in2(_gnd_net_),
            .in3(N__17199),
            .lcout(\ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_23_6 .LUT_INIT=16'b1111101011110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_23_6  (
            .in0(N__17183),
            .in1(N__16370),
            .in2(N__23535),
            .in3(N__21056),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23821),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_8_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_8_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_8_23_7 .LUT_INIT=16'b1100001111010011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_8_23_7  (
            .in0(N__17865),
            .in1(N__19859),
            .in2(N__19826),
            .in3(N__17182),
            .lcout(\ppm_encoder_1.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNI4IMS_12_LC_8_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNI4IMS_12_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNI4IMS_12_LC_8_24_0 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \ppm_encoder_1.aileron_RNI4IMS_12_LC_8_24_0  (
            .in0(N__20243),
            .in1(_gnd_net_),
            .in2(N__19088),
            .in3(N__20133),
            .lcout(),
            .ltout(\ppm_encoder_1.N_407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIIORA2_12_LC_8_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIIORA2_12_LC_8_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIIORA2_12_LC_8_24_1 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.rudder_RNIIORA2_12_LC_8_24_1  (
            .in0(N__16338),
            .in1(N__20398),
            .in2(N__16332),
            .in3(N__18494),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIUETK_2_LC_8_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIUETK_2_LC_8_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIUETK_2_LC_8_24_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.throttle_RNIUETK_2_LC_8_24_2  (
            .in0(N__20615),
            .in1(N__20132),
            .in2(_gnd_net_),
            .in3(N__18740),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7NRJ2_2_LC_8_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7NRJ2_2_LC_8_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7NRJ2_2_LC_8_24_3 .LUT_INIT=16'b1001100101101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7NRJ2_2_LC_8_24_3  (
            .in0(N__20540),
            .in1(N__17687),
            .in2(N__16329),
            .in3(N__17036),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIE48O3_2_LC_8_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIE48O3_2_LC_8_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIE48O3_2_LC_8_24_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIE48O3_2_LC_8_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16326),
            .in3(N__18040),
            .lcout(\ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIKMK32_14_LC_8_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIKMK32_14_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIKMK32_14_LC_8_24_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIKMK32_14_LC_8_24_5  (
            .in0(N__21540),
            .in1(N__20399),
            .in2(_gnd_net_),
            .in3(N__17037),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_8_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI81081_4_LC_8_24_6 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI81081_4_LC_8_24_6  (
            .in0(N__17805),
            .in1(N__22639),
            .in2(N__19620),
            .in3(N__21083),
            .lcout(\ppm_encoder_1.N_251_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_8_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_8_24_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_8_24_7 .LUT_INIT=16'b0100010100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_8_24_7  (
            .in0(N__23512),
            .in1(N__21167),
            .in2(N__18654),
            .in3(N__17806),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23816),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPNS41_13_LC_8_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPNS41_13_LC_8_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPNS41_13_LC_8_25_0 .LUT_INIT=16'b1101001011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPNS41_13_LC_8_25_0  (
            .in0(N__19713),
            .in1(N__21062),
            .in2(N__21336),
            .in3(N__19626),
            .lcout(\ppm_encoder_1.N_259_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI14O81_14_LC_8_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI14O81_14_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI14O81_14_LC_8_25_1 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI14O81_14_LC_8_25_1  (
            .in0(N__20222),
            .in1(N__16428),
            .in2(N__16419),
            .in3(N__20115),
            .lcout(\ppm_encoder_1.pulses2count_9_i_o2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICOM64_12_LC_8_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICOM64_12_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICOM64_12_LC_8_25_2 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICOM64_12_LC_8_25_2  (
            .in0(N__16398),
            .in1(N__17669),
            .in2(N__19337),
            .in3(N__17058),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI5FJB5_12_LC_8_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5FJB5_12_LC_8_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5FJB5_12_LC_8_25_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5FJB5_12_LC_8_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16392),
            .in3(N__19295),
            .lcout(\ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDCUU1_6_LC_8_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCUU1_6_LC_8_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCUU1_6_LC_8_25_4 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCUU1_6_LC_8_25_4  (
            .in0(N__17668),
            .in1(N__21064),
            .in2(N__19180),
            .in3(N__17748),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI69BV2_6_LC_8_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI69BV2_6_LC_8_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI69BV2_6_LC_8_25_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI69BV2_6_LC_8_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16383),
            .in3(N__17916),
            .lcout(\ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPSC01_6_LC_8_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPSC01_6_LC_8_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPSC01_6_LC_8_25_6 .LUT_INIT=16'b1001101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPSC01_6_LC_8_25_6  (
            .in0(N__19170),
            .in1(N__21061),
            .in2(N__17813),
            .in3(N__19822),
            .lcout(\ppm_encoder_1.N_253_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_8_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_8_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_8_25_7 .LUT_INIT=16'b1011111101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_8_25_7  (
            .in0(N__21063),
            .in1(N__17802),
            .in2(N__19632),
            .in3(N__17304),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIKON03_13_LC_8_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIKON03_13_LC_8_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIKON03_13_LC_8_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIKON03_13_LC_8_26_1  (
            .in0(_gnd_net_),
            .in1(N__18131),
            .in2(_gnd_net_),
            .in3(N__16530),
            .lcout(\ppm_encoder_1.init_pulses_RNIKON03Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_8_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_8_26_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_8_26_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_8_26_2  (
            .in0(N__16786),
            .in1(N__18111),
            .in2(N__16878),
            .in3(N__16518),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23804),
            .ce(),
            .sr(N__23379));
    defparam \ppm_encoder_1.init_pulses_17_LC_8_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_26_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_26_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_8_26_3  (
            .in0(N__16863),
            .in1(N__16789),
            .in2(N__18354),
            .in3(N__16509),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23804),
            .ce(),
            .sr(N__23379));
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_8_26_4  (
            .in0(N__16788),
            .in1(N__18336),
            .in2(N__16880),
            .in3(N__16503),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23804),
            .ce(),
            .sr(N__23379));
    defparam \ppm_encoder_1.init_pulses_1_LC_8_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_8_26_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_8_26_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_8_26_5  (
            .in0(N__18069),
            .in1(N__16790),
            .in2(N__16881),
            .in3(N__16497),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23804),
            .ce(),
            .sr(N__23379));
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_8_26_6  (
            .in0(N__16787),
            .in1(N__18378),
            .in2(N__16879),
            .in3(N__16485),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23804),
            .ce(),
            .sr(N__23379));
    defparam \ppm_encoder_1.init_pulses_RNISPS41_15_LC_8_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISPS41_15_LC_8_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISPS41_15_LC_8_26_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISPS41_15_LC_8_26_7  (
            .in0(N__19746),
            .in1(N__20342),
            .in2(N__21817),
            .in3(N__21145),
            .lcout(\ppm_encoder_1.N_245_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_8_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_8_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIF6081_9_LC_8_27_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIF6081_9_LC_8_27_0  (
            .in0(N__21211),
            .in1(N__24147),
            .in2(N__19765),
            .in3(N__20343),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_8_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_8_27_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_8_27_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_8_27_1  (
            .in0(N__16782),
            .in1(N__18213),
            .in2(N__16877),
            .in3(N__16461),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23797),
            .ce(),
            .sr(N__23385));
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_27_2 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_27_2  (
            .in0(N__21212),
            .in1(N__22512),
            .in2(N__19766),
            .in3(N__20344),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_8_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_27_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_27_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_8_27_3  (
            .in0(N__16780),
            .in1(N__16596),
            .in2(N__16875),
            .in3(N__18198),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23797),
            .ce(),
            .sr(N__23385));
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_27_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_27_4  (
            .in0(N__21213),
            .in1(N__20014),
            .in2(N__19767),
            .in3(N__20345),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_11_LC_8_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_8_27_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_8_27_5 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_8_27_5  (
            .in0(N__18180),
            .in1(N__16853),
            .in2(N__16800),
            .in3(N__16587),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23797),
            .ce(),
            .sr(N__23385));
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_0_12_LC_8_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_0_12_LC_8_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_0_12_LC_8_27_6 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPMS41_0_12_LC_8_27_6  (
            .in0(N__21214),
            .in1(N__19318),
            .in2(N__19768),
            .in3(N__20346),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_12_LC_8_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_8_27_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_8_27_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_8_27_7  (
            .in0(N__16781),
            .in1(N__18165),
            .in2(N__16876),
            .in3(N__16578),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23797),
            .ce(),
            .sr(N__23385));
    defparam \ppm_encoder_1.init_pulses_2_LC_8_28_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_8_28_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_8_28_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_8_28_0  (
            .in0(N__16794),
            .in1(N__18018),
            .in2(N__16919),
            .in3(N__16569),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam \ppm_encoder_1.init_pulses_3_LC_8_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_8_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_8_28_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_8_28_1  (
            .in0(N__16910),
            .in1(N__17997),
            .in2(N__16557),
            .in3(N__16799),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam \ppm_encoder_1.init_pulses_5_LC_8_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_8_28_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_8_28_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_8_28_2  (
            .in0(N__16795),
            .in1(N__17952),
            .in2(N__16920),
            .in3(N__16542),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam \ppm_encoder_1.init_pulses_6_LC_8_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_8_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_8_28_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_8_28_3  (
            .in0(N__17895),
            .in1(N__16797),
            .in2(N__16922),
            .in3(N__16947),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam \ppm_encoder_1.init_pulses_7_LC_8_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_8_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_8_28_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_8_28_4  (
            .in0(N__16796),
            .in1(N__18243),
            .in2(N__16921),
            .in3(N__16935),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam \ppm_encoder_1.init_pulses_8_LC_8_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_8_28_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_8_28_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_8_28_5  (
            .in0(N__16914),
            .in1(N__16798),
            .in2(N__18231),
            .in3(N__16722),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23792),
            .ce(),
            .sr(N__23393));
    defparam CONSTANT_ONE_LUT4_LC_9_19_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_19_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_8_LC_9_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_9_21_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_9_21_2  (
            .in0(N__16710),
            .in1(N__16698),
            .in2(N__18555),
            .in3(N__17459),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23827),
            .ce(),
            .sr(N__23357));
    defparam \ppm_encoder_1.throttle_7_LC_9_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_9_21_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_9_21_5  (
            .in0(N__16674),
            .in1(N__16656),
            .in2(N__17509),
            .in3(N__18534),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23827),
            .ce(),
            .sr(N__23357));
    defparam \ppm_encoder_1.rudder_7_LC_9_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_9_21_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_9_21_6  (
            .in0(N__16638),
            .in1(N__16623),
            .in2(N__22283),
            .in3(N__17458),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23827),
            .ce(),
            .sr(N__23357));
    defparam \ppm_encoder_1.rudder_RNITHN71_7_LC_9_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNITHN71_7_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNITHN71_7_LC_9_22_0 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \ppm_encoder_1.rudder_RNITHN71_7_LC_9_22_0  (
            .in0(N__19552),
            .in1(N__18739),
            .in2(N__22279),
            .in3(N__18901),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5QED3_7_LC_9_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5QED3_7_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5QED3_7_LC_9_22_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5QED3_7_LC_9_22_1  (
            .in0(N__18512),
            .in1(_gnd_net_),
            .in2(N__16599),
            .in3(N__17133),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_0_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJ7DC5_7_LC_9_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJ7DC5_7_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJ7DC5_7_LC_9_22_2 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJ7DC5_7_LC_9_22_2  (
            .in0(N__19467),
            .in1(N__17703),
            .in2(N__17202),
            .in3(N__17029),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFL141_7_LC_9_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFL141_7_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFL141_7_LC_9_22_4 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIFL141_7_LC_9_22_4  (
            .in0(N__17184),
            .in1(N__17087),
            .in2(N__17151),
            .in3(N__17872),
            .lcout(\ppm_encoder_1.pulses2count_9_i_o2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIPIL11_7_LC_9_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIPIL11_7_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIPIL11_7_LC_9_22_5 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \ppm_encoder_1.throttle_RNIPIL11_7_LC_9_22_5  (
            .in0(N__18532),
            .in1(N__22269),
            .in2(_gnd_net_),
            .in3(N__19551),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_rn_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_9_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_9_22_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_9_22_6  (
            .in0(N__17127),
            .in1(N__17112),
            .in2(N__17535),
            .in3(N__17088),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23822),
            .ce(),
            .sr(N__23361));
    defparam \ppm_encoder_1.init_pulses_RNI4LRJ2_1_LC_9_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI4LRJ2_1_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4LRJ2_1_LC_9_23_0 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4LRJ2_1_LC_9_23_0  (
            .in0(N__17067),
            .in1(N__17306),
            .in2(N__17704),
            .in3(N__17027),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOC8K3_1_LC_9_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOC8K3_1_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOC8K3_1_LC_9_23_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOC8K3_1_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17079),
            .in3(N__17276),
            .lcout(\ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNISDTK_1_LC_9_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNISDTK_1_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNISDTK_1_LC_9_23_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.throttle_RNISDTK_1_LC_9_23_2  (
            .in0(N__20770),
            .in1(N__18735),
            .in2(_gnd_net_),
            .in3(N__18899),
            .lcout(\ppm_encoder_1.N_426 ),
            .ltout(\ppm_encoder_1.N_426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI6NRJ2_3_LC_9_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI6NRJ2_3_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI6NRJ2_3_LC_9_23_3 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI6NRJ2_3_LC_9_23_3  (
            .in0(N__17028),
            .in1(N__20586),
            .in2(N__16962),
            .in3(N__17666),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISG8K3_3_LC_9_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISG8K3_3_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISG8K3_3_LC_9_23_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISG8K3_3_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16959),
            .in3(N__17258),
            .lcout(\ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_1_LC_9_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_9_23_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__17563),
            .in2(_gnd_net_),
            .in3(N__20771),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23817),
            .ce(),
            .sr(N__23365));
    defparam \ppm_encoder_1.init_pulses_RNIKNC01_1_LC_9_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIKNC01_1_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIKNC01_1_LC_9_23_6 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIKNC01_1_LC_9_23_6  (
            .in0(N__17803),
            .in1(N__19820),
            .in2(N__21130),
            .in3(N__17305),
            .lcout(\ppm_encoder_1.N_248_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIMPC01_3_LC_9_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIMPC01_3_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIMPC01_3_LC_9_23_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIMPC01_3_LC_9_23_7  (
            .in0(N__19821),
            .in1(N__17804),
            .in2(N__20591),
            .in3(N__21060),
            .lcout(\ppm_encoder_1.N_250_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIB4081_7_LC_9_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIB4081_7_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIB4081_7_LC_9_24_0 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIB4081_7_LC_9_24_0  (
            .in0(N__21085),
            .in1(N__19593),
            .in2(N__19475),
            .in3(N__17811),
            .lcout(\ppm_encoder_1.N_254_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_9_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_9_24_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19425),
            .in3(N__22835),
            .lcout(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0 ),
            .ltout(\ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIE6081_9_LC_9_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIE6081_9_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIE6081_9_LC_9_24_2 .LUT_INIT=16'b1010011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIE6081_9_LC_9_24_2  (
            .in0(N__24157),
            .in1(N__19686),
            .in2(N__17223),
            .in3(N__19592),
            .lcout(\ppm_encoder_1.N_246_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17J_3_LC_9_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17J_3_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17J_3_LC_9_24_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17J_3_LC_9_24_3  (
            .in0(N__19858),
            .in1(N__19816),
            .in2(N__24405),
            .in3(N__22836),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_9_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_9_24_4 .LUT_INIT=16'b0101000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_9_24_4  (
            .in0(N__23506),
            .in1(N__18640),
            .in2(N__19866),
            .in3(N__21204),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_9_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_9_24_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_9_24_5  (
            .in0(N__21202),
            .in1(N__23507),
            .in2(N__18290),
            .in3(N__19817),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_9_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_9_24_6 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_9_24_6  (
            .in0(N__21973),
            .in1(N__17871),
            .in2(N__23531),
            .in3(N__21203),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIMKS41_10_LC_9_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIMKS41_10_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIMKS41_10_LC_9_24_7 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIMKS41_10_LC_9_24_7  (
            .in0(N__19591),
            .in1(N__22525),
            .in2(N__19706),
            .in3(N__21084),
            .lcout(\ppm_encoder_1.N_256_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_9_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI70081_3_LC_9_25_0 .LUT_INIT=16'b1100011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI70081_3_LC_9_25_0  (
            .in0(N__17812),
            .in1(N__20587),
            .in2(N__21169),
            .in3(N__19630),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_9_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_9_25_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_9_25_1  (
            .in0(N__21772),
            .in1(N__24004),
            .in2(N__21271),
            .in3(N__21099),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI98UU1_2_LC_9_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98UU1_2_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98UU1_2_LC_9_25_2 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98UU1_2_LC_9_25_2  (
            .in0(N__20532),
            .in1(N__17744),
            .in2(N__21168),
            .in3(N__17667),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGLA33_2_LC_9_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGLA33_2_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGLA33_2_LC_9_25_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGLA33_2_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17586),
            .in3(N__18039),
            .lcout(\ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIROS41_14_LC_9_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIROS41_14_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIROS41_14_LC_9_25_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIROS41_14_LC_9_25_4  (
            .in0(N__21097),
            .in1(N__21507),
            .in2(N__19714),
            .in3(N__20391),
            .lcout(\ppm_encoder_1.N_260_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_9_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA2081_5_LC_9_25_5 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA2081_5_LC_9_25_5  (
            .in0(N__19631),
            .in1(N__19701),
            .in2(N__22577),
            .in3(N__21098),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI4RFR_0_LC_9_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI4RFR_0_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI4RFR_0_LC_9_25_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_RNI4RFR_0_LC_9_25_6  (
            .in0(N__19862),
            .in1(N__19818),
            .in2(N__20539),
            .in3(N__19424),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7DC41_2_LC_9_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7DC41_2_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7DC41_2_LC_9_25_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7DC41_2_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__20531),
            .in2(N__18090),
            .in3(N__22837),
            .lcout(\ppm_encoder_1.N_249_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUUR33_0_LC_9_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIUUR33_0_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUUR33_0_LC_9_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUUR33_0_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__18087),
            .in2(N__20440),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_9_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__18075),
            .in2(_gnd_net_),
            .in3(N__18063),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_9_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_9_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__18060),
            .in2(N__18047),
            .in3(N__18006),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_9_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_9_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(N__18003),
            .in2(_gnd_net_),
            .in3(N__17988),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_9_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_9_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(N__17985),
            .in2(_gnd_net_),
            .in3(N__17961),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_9_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_9_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(N__17958),
            .in2(_gnd_net_),
            .in3(N__17943),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_9_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_9_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__17940),
            .in2(N__17929),
            .in3(N__17886),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_9_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_9_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__19431),
            .in2(_gnd_net_),
            .in3(N__18234),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_9_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_9_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__18666),
            .in2(_gnd_net_),
            .in3(N__18222),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_9_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_9_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__18219),
            .in2(_gnd_net_),
            .in3(N__18207),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_9_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_9_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__18204),
            .in2(_gnd_net_),
            .in3(N__18192),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_9_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_9_27_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18189),
            .in3(N__18174),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_9_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_9_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__18171),
            .in2(_gnd_net_),
            .in3(N__18159),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_9_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_9_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__18152),
            .in2(N__18120),
            .in3(N__18105),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_LUT4_0_LC_9_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_LUT4_0_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_LUT4_0_LC_9_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_LUT4_0_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18317),
            .in3(N__18093),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_9_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_9_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__20625),
            .in2(_gnd_net_),
            .in3(N__18372),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_9_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_9_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__18327),
            .in2(_gnd_net_),
            .in3(N__18357),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_9_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_9_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__18300),
            .in2(_gnd_net_),
            .in3(N__18342),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_9_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_9_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__19968),
            .in2(_gnd_net_),
            .in3(N__18339),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_28_3 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_28_3  (
            .in0(N__21218),
            .in1(N__23522),
            .in2(N__18273),
            .in3(N__23961),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23788),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_9_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVM131_16_LC_9_28_5 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVM131_16_LC_9_28_5  (
            .in0(N__21216),
            .in1(N__23959),
            .in2(N__21272),
            .in3(N__21685),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_28_6 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_28_6  (
            .in0(N__21684),
            .in1(N__21511),
            .in2(N__24002),
            .in3(N__21215),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_9_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0O131_17_LC_9_28_7 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0O131_17_LC_9_28_7  (
            .in0(N__21217),
            .in1(N__23960),
            .in2(N__20926),
            .in3(N__21686),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_0_0_LC_9_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_0_0_LC_9_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_0_0_LC_9_29_2 .LUT_INIT=16'b0000011110001000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_0_0_LC_9_29_2  (
            .in0(N__22097),
            .in1(N__21965),
            .in2(N__21734),
            .in3(N__20396),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_9_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_9_29_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_9_29_6 .LUT_INIT=16'b1111011100001111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_9_29_6  (
            .in0(N__22096),
            .in1(N__21964),
            .in2(N__21733),
            .in3(N__20395),
            .lcout(\ppm_encoder_1.N_204 ),
            .ltout(\ppm_encoder_1.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_9_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_9_29_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_9_29_7 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_9_29_7  (
            .in0(N__23511),
            .in1(N__21702),
            .in2(N__18597),
            .in3(N__21219),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23785),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_0 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_0  (
            .in0(N__18594),
            .in1(N__20159),
            .in2(N__20273),
            .in3(N__18576),
            .lcout(),
            .ltout(\ppm_encoder_1.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_1 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__20419),
            .in2(N__18558),
            .in3(N__18551),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_10_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_10_20_5 .LUT_INIT=16'b1100010111001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_10_20_5  (
            .in0(N__18533),
            .in1(N__18516),
            .in2(N__18789),
            .in3(N__18903),
            .lcout(\ppm_encoder_1.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_10_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_10_20_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_10_20_6  (
            .in0(N__20420),
            .in1(N__18501),
            .in2(N__20274),
            .in3(N__20160),
            .lcout(\ppm_encoder_1.N_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_10_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_10_21_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_10_21_0  (
            .in0(N__22116),
            .in1(N__21975),
            .in2(N__18387),
            .in3(N__18468),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_10_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_10_21_2 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_10_21_2  (
            .in0(N__22117),
            .in1(N__21976),
            .in2(N__18444),
            .in3(N__18435),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_10_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_10_21_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_10_21_7  (
            .in0(N__20158),
            .in1(N__18414),
            .in2(N__20421),
            .in3(N__20272),
            .lcout(\ppm_encoder_1.N_391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_10_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_10_22_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_10_22_0  (
            .in0(N__22118),
            .in1(N__21991),
            .in2(N__19092),
            .in3(N__24025),
            .lcout(\ppm_encoder_1.N_393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIHVID1_1_LC_10_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIHVID1_1_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIHVID1_1_LC_10_22_1 .LUT_INIT=16'b1111101011110100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIHVID1_1_LC_10_22_1  (
            .in0(N__21993),
            .in1(N__20418),
            .in2(N__21786),
            .in3(N__22120),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_22_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_22_2  (
            .in0(N__22119),
            .in1(N__21992),
            .in2(N__19059),
            .in3(N__19047),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_10_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_10_22_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_10_22_3  (
            .in0(N__20257),
            .in1(N__20157),
            .in2(_gnd_net_),
            .in3(N__19014),
            .lcout(),
            .ltout(\ppm_encoder_1.N_327_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_10_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_10_22_4 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_10_22_4  (
            .in0(N__18984),
            .in1(N__24024),
            .in2(N__18972),
            .in3(N__18969),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_10_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_10_22_6 .LUT_INIT=16'b1100110001011100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_10_22_6  (
            .in0(N__18939),
            .in1(N__18921),
            .in2(N__18900),
            .in3(N__18787),
            .lcout(\ppm_encoder_1.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNID5081_0_8_LC_10_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID5081_0_8_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID5081_0_8_LC_10_23_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID5081_0_8_LC_10_23_0  (
            .in0(N__19690),
            .in1(N__19623),
            .in2(N__22703),
            .in3(N__21089),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_10_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_10_23_1 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_10_23_1  (
            .in0(N__21090),
            .in1(N__23520),
            .in2(N__18653),
            .in3(N__19691),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23805),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNID5081_8_LC_10_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID5081_8_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID5081_8_LC_10_23_2 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID5081_8_LC_10_23_2  (
            .in0(N__19688),
            .in1(N__19622),
            .in2(N__22702),
            .in3(N__21087),
            .lcout(\ppm_encoder_1.N_255_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_10_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_10_23_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_10_23_3  (
            .in0(N__20828),
            .in1(N__19336),
            .in2(N__24253),
            .in3(N__19374),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_10_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_10_23_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_10_23_4  (
            .in0(N__19689),
            .in1(N__20407),
            .in2(N__19338),
            .in3(N__21088),
            .lcout(\ppm_encoder_1.N_258_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_10_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_10_23_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_10_23_6  (
            .in0(N__19687),
            .in1(N__20406),
            .in2(N__20039),
            .in3(N__21086),
            .lcout(\ppm_encoder_1.N_257_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_10_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_10_23_7 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_10_23_7  (
            .in0(N__20408),
            .in1(N__21781),
            .in2(N__21609),
            .in3(N__19239),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_10_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_10_24_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_10_24_0  (
            .in0(N__19143),
            .in1(N__22384),
            .in2(N__19128),
            .in3(N__22327),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_10_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_10_24_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_10_24_1  (
            .in0(N__19209),
            .in1(N__19203),
            .in2(N__19188),
            .in3(N__24236),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23799),
            .ce(N__23569),
            .sr(N__23371));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_10_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_10_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_10_24_2 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_10_24_2  (
            .in0(N__24235),
            .in1(N__19137),
            .in2(N__22251),
            .in3(N__19471),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23799),
            .ce(N__23569),
            .sr(N__23371));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_10_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_10_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_10_24_5  (
            .in0(N__21407),
            .in1(N__19119),
            .in2(N__19113),
            .in3(N__19101),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23799),
            .ce(N__23569),
            .sr(N__23371));
    defparam \ppm_encoder_1.init_pulses_RNILB4M_0_LC_10_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILB4M_0_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILB4M_0_LC_10_25_0 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILB4M_0_LC_10_25_0  (
            .in0(N__24393),
            .in1(N__19861),
            .in2(N__22235),
            .in3(N__19819),
            .lcout(\ppm_encoder_1.init_pulses_RNILB4MZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC4081_7_LC_10_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC4081_7_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC4081_7_LC_10_25_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC4081_7_LC_10_25_1  (
            .in0(N__19705),
            .in1(N__19621),
            .in2(N__19479),
            .in3(N__21100),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_10_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_fast_0_LC_10_25_2 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_0_LC_10_25_2  (
            .in0(N__22840),
            .in1(N__24529),
            .in2(N__22872),
            .in3(N__24579),
            .lcout(\ppm_encoder_1.PPM_STATE_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23794),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNII3AF_1_LC_10_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNII3AF_1_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNII3AF_1_LC_10_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNII3AF_1_LC_10_25_3  (
            .in0(N__24345),
            .in1(N__22186),
            .in2(N__22469),
            .in3(N__22839),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_10_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_10_25_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ppm_encoder_1.counter_RNIS9KG_2_LC_10_25_4  (
            .in0(N__20753),
            .in1(N__20732),
            .in2(N__22770),
            .in3(N__22733),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_10_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_10_25_5 .LUT_INIT=16'b0000101000001011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_10_25_5  (
            .in0(N__24578),
            .in1(N__22868),
            .in2(N__24534),
            .in3(N__22841),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23794),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_10_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_10_25_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_10_25_6  (
            .in0(N__24394),
            .in1(N__24528),
            .in2(_gnd_net_),
            .in3(N__24577),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23794),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_10_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_10_26_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_10_26_1  (
            .in0(N__24346),
            .in1(N__22194),
            .in2(N__22470),
            .in3(N__24401),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_10_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_10_26_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_10_26_2  (
            .in0(N__22072),
            .in1(N__21942),
            .in2(N__24086),
            .in3(N__19410),
            .lcout(\ppm_encoder_1.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_LC_10_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIMR0V_0_LC_10_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIMR0V_0_LC_10_26_4  (
            .in0(N__22231),
            .in1(N__20466),
            .in2(_gnd_net_),
            .in3(N__22838),
            .lcout(\ppm_encoder_1.N_247_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNI1UMR_LC_10_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNI1UMR_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNI1UMR_LC_10_26_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNI1UMR_LC_10_26_5  (
            .in0(N__20414),
            .in1(N__20255),
            .in2(_gnd_net_),
            .in3(N__20143),
            .lcout(\ppm_encoder_1.N_441 ),
            .ltout(\ppm_encoder_1.N_441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_10_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_10_26_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_10_26_6  (
            .in0(N__20816),
            .in1(N__20032),
            .in2(N__19995),
            .in3(N__19992),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIM3KG_18_LC_10_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIM3KG_18_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIM3KG_18_LC_10_26_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ppm_encoder_1.counter_RNIM3KG_18_LC_10_26_7  (
            .in0(N__21450),
            .in1(N__22990),
            .in2(N__22428),
            .in3(N__22155),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_3_18_LC_10_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_3_18_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_3_18_LC_10_27_0 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_3_18_LC_10_27_0  (
            .in0(N__21761),
            .in1(N__20885),
            .in2(N__24005),
            .in3(N__21221),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_27_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_27_1  (
            .in0(N__22059),
            .in1(N__21980),
            .in2(_gnd_net_),
            .in3(N__19962),
            .lcout(),
            .ltout(\ppm_encoder_1.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_10_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_10_27_2 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_10_27_2  (
            .in0(N__19932),
            .in1(N__19902),
            .in2(N__19890),
            .in3(N__23981),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_10_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_10_27_3 .LUT_INIT=16'b0010000100110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_10_27_3  (
            .in0(N__21222),
            .in1(N__23521),
            .in2(N__22098),
            .in3(N__21981),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23786),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_10_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_10_27_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_10_27_5  (
            .in0(N__22058),
            .in1(N__21979),
            .in2(_gnd_net_),
            .in3(N__19887),
            .lcout(),
            .ltout(\ppm_encoder_1.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_27_6 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_27_6  (
            .in0(N__20700),
            .in1(N__23980),
            .in2(N__20688),
            .in3(N__20685),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_10_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_10_27_7 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_10_27_7  (
            .in0(N__23982),
            .in1(N__21762),
            .in2(N__21621),
            .in3(N__20664),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_0_1_LC_10_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_0_1_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_0_1_LC_10_28_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_0_1_LC_10_28_1  (
            .in0(N__21703),
            .in1(N__22068),
            .in2(N__24003),
            .in3(N__21966),
            .lcout(\ppm_encoder_1.N_247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_10_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUL131_15_LC_10_28_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUL131_15_LC_10_28_4  (
            .in0(N__21687),
            .in1(N__23962),
            .in2(N__21830),
            .in3(N__21220),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_11_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_11_21_4 .LUT_INIT=16'b0000001000000110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_11_21_4  (
            .in0(N__22123),
            .in1(N__21977),
            .in2(N__24085),
            .in3(N__20619),
            .lcout(\ppm_encoder_1.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_22_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_11_22_1  (
            .in0(N__20472),
            .in1(N__24255),
            .in2(N__20502),
            .in3(N__20592),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23806),
            .ce(N__23564),
            .sr(N__23366));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_11_23_1 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_11_23_1  (
            .in0(N__20556),
            .in1(N__24260),
            .in2(N__20547),
            .in3(N__20501),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23800),
            .ce(N__23567),
            .sr(N__23372));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_23_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_23_2  (
            .in0(N__20731),
            .in1(N__20487),
            .in2(N__20481),
            .in3(N__20752),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_23_5 .LUT_INIT=16'b0000011000000010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_23_5  (
            .in0(N__22124),
            .in1(N__21978),
            .in2(N__24089),
            .in3(N__20777),
            .lcout(\ppm_encoder_1.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_23_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_11_23_7  (
            .in0(N__21408),
            .in1(N__20829),
            .in2(N__20793),
            .in3(N__20778),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23800),
            .ce(N__23567),
            .sr(N__23372));
    defparam \ppm_encoder_1.counter_0_LC_11_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_11_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__22154),
            .in2(N__21227),
            .in3(N__21201),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_1_LC_11_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_11_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__22187),
            .in2(_gnd_net_),
            .in3(N__20757),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_2_LC_11_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_11_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_11_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__20754),
            .in2(_gnd_net_),
            .in3(N__20736),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_3_LC_11_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_11_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__20733),
            .in2(_gnd_net_),
            .in3(N__20715),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_4_LC_11_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_11_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__21449),
            .in2(_gnd_net_),
            .in3(N__20712),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_5_LC_11_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_11_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__22368),
            .in2(_gnd_net_),
            .in3(N__20709),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_6_LC_11_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_11_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__22329),
            .in2(_gnd_net_),
            .in3(N__20706),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_7_LC_11_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_11_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__22386),
            .in2(_gnd_net_),
            .in3(N__20703),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__23795),
            .ce(),
            .sr(N__21423));
    defparam \ppm_encoder_1.counter_8_LC_11_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_11_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__24299),
            .in2(_gnd_net_),
            .in3(N__20856),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_9_LC_11_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_11_25_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_11_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_11_25_1  (
            .in0(_gnd_net_),
            .in1(N__24347),
            .in2(_gnd_net_),
            .in3(N__20853),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_10_LC_11_25_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_11_25_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_11_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(N__22427),
            .in2(_gnd_net_),
            .in3(N__20850),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_11_LC_11_25_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_11_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(N__22468),
            .in2(_gnd_net_),
            .in3(N__20847),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_12_LC_11_25_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_11_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__23019),
            .in2(_gnd_net_),
            .in3(N__20844),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_13_LC_11_25_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_11_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(N__22938),
            .in2(_gnd_net_),
            .in3(N__20841),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_14_LC_11_25_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_11_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_11_25_6  (
            .in0(_gnd_net_),
            .in1(N__22349),
            .in2(_gnd_net_),
            .in3(N__20838),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_15_LC_11_25_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_11_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__22968),
            .in2(_gnd_net_),
            .in3(N__20835),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__23790),
            .ce(),
            .sr(N__21422));
    defparam \ppm_encoder_1.counter_16_LC_11_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_11_26_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_11_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_11_26_0  (
            .in0(_gnd_net_),
            .in1(N__22734),
            .in2(_gnd_net_),
            .in3(N__20832),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__23787),
            .ce(),
            .sr(N__21421));
    defparam \ppm_encoder_1.counter_17_LC_11_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_11_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__22766),
            .in2(_gnd_net_),
            .in3(N__21429),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__23787),
            .ce(),
            .sr(N__21421));
    defparam \ppm_encoder_1.counter_18_LC_11_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_11_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_11_26_2  (
            .in0(_gnd_net_),
            .in1(N__22994),
            .in2(_gnd_net_),
            .in3(N__21426),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23787),
            .ce(),
            .sr(N__21421));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_11_27_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_11_27_4  (
            .in0(N__21394),
            .in1(N__21381),
            .in2(N__21375),
            .in3(N__21366),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23784),
            .ce(N__23570),
            .sr(N__23396));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_27_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_27_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_11_27_5  (
            .in0(N__24225),
            .in1(N__21350),
            .in2(N__21303),
            .in3(N__21294),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23784),
            .ce(N__23570),
            .sr(N__23396));
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_28_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_11_28_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_16_LC_11_28_7  (
            .in0(N__24017),
            .in1(N__21622),
            .in2(N__21276),
            .in3(N__21760),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23782),
            .ce(N__23571),
            .sr(N__23401));
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_LC_12_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_LC_12_12_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__23490),
            .in2(_gnd_net_),
            .in3(N__21234),
            .lcout(\ppm_encoder_1.N_238_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_12_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_12_22_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_17_LC_12_22_2  (
            .in0(N__24068),
            .in1(N__20930),
            .in2(N__21624),
            .in3(N__21777),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23798),
            .ce(N__23562),
            .sr(N__23373));
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_12_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_12_22_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_18_LC_12_22_3  (
            .in0(N__21776),
            .in1(N__21614),
            .in2(N__20889),
            .in3(N__24069),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23798),
            .ce(N__23562),
            .sr(N__23373));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_12_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_12_22_6 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_12_22_6  (
            .in0(N__24067),
            .in1(N__21775),
            .in2(N__21623),
            .in3(N__22311),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_22_7 .LUT_INIT=16'b1110111010101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_22_7  (
            .in0(N__21774),
            .in1(N__24066),
            .in2(N__22287),
            .in3(N__21610),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_12_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_12_23_0 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_12_23_0  (
            .in0(N__21989),
            .in1(N__24073),
            .in2(N__22133),
            .in3(N__22236),
            .lcout(\ppm_encoder_1.pulses2count_9_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_12_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_12_23_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_12_23_2  (
            .in0(N__22185),
            .in1(N__23889),
            .in2(N__22164),
            .in3(N__22150),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_1_LC_12_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_1_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_1_LC_12_23_3 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_1_LC_12_23_3  (
            .in0(N__21778),
            .in1(N__22125),
            .in2(N__24087),
            .in3(N__21990),
            .lcout(\ppm_encoder_1.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_12_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_12_23_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_15_LC_12_23_4  (
            .in0(N__21619),
            .in1(N__21780),
            .in2(N__21831),
            .in3(N__24077),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23793),
            .ce(N__23563),
            .sr(N__23380));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_23_5 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_23_5  (
            .in0(N__21779),
            .in1(N__21618),
            .in2(N__24088),
            .in3(N__21539),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_12_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_12_23_6 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_12_23_6  (
            .in0(N__21513),
            .in1(N__24261),
            .in2(N__21471),
            .in3(N__21468),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23793),
            .ce(N__23563),
            .sr(N__23380));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_12_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_12_24_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_12_24_0  (
            .in0(N__22366),
            .in1(N__22608),
            .in2(N__22539),
            .in3(N__21445),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_12_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_12_24_1 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_12_24_1  (
            .in0(N__22656),
            .in1(N__24259),
            .in2(N__24125),
            .in3(N__22644),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23789),
            .ce(N__23566),
            .sr(N__23386));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_12_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_12_24_2 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_12_24_2  (
            .in0(N__24257),
            .in1(N__22602),
            .in2(N__22590),
            .in3(N__22578),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23789),
            .ce(N__23566),
            .sr(N__23386));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_12_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_12_24_3 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_12_24_3  (
            .in0(N__24118),
            .in1(N__24258),
            .in2(N__22530),
            .in3(N__22488),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23789),
            .ce(N__23566),
            .sr(N__23386));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_12_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_12_24_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_12_24_4  (
            .in0(N__22476),
            .in1(N__22461),
            .in2(N__22440),
            .in3(N__22423),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_12_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_12_25_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_12_25_0  (
            .in0(N__24554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24407),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_25_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_25_1  (
            .in0(N__22966),
            .in1(N__22407),
            .in2(N__22398),
            .in3(N__22345),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIGV08_5_LC_12_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIGV08_5_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIGV08_5_LC_12_25_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIGV08_5_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__22385),
            .in2(_gnd_net_),
            .in3(N__22367),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUBKG_6_LC_12_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUBKG_6_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUBKG_6_LC_12_25_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUBKG_6_LC_12_25_3  (
            .in0(N__23018),
            .in1(N__24298),
            .in2(N__22350),
            .in3(N__22328),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4 ),
            .ltout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI09RH2_1_LC_12_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI09RH2_1_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI09RH2_1_LC_12_25_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNI09RH2_1_LC_12_25_4  (
            .in0(N__22895),
            .in1(N__23055),
            .in2(N__23046),
            .in3(N__22920),
            .lcout(\ppm_encoder_1.N_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_12_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_12_25_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_12_25_6  (
            .in0(N__23043),
            .in1(N__22936),
            .in2(N__23031),
            .in3(N__23017),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_12_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_12_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_12_25_7  (
            .in0(_gnd_net_),
            .in1(N__23004),
            .in2(_gnd_net_),
            .in3(N__22995),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIKF811_13_LC_12_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIKF811_13_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIKF811_13_LC_12_26_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIKF811_13_LC_12_26_2  (
            .in0(N__22974),
            .in1(N__22967),
            .in2(N__22950),
            .in3(N__22937),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2 ),
            .ltout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_26_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_26_3  (
            .in0(N__22914),
            .in1(N__22905),
            .in2(N__22899),
            .in3(N__22896),
            .lcout(),
            .ltout(\ppm_encoder_1.N_431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_26_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_26_4 .LUT_INIT=16'b1010001110101011;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_12_26_4  (
            .in0(N__22787),
            .in1(N__22862),
            .in2(N__22851),
            .in3(N__22848),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23783),
            .ce(),
            .sr(N__23397));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_12_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_12_27_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_12_27_5  (
            .in0(N__22776),
            .in1(N__22762),
            .in2(N__22746),
            .in3(N__22732),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_13_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_13_22_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_13_22_0 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_13_22_0  (
            .in0(N__24254),
            .in1(N__22716),
            .in2(N__24126),
            .in3(N__22704),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23807),
            .ce(N__23565),
            .sr(N__23381));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_13_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_13_23_2 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_13_23_2  (
            .in0(N__24273),
            .in1(N__24256),
            .in2(N__24165),
            .in3(N__24117),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23801),
            .ce(N__23568),
            .sr(N__23387));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_13_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_13_23_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_13_23_3  (
            .in0(N__24116),
            .in1(N__24096),
            .in2(_gnd_net_),
            .in3(N__24078),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23801),
            .ce(N__23568),
            .sr(N__23387));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_13_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_13_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__23094),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_13_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_13_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__23088),
            .in2(N__24747),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_13_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_13_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__23076),
            .in2(N__24741),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_13_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_13_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__23070),
            .in2(N__24744),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_13_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_13_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__24279),
            .in2(N__24742),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_13_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_13_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__23061),
            .in2(N__24745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_13_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_13_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__24801),
            .in2(N__24743),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_13_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_13_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__24795),
            .in2(N__24746),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_13_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_13_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__24712),
            .in2(N__24789),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_13_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_13_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__24777),
            .in2(N__24748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_13_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_13_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24582),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_25_5 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_25_5  (
            .in0(N__24569),
            .in1(N__24550),
            .in2(N__24533),
            .in3(N__24406),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_13_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_13_25_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_13_25_6  (
            .in0(N__24348),
            .in1(N__24321),
            .in2(N__24312),
            .in3(N__24300),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // Pc2Drone
