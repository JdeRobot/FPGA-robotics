//---- Felipe Machado -------------------------------
//---- Area de Tecnologia Electronica ---------------
//---- Universidad Rey Juan Carlos ------------------
//---- https://github.com/felipe-m ------------------
//---------------------------------------------------
//---- Autcmatically generated verilog ROM blockfrom a VHDL file----
//  Original VHDL file name: rom_red_square_80x60_rgb_9b.vhd
//  Constant VHDL name: filaimg
//  Memory with non-blocking assignments (<=)

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module rom_red_square_80x60_rgb_9b
  (
     input     clk,   // clock
     input      [13-1:0] addr,  //4800 memory positions
     output reg  [9-1:0] filaimg  // memory data width
  );


//  Memory with clock

  always @(posedge clk)
  begin
    case(addr)
            //"RRRGGGBBB"
      13'h0: filaimg <= 9'b101110110;
      13'h1: filaimg <= 9'b101110110;
      13'h2: filaimg <= 9'b101110110;
      13'h3: filaimg <= 9'b101110110;
      13'h4: filaimg <= 9'b101110110;
      13'h5: filaimg <= 9'b101110110;
      13'h6: filaimg <= 9'b101110110;
      13'h7: filaimg <= 9'b101110110;
      13'h8: filaimg <= 9'b101110110;
      13'h9: filaimg <= 9'b101110110;
      13'hA: filaimg <= 9'b101110110;
      13'hB: filaimg <= 9'b101110110;
      13'hC: filaimg <= 9'b101110110;
      13'hD: filaimg <= 9'b101110110;
      13'hE: filaimg <= 9'b101110110;
      13'hF: filaimg <= 9'b101110110;
      13'h10: filaimg <= 9'b101110110;
      13'h11: filaimg <= 9'b101110110;
      13'h12: filaimg <= 9'b101110110;
      13'h13: filaimg <= 9'b101110110;
      13'h14: filaimg <= 9'b101110110;
      13'h15: filaimg <= 9'b101110110;
      13'h16: filaimg <= 9'b101110110;
      13'h17: filaimg <= 9'b101110110;
      13'h18: filaimg <= 9'b101110110;
      13'h19: filaimg <= 9'b101110110;
      13'h1A: filaimg <= 9'b101110110;
      13'h1B: filaimg <= 9'b101110110;
      13'h1C: filaimg <= 9'b101110110;
      13'h1D: filaimg <= 9'b101110110;
      13'h1E: filaimg <= 9'b101110110;
      13'h1F: filaimg <= 9'b101110110;
      13'h20: filaimg <= 9'b101110110;
      13'h21: filaimg <= 9'b101110110;
      13'h22: filaimg <= 9'b101110110;
      13'h23: filaimg <= 9'b101110110;
      13'h24: filaimg <= 9'b101110110;
      13'h25: filaimg <= 9'b101110110;
      13'h26: filaimg <= 9'b101110110;
      13'h27: filaimg <= 9'b101110110;
      13'h28: filaimg <= 9'b101110110;
      13'h29: filaimg <= 9'b101110110;
      13'h2A: filaimg <= 9'b101110110;
      13'h2B: filaimg <= 9'b101110110;
      13'h2C: filaimg <= 9'b101110110;
      13'h2D: filaimg <= 9'b101110110;
      13'h2E: filaimg <= 9'b101110110;
      13'h2F: filaimg <= 9'b101110110;
      13'h30: filaimg <= 9'b101110110;
      13'h31: filaimg <= 9'b101110110;
      13'h32: filaimg <= 9'b101110110;
      13'h33: filaimg <= 9'b101110110;
      13'h34: filaimg <= 9'b101110110;
      13'h35: filaimg <= 9'b101110110;
      13'h36: filaimg <= 9'b101110110;
      13'h37: filaimg <= 9'b101110110;
      13'h38: filaimg <= 9'b101110110;
      13'h39: filaimg <= 9'b101110110;
      13'h3A: filaimg <= 9'b101110110;
      13'h3B: filaimg <= 9'b101110110;
      13'h3C: filaimg <= 9'b101110110;
      13'h3D: filaimg <= 9'b101110110;
      13'h3E: filaimg <= 9'b101110110;
      13'h3F: filaimg <= 9'b101110110;
      13'h40: filaimg <= 9'b101110110;
      13'h41: filaimg <= 9'b101110110;
      13'h42: filaimg <= 9'b101110110;
      13'h43: filaimg <= 9'b101110110;
      13'h44: filaimg <= 9'b101110110;
      13'h45: filaimg <= 9'b101110110;
      13'h46: filaimg <= 9'b101110110;
      13'h47: filaimg <= 9'b101110110;
      13'h48: filaimg <= 9'b101110110;
      13'h49: filaimg <= 9'b101110110;
      13'h4A: filaimg <= 9'b101110110;
      13'h4B: filaimg <= 9'b101110110;
      13'h4C: filaimg <= 9'b101110110;
      13'h4D: filaimg <= 9'b101110110;
      13'h4E: filaimg <= 9'b101110110;
      13'h4F: filaimg <= 9'b101110110;
      13'h50: filaimg <= 9'b101110110;
      13'h51: filaimg <= 9'b101110110;
      13'h52: filaimg <= 9'b101110110;
      13'h53: filaimg <= 9'b101110110;
      13'h54: filaimg <= 9'b101110110;
      13'h55: filaimg <= 9'b101110110;
      13'h56: filaimg <= 9'b101110110;
      13'h57: filaimg <= 9'b101110110;
      13'h58: filaimg <= 9'b101110110;
      13'h59: filaimg <= 9'b101110110;
      13'h5A: filaimg <= 9'b101110110;
      13'h5B: filaimg <= 9'b101110110;
      13'h5C: filaimg <= 9'b101110110;
      13'h5D: filaimg <= 9'b101110110;
      13'h5E: filaimg <= 9'b101110110;
      13'h5F: filaimg <= 9'b101110110;
      13'h60: filaimg <= 9'b101110110;
      13'h61: filaimg <= 9'b101110110;
      13'h62: filaimg <= 9'b101110110;
      13'h63: filaimg <= 9'b101110110;
      13'h64: filaimg <= 9'b101110110;
      13'h65: filaimg <= 9'b101110110;
      13'h66: filaimg <= 9'b101110110;
      13'h67: filaimg <= 9'b101110110;
      13'h68: filaimg <= 9'b101110110;
      13'h69: filaimg <= 9'b101110110;
      13'h6A: filaimg <= 9'b101110110;
      13'h6B: filaimg <= 9'b101110110;
      13'h6C: filaimg <= 9'b101110110;
      13'h6D: filaimg <= 9'b101110110;
      13'h6E: filaimg <= 9'b101110110;
      13'h6F: filaimg <= 9'b101110110;
      13'h70: filaimg <= 9'b101110110;
      13'h71: filaimg <= 9'b101110110;
      13'h72: filaimg <= 9'b101110110;
      13'h73: filaimg <= 9'b101110110;
      13'h74: filaimg <= 9'b101110110;
      13'h75: filaimg <= 9'b101110110;
      13'h76: filaimg <= 9'b101110110;
      13'h77: filaimg <= 9'b101110110;
      13'h78: filaimg <= 9'b101110110;
      13'h79: filaimg <= 9'b101110110;
      13'h7A: filaimg <= 9'b101110110;
      13'h7B: filaimg <= 9'b101110110;
      13'h7C: filaimg <= 9'b101110110;
      13'h7D: filaimg <= 9'b101110110;
      13'h7E: filaimg <= 9'b101110110;
      13'h7F: filaimg <= 9'b101110110;
      13'h80: filaimg <= 9'b101110110;
      13'h81: filaimg <= 9'b101110110;
      13'h82: filaimg <= 9'b101110110;
      13'h83: filaimg <= 9'b101110110;
      13'h84: filaimg <= 9'b101110110;
      13'h85: filaimg <= 9'b101110110;
      13'h86: filaimg <= 9'b101110110;
      13'h87: filaimg <= 9'b101110110;
      13'h88: filaimg <= 9'b101110110;
      13'h89: filaimg <= 9'b101110110;
      13'h8A: filaimg <= 9'b101110110;
      13'h8B: filaimg <= 9'b101110110;
      13'h8C: filaimg <= 9'b101110110;
      13'h8D: filaimg <= 9'b101110110;
      13'h8E: filaimg <= 9'b101110110;
      13'h8F: filaimg <= 9'b101110110;
      13'h90: filaimg <= 9'b101110110;
      13'h91: filaimg <= 9'b101110110;
      13'h92: filaimg <= 9'b101110110;
      13'h93: filaimg <= 9'b101110110;
      13'h94: filaimg <= 9'b101110110;
      13'h95: filaimg <= 9'b101110110;
      13'h96: filaimg <= 9'b101110110;
      13'h97: filaimg <= 9'b101110110;
      13'h98: filaimg <= 9'b101110110;
      13'h99: filaimg <= 9'b101110110;
      13'h9A: filaimg <= 9'b101110110;
      13'h9B: filaimg <= 9'b101110110;
      13'h9C: filaimg <= 9'b101110110;
      13'h9D: filaimg <= 9'b101110110;
      13'h9E: filaimg <= 9'b101110110;
      13'h9F: filaimg <= 9'b101110110;
      13'hA0: filaimg <= 9'b101110110;
      13'hA1: filaimg <= 9'b101110110;
      13'hA2: filaimg <= 9'b101110110;
      13'hA3: filaimg <= 9'b101110110;
      13'hA4: filaimg <= 9'b101110110;
      13'hA5: filaimg <= 9'b101110110;
      13'hA6: filaimg <= 9'b101110110;
      13'hA7: filaimg <= 9'b101110110;
      13'hA8: filaimg <= 9'b101110110;
      13'hA9: filaimg <= 9'b101110110;
      13'hAA: filaimg <= 9'b101110110;
      13'hAB: filaimg <= 9'b101110110;
      13'hAC: filaimg <= 9'b101110110;
      13'hAD: filaimg <= 9'b101110110;
      13'hAE: filaimg <= 9'b101110110;
      13'hAF: filaimg <= 9'b101110110;
      13'hB0: filaimg <= 9'b101110110;
      13'hB1: filaimg <= 9'b101110110;
      13'hB2: filaimg <= 9'b101110110;
      13'hB3: filaimg <= 9'b101110110;
      13'hB4: filaimg <= 9'b101110110;
      13'hB5: filaimg <= 9'b101110110;
      13'hB6: filaimg <= 9'b101110110;
      13'hB7: filaimg <= 9'b101110110;
      13'hB8: filaimg <= 9'b101110110;
      13'hB9: filaimg <= 9'b101110110;
      13'hBA: filaimg <= 9'b101110110;
      13'hBB: filaimg <= 9'b101110110;
      13'hBC: filaimg <= 9'b101110110;
      13'hBD: filaimg <= 9'b101110110;
      13'hBE: filaimg <= 9'b101110110;
      13'hBF: filaimg <= 9'b101110110;
      13'hC0: filaimg <= 9'b101110110;
      13'hC1: filaimg <= 9'b101110110;
      13'hC2: filaimg <= 9'b101110110;
      13'hC3: filaimg <= 9'b101110110;
      13'hC4: filaimg <= 9'b101110110;
      13'hC5: filaimg <= 9'b101110110;
      13'hC6: filaimg <= 9'b101110110;
      13'hC7: filaimg <= 9'b101110110;
      13'hC8: filaimg <= 9'b101110110;
      13'hC9: filaimg <= 9'b101110110;
      13'hCA: filaimg <= 9'b101110110;
      13'hCB: filaimg <= 9'b101110110;
      13'hCC: filaimg <= 9'b101110110;
      13'hCD: filaimg <= 9'b101110110;
      13'hCE: filaimg <= 9'b101110110;
      13'hCF: filaimg <= 9'b101110110;
      13'hD0: filaimg <= 9'b101110110;
      13'hD1: filaimg <= 9'b101110110;
      13'hD2: filaimg <= 9'b101110110;
      13'hD3: filaimg <= 9'b101110110;
      13'hD4: filaimg <= 9'b101110110;
      13'hD5: filaimg <= 9'b101110110;
      13'hD6: filaimg <= 9'b101110110;
      13'hD7: filaimg <= 9'b101110110;
      13'hD8: filaimg <= 9'b101110110;
      13'hD9: filaimg <= 9'b101110110;
      13'hDA: filaimg <= 9'b101110110;
      13'hDB: filaimg <= 9'b101110110;
      13'hDC: filaimg <= 9'b101110110;
      13'hDD: filaimg <= 9'b101110110;
      13'hDE: filaimg <= 9'b101110110;
      13'hDF: filaimg <= 9'b101110110;
      13'hE0: filaimg <= 9'b101110110;
      13'hE1: filaimg <= 9'b101110110;
      13'hE2: filaimg <= 9'b101110110;
      13'hE3: filaimg <= 9'b101110110;
      13'hE4: filaimg <= 9'b101110110;
      13'hE5: filaimg <= 9'b101110110;
      13'hE6: filaimg <= 9'b101110110;
      13'hE7: filaimg <= 9'b101110110;
      13'hE8: filaimg <= 9'b101110110;
      13'hE9: filaimg <= 9'b101110110;
      13'hEA: filaimg <= 9'b101110110;
      13'hEB: filaimg <= 9'b101110110;
      13'hEC: filaimg <= 9'b101110110;
      13'hED: filaimg <= 9'b101110110;
      13'hEE: filaimg <= 9'b101110110;
      13'hEF: filaimg <= 9'b101110110;
      13'hF0: filaimg <= 9'b101110110;
      13'hF1: filaimg <= 9'b101110110;
      13'hF2: filaimg <= 9'b101110110;
      13'hF3: filaimg <= 9'b101110110;
      13'hF4: filaimg <= 9'b101110110;
      13'hF5: filaimg <= 9'b101110110;
      13'hF6: filaimg <= 9'b101110110;
      13'hF7: filaimg <= 9'b101110110;
      13'hF8: filaimg <= 9'b101110110;
      13'hF9: filaimg <= 9'b101110110;
      13'hFA: filaimg <= 9'b101110110;
      13'hFB: filaimg <= 9'b101110110;
      13'hFC: filaimg <= 9'b101110110;
      13'hFD: filaimg <= 9'b101110110;
      13'hFE: filaimg <= 9'b101110110;
      13'hFF: filaimg <= 9'b101110110;
      13'h100: filaimg <= 9'b101110110;
      13'h101: filaimg <= 9'b101110110;
      13'h102: filaimg <= 9'b101110110;
      13'h103: filaimg <= 9'b101110110;
      13'h104: filaimg <= 9'b101110110;
      13'h105: filaimg <= 9'b101110110;
      13'h106: filaimg <= 9'b101110110;
      13'h107: filaimg <= 9'b101110110;
      13'h108: filaimg <= 9'b101110110;
      13'h109: filaimg <= 9'b101110110;
      13'h10A: filaimg <= 9'b101110110;
      13'h10B: filaimg <= 9'b101110110;
      13'h10C: filaimg <= 9'b101110110;
      13'h10D: filaimg <= 9'b101110110;
      13'h10E: filaimg <= 9'b101110110;
      13'h10F: filaimg <= 9'b101110110;
      13'h110: filaimg <= 9'b101110110;
      13'h111: filaimg <= 9'b101110110;
      13'h112: filaimg <= 9'b101110110;
      13'h113: filaimg <= 9'b101110110;
      13'h114: filaimg <= 9'b101110110;
      13'h115: filaimg <= 9'b101110110;
      13'h116: filaimg <= 9'b101110110;
      13'h117: filaimg <= 9'b101110110;
      13'h118: filaimg <= 9'b101110110;
      13'h119: filaimg <= 9'b101110110;
      13'h11A: filaimg <= 9'b101110110;
      13'h11B: filaimg <= 9'b101110110;
      13'h11C: filaimg <= 9'b101110110;
      13'h11D: filaimg <= 9'b101110110;
      13'h11E: filaimg <= 9'b101110110;
      13'h11F: filaimg <= 9'b101110110;
      13'h120: filaimg <= 9'b101110110;
      13'h121: filaimg <= 9'b101110110;
      13'h122: filaimg <= 9'b101110110;
      13'h123: filaimg <= 9'b101110110;
      13'h124: filaimg <= 9'b101110110;
      13'h125: filaimg <= 9'b101110110;
      13'h126: filaimg <= 9'b101110110;
      13'h127: filaimg <= 9'b101110110;
      13'h128: filaimg <= 9'b101110110;
      13'h129: filaimg <= 9'b101110110;
      13'h12A: filaimg <= 9'b101110110;
      13'h12B: filaimg <= 9'b101110110;
      13'h12C: filaimg <= 9'b101110110;
      13'h12D: filaimg <= 9'b101110110;
      13'h12E: filaimg <= 9'b101110110;
      13'h12F: filaimg <= 9'b101110110;
      13'h130: filaimg <= 9'b101110110;
      13'h131: filaimg <= 9'b101110110;
      13'h132: filaimg <= 9'b101110110;
      13'h133: filaimg <= 9'b101110110;
      13'h134: filaimg <= 9'b101110110;
      13'h135: filaimg <= 9'b101110110;
      13'h136: filaimg <= 9'b101110110;
      13'h137: filaimg <= 9'b101110110;
      13'h138: filaimg <= 9'b101110110;
      13'h139: filaimg <= 9'b101110110;
      13'h13A: filaimg <= 9'b101110110;
      13'h13B: filaimg <= 9'b101110110;
      13'h13C: filaimg <= 9'b101110110;
      13'h13D: filaimg <= 9'b101110110;
      13'h13E: filaimg <= 9'b101110110;
      13'h13F: filaimg <= 9'b101110110;
      13'h140: filaimg <= 9'b101110110;
      13'h141: filaimg <= 9'b101110110;
      13'h142: filaimg <= 9'b101110110;
      13'h143: filaimg <= 9'b101110110;
      13'h144: filaimg <= 9'b101110110;
      13'h145: filaimg <= 9'b101110110;
      13'h146: filaimg <= 9'b101110110;
      13'h147: filaimg <= 9'b101110110;
      13'h148: filaimg <= 9'b101110110;
      13'h149: filaimg <= 9'b101110110;
      13'h14A: filaimg <= 9'b101110110;
      13'h14B: filaimg <= 9'b101110110;
      13'h14C: filaimg <= 9'b101110110;
      13'h14D: filaimg <= 9'b101110110;
      13'h14E: filaimg <= 9'b101110110;
      13'h14F: filaimg <= 9'b101110110;
      13'h150: filaimg <= 9'b101110110;
      13'h151: filaimg <= 9'b101110110;
      13'h152: filaimg <= 9'b101110110;
      13'h153: filaimg <= 9'b101110110;
      13'h154: filaimg <= 9'b101110110;
      13'h155: filaimg <= 9'b101110110;
      13'h156: filaimg <= 9'b101110110;
      13'h157: filaimg <= 9'b101110110;
      13'h158: filaimg <= 9'b101110110;
      13'h159: filaimg <= 9'b101110110;
      13'h15A: filaimg <= 9'b101110110;
      13'h15B: filaimg <= 9'b101110110;
      13'h15C: filaimg <= 9'b101110110;
      13'h15D: filaimg <= 9'b101110110;
      13'h15E: filaimg <= 9'b101110110;
      13'h15F: filaimg <= 9'b101110110;
      13'h160: filaimg <= 9'b101110110;
      13'h161: filaimg <= 9'b101110110;
      13'h162: filaimg <= 9'b101110110;
      13'h163: filaimg <= 9'b101110110;
      13'h164: filaimg <= 9'b101110110;
      13'h165: filaimg <= 9'b101110110;
      13'h166: filaimg <= 9'b101110110;
      13'h167: filaimg <= 9'b101110110;
      13'h168: filaimg <= 9'b101110110;
      13'h169: filaimg <= 9'b101110110;
      13'h16A: filaimg <= 9'b101110110;
      13'h16B: filaimg <= 9'b101110110;
      13'h16C: filaimg <= 9'b101110110;
      13'h16D: filaimg <= 9'b101110110;
      13'h16E: filaimg <= 9'b101110110;
      13'h16F: filaimg <= 9'b101110110;
      13'h170: filaimg <= 9'b101110110;
      13'h171: filaimg <= 9'b101110110;
      13'h172: filaimg <= 9'b101110110;
      13'h173: filaimg <= 9'b101110110;
      13'h174: filaimg <= 9'b101110110;
      13'h175: filaimg <= 9'b101110110;
      13'h176: filaimg <= 9'b101110110;
      13'h177: filaimg <= 9'b101110110;
      13'h178: filaimg <= 9'b101110110;
      13'h179: filaimg <= 9'b101110110;
      13'h17A: filaimg <= 9'b101110110;
      13'h17B: filaimg <= 9'b101110110;
      13'h17C: filaimg <= 9'b101110110;
      13'h17D: filaimg <= 9'b101110110;
      13'h17E: filaimg <= 9'b101110110;
      13'h17F: filaimg <= 9'b101110110;
      13'h180: filaimg <= 9'b101110110;
      13'h181: filaimg <= 9'b101110110;
      13'h182: filaimg <= 9'b101110110;
      13'h183: filaimg <= 9'b101110110;
      13'h184: filaimg <= 9'b101110110;
      13'h185: filaimg <= 9'b101110110;
      13'h186: filaimg <= 9'b101110110;
      13'h187: filaimg <= 9'b101110110;
      13'h188: filaimg <= 9'b101110110;
      13'h189: filaimg <= 9'b101110110;
      13'h18A: filaimg <= 9'b101110110;
      13'h18B: filaimg <= 9'b101110110;
      13'h18C: filaimg <= 9'b101110110;
      13'h18D: filaimg <= 9'b101110110;
      13'h18E: filaimg <= 9'b101110110;
      13'h18F: filaimg <= 9'b101110110;
      13'h190: filaimg <= 9'b101110110;
      13'h191: filaimg <= 9'b101110110;
      13'h192: filaimg <= 9'b101110110;
      13'h193: filaimg <= 9'b101110110;
      13'h194: filaimg <= 9'b101110110;
      13'h195: filaimg <= 9'b101110110;
      13'h196: filaimg <= 9'b101110110;
      13'h197: filaimg <= 9'b101110110;
      13'h198: filaimg <= 9'b101110110;
      13'h199: filaimg <= 9'b101110110;
      13'h19A: filaimg <= 9'b101110110;
      13'h19B: filaimg <= 9'b101110110;
      13'h19C: filaimg <= 9'b101110110;
      13'h19D: filaimg <= 9'b101110110;
      13'h19E: filaimg <= 9'b101110110;
      13'h19F: filaimg <= 9'b101110110;
      13'h1A0: filaimg <= 9'b101110110;
      13'h1A1: filaimg <= 9'b101110110;
      13'h1A2: filaimg <= 9'b101110110;
      13'h1A3: filaimg <= 9'b101110110;
      13'h1A4: filaimg <= 9'b101110110;
      13'h1A5: filaimg <= 9'b101110110;
      13'h1A6: filaimg <= 9'b101110110;
      13'h1A7: filaimg <= 9'b101110110;
      13'h1A8: filaimg <= 9'b101110110;
      13'h1A9: filaimg <= 9'b101110110;
      13'h1AA: filaimg <= 9'b101110110;
      13'h1AB: filaimg <= 9'b101110110;
      13'h1AC: filaimg <= 9'b101110110;
      13'h1AD: filaimg <= 9'b101110110;
      13'h1AE: filaimg <= 9'b101110110;
      13'h1AF: filaimg <= 9'b101110110;
      13'h1B0: filaimg <= 9'b101110110;
      13'h1B1: filaimg <= 9'b101110110;
      13'h1B2: filaimg <= 9'b101110110;
      13'h1B3: filaimg <= 9'b101110110;
      13'h1B4: filaimg <= 9'b101110110;
      13'h1B5: filaimg <= 9'b101110110;
      13'h1B6: filaimg <= 9'b101110110;
      13'h1B7: filaimg <= 9'b101110110;
      13'h1B8: filaimg <= 9'b101110110;
      13'h1B9: filaimg <= 9'b101110110;
      13'h1BA: filaimg <= 9'b101110110;
      13'h1BB: filaimg <= 9'b101110110;
      13'h1BC: filaimg <= 9'b101110110;
      13'h1BD: filaimg <= 9'b101110110;
      13'h1BE: filaimg <= 9'b101110110;
      13'h1BF: filaimg <= 9'b101110110;
      13'h1C0: filaimg <= 9'b101110110;
      13'h1C1: filaimg <= 9'b101110110;
      13'h1C2: filaimg <= 9'b101110110;
      13'h1C3: filaimg <= 9'b101110110;
      13'h1C4: filaimg <= 9'b101110110;
      13'h1C5: filaimg <= 9'b101110110;
      13'h1C6: filaimg <= 9'b101110110;
      13'h1C7: filaimg <= 9'b101110110;
      13'h1C8: filaimg <= 9'b101110110;
      13'h1C9: filaimg <= 9'b101110110;
      13'h1CA: filaimg <= 9'b101110110;
      13'h1CB: filaimg <= 9'b101110110;
      13'h1CC: filaimg <= 9'b101110110;
      13'h1CD: filaimg <= 9'b101110110;
      13'h1CE: filaimg <= 9'b101110110;
      13'h1CF: filaimg <= 9'b101110110;
      13'h1D0: filaimg <= 9'b101110110;
      13'h1D1: filaimg <= 9'b101110110;
      13'h1D2: filaimg <= 9'b101110110;
      13'h1D3: filaimg <= 9'b101110110;
      13'h1D4: filaimg <= 9'b101110110;
      13'h1D5: filaimg <= 9'b101110110;
      13'h1D6: filaimg <= 9'b101110110;
      13'h1D7: filaimg <= 9'b101110110;
      13'h1D8: filaimg <= 9'b101110110;
      13'h1D9: filaimg <= 9'b101110110;
      13'h1DA: filaimg <= 9'b101110110;
      13'h1DB: filaimg <= 9'b101110110;
      13'h1DC: filaimg <= 9'b101110110;
      13'h1DD: filaimg <= 9'b101110110;
      13'h1DE: filaimg <= 9'b101110110;
      13'h1DF: filaimg <= 9'b101110110;
      13'h1E0: filaimg <= 9'b101110110;
      13'h1E1: filaimg <= 9'b101110110;
      13'h1E2: filaimg <= 9'b101110110;
      13'h1E3: filaimg <= 9'b101110110;
      13'h1E4: filaimg <= 9'b101110110;
      13'h1E5: filaimg <= 9'b101110110;
      13'h1E6: filaimg <= 9'b101110110;
      13'h1E7: filaimg <= 9'b101110110;
      13'h1E8: filaimg <= 9'b101110110;
      13'h1E9: filaimg <= 9'b101110110;
      13'h1EA: filaimg <= 9'b101110110;
      13'h1EB: filaimg <= 9'b101110110;
      13'h1EC: filaimg <= 9'b101110110;
      13'h1ED: filaimg <= 9'b101110110;
      13'h1EE: filaimg <= 9'b101110110;
      13'h1EF: filaimg <= 9'b101110110;
      13'h1F0: filaimg <= 9'b101110110;
      13'h1F1: filaimg <= 9'b101110110;
      13'h1F2: filaimg <= 9'b101110110;
      13'h1F3: filaimg <= 9'b101110110;
      13'h1F4: filaimg <= 9'b101110110;
      13'h1F5: filaimg <= 9'b101110110;
      13'h1F6: filaimg <= 9'b101110110;
      13'h1F7: filaimg <= 9'b101110110;
      13'h1F8: filaimg <= 9'b101110110;
      13'h1F9: filaimg <= 9'b101110110;
      13'h1FA: filaimg <= 9'b101110110;
      13'h1FB: filaimg <= 9'b101110110;
      13'h1FC: filaimg <= 9'b101110110;
      13'h1FD: filaimg <= 9'b101110110;
      13'h1FE: filaimg <= 9'b101110110;
      13'h1FF: filaimg <= 9'b101110110;
      13'h200: filaimg <= 9'b101110110;
      13'h201: filaimg <= 9'b101110110;
      13'h202: filaimg <= 9'b101110110;
      13'h203: filaimg <= 9'b101110110;
      13'h204: filaimg <= 9'b101110110;
      13'h205: filaimg <= 9'b101110110;
      13'h206: filaimg <= 9'b101110110;
      13'h207: filaimg <= 9'b101110110;
      13'h208: filaimg <= 9'b101110110;
      13'h209: filaimg <= 9'b101110110;
      13'h20A: filaimg <= 9'b101110110;
      13'h20B: filaimg <= 9'b101110110;
      13'h20C: filaimg <= 9'b101110110;
      13'h20D: filaimg <= 9'b101110110;
      13'h20E: filaimg <= 9'b101110110;
      13'h20F: filaimg <= 9'b101110110;
      13'h210: filaimg <= 9'b101110110;
      13'h211: filaimg <= 9'b101110110;
      13'h212: filaimg <= 9'b101110110;
      13'h213: filaimg <= 9'b101110110;
      13'h214: filaimg <= 9'b101110110;
      13'h215: filaimg <= 9'b101110110;
      13'h216: filaimg <= 9'b101110110;
      13'h217: filaimg <= 9'b101110110;
      13'h218: filaimg <= 9'b101110110;
      13'h219: filaimg <= 9'b101110110;
      13'h21A: filaimg <= 9'b101110110;
      13'h21B: filaimg <= 9'b101110110;
      13'h21C: filaimg <= 9'b101110110;
      13'h21D: filaimg <= 9'b101110110;
      13'h21E: filaimg <= 9'b101110110;
      13'h21F: filaimg <= 9'b101110110;
      13'h220: filaimg <= 9'b101110110;
      13'h221: filaimg <= 9'b101110110;
      13'h222: filaimg <= 9'b101110110;
      13'h223: filaimg <= 9'b101110110;
      13'h224: filaimg <= 9'b101110110;
      13'h225: filaimg <= 9'b101110110;
      13'h226: filaimg <= 9'b101110110;
      13'h227: filaimg <= 9'b101110110;
      13'h228: filaimg <= 9'b101110110;
      13'h229: filaimg <= 9'b101110110;
      13'h22A: filaimg <= 9'b101110110;
      13'h22B: filaimg <= 9'b101110110;
      13'h22C: filaimg <= 9'b101110110;
      13'h22D: filaimg <= 9'b101110110;
      13'h22E: filaimg <= 9'b101110110;
      13'h22F: filaimg <= 9'b101110110;
      13'h230: filaimg <= 9'b101110110;
      13'h231: filaimg <= 9'b101110110;
      13'h232: filaimg <= 9'b101110110;
      13'h233: filaimg <= 9'b101110110;
      13'h234: filaimg <= 9'b101110110;
      13'h235: filaimg <= 9'b101110110;
      13'h236: filaimg <= 9'b101110110;
      13'h237: filaimg <= 9'b101110110;
      13'h238: filaimg <= 9'b101110110;
      13'h239: filaimg <= 9'b101110110;
      13'h23A: filaimg <= 9'b101110110;
      13'h23B: filaimg <= 9'b101110110;
      13'h23C: filaimg <= 9'b101110110;
      13'h23D: filaimg <= 9'b101110110;
      13'h23E: filaimg <= 9'b101110110;
      13'h23F: filaimg <= 9'b101110110;
      13'h240: filaimg <= 9'b101110110;
      13'h241: filaimg <= 9'b101110110;
      13'h242: filaimg <= 9'b101110110;
      13'h243: filaimg <= 9'b101110110;
      13'h244: filaimg <= 9'b101110110;
      13'h245: filaimg <= 9'b101110110;
      13'h246: filaimg <= 9'b101110110;
      13'h247: filaimg <= 9'b101110110;
      13'h248: filaimg <= 9'b101110110;
      13'h249: filaimg <= 9'b101110110;
      13'h24A: filaimg <= 9'b101110110;
      13'h24B: filaimg <= 9'b101110110;
      13'h24C: filaimg <= 9'b101110110;
      13'h24D: filaimg <= 9'b101110110;
      13'h24E: filaimg <= 9'b101110110;
      13'h24F: filaimg <= 9'b101110110;
      13'h250: filaimg <= 9'b101110110;
      13'h251: filaimg <= 9'b101110110;
      13'h252: filaimg <= 9'b101110110;
      13'h253: filaimg <= 9'b101110110;
      13'h254: filaimg <= 9'b101110110;
      13'h255: filaimg <= 9'b101110110;
      13'h256: filaimg <= 9'b101110110;
      13'h257: filaimg <= 9'b101110110;
      13'h258: filaimg <= 9'b101110110;
      13'h259: filaimg <= 9'b101110110;
      13'h25A: filaimg <= 9'b101110110;
      13'h25B: filaimg <= 9'b101110110;
      13'h25C: filaimg <= 9'b101110110;
      13'h25D: filaimg <= 9'b101110110;
      13'h25E: filaimg <= 9'b101110110;
      13'h25F: filaimg <= 9'b101110110;
      13'h260: filaimg <= 9'b101110110;
      13'h261: filaimg <= 9'b101110110;
      13'h262: filaimg <= 9'b101110110;
      13'h263: filaimg <= 9'b101110110;
      13'h264: filaimg <= 9'b101110110;
      13'h265: filaimg <= 9'b101110110;
      13'h266: filaimg <= 9'b101110110;
      13'h267: filaimg <= 9'b101110110;
      13'h268: filaimg <= 9'b101110110;
      13'h269: filaimg <= 9'b101110110;
      13'h26A: filaimg <= 9'b101110110;
      13'h26B: filaimg <= 9'b101110110;
      13'h26C: filaimg <= 9'b101110110;
      13'h26D: filaimg <= 9'b101110110;
      13'h26E: filaimg <= 9'b101110110;
      13'h26F: filaimg <= 9'b101110110;
      13'h270: filaimg <= 9'b101110110;
      13'h271: filaimg <= 9'b101110110;
      13'h272: filaimg <= 9'b101110110;
      13'h273: filaimg <= 9'b101110110;
      13'h274: filaimg <= 9'b101110110;
      13'h275: filaimg <= 9'b101110110;
      13'h276: filaimg <= 9'b101110110;
      13'h277: filaimg <= 9'b101110110;
      13'h278: filaimg <= 9'b101110110;
      13'h279: filaimg <= 9'b101110110;
      13'h27A: filaimg <= 9'b101110110;
      13'h27B: filaimg <= 9'b101110110;
      13'h27C: filaimg <= 9'b101110110;
      13'h27D: filaimg <= 9'b101110110;
      13'h27E: filaimg <= 9'b101110110;
      13'h27F: filaimg <= 9'b101110110;
      13'h280: filaimg <= 9'b101110110;
      13'h281: filaimg <= 9'b101110110;
      13'h282: filaimg <= 9'b101110110;
      13'h283: filaimg <= 9'b101110110;
      13'h284: filaimg <= 9'b101110110;
      13'h285: filaimg <= 9'b101110110;
      13'h286: filaimg <= 9'b101110110;
      13'h287: filaimg <= 9'b101110110;
      13'h288: filaimg <= 9'b101110110;
      13'h289: filaimg <= 9'b101110110;
      13'h28A: filaimg <= 9'b101110110;
      13'h28B: filaimg <= 9'b101110110;
      13'h28C: filaimg <= 9'b101110110;
      13'h28D: filaimg <= 9'b101110110;
      13'h28E: filaimg <= 9'b101110110;
      13'h28F: filaimg <= 9'b101110110;
      13'h290: filaimg <= 9'b101110110;
      13'h291: filaimg <= 9'b101110110;
      13'h292: filaimg <= 9'b101110110;
      13'h293: filaimg <= 9'b101110110;
      13'h294: filaimg <= 9'b101110110;
      13'h295: filaimg <= 9'b101110110;
      13'h296: filaimg <= 9'b101110110;
      13'h297: filaimg <= 9'b101110110;
      13'h298: filaimg <= 9'b101110110;
      13'h299: filaimg <= 9'b101110110;
      13'h29A: filaimg <= 9'b101110110;
      13'h29B: filaimg <= 9'b101110110;
      13'h29C: filaimg <= 9'b101110110;
      13'h29D: filaimg <= 9'b101110110;
      13'h29E: filaimg <= 9'b101110110;
      13'h29F: filaimg <= 9'b101110110;
      13'h2A0: filaimg <= 9'b101110110;
      13'h2A1: filaimg <= 9'b101110110;
      13'h2A2: filaimg <= 9'b101110110;
      13'h2A3: filaimg <= 9'b101110110;
      13'h2A4: filaimg <= 9'b101110110;
      13'h2A5: filaimg <= 9'b101110110;
      13'h2A6: filaimg <= 9'b101110110;
      13'h2A7: filaimg <= 9'b101110110;
      13'h2A8: filaimg <= 9'b101110110;
      13'h2A9: filaimg <= 9'b101110110;
      13'h2AA: filaimg <= 9'b101110110;
      13'h2AB: filaimg <= 9'b101110110;
      13'h2AC: filaimg <= 9'b101110110;
      13'h2AD: filaimg <= 9'b101110110;
      13'h2AE: filaimg <= 9'b101110110;
      13'h2AF: filaimg <= 9'b101110110;
      13'h2B0: filaimg <= 9'b101110110;
      13'h2B1: filaimg <= 9'b101110110;
      13'h2B2: filaimg <= 9'b101110110;
      13'h2B3: filaimg <= 9'b101110110;
      13'h2B4: filaimg <= 9'b101110110;
      13'h2B5: filaimg <= 9'b101110110;
      13'h2B6: filaimg <= 9'b101110110;
      13'h2B7: filaimg <= 9'b101110110;
      13'h2B8: filaimg <= 9'b101110110;
      13'h2B9: filaimg <= 9'b101110110;
      13'h2BA: filaimg <= 9'b101110110;
      13'h2BB: filaimg <= 9'b101110110;
      13'h2BC: filaimg <= 9'b101110110;
      13'h2BD: filaimg <= 9'b101110110;
      13'h2BE: filaimg <= 9'b101110110;
      13'h2BF: filaimg <= 9'b101110110;
      13'h2C0: filaimg <= 9'b101110110;
      13'h2C1: filaimg <= 9'b101110110;
      13'h2C2: filaimg <= 9'b101110110;
      13'h2C3: filaimg <= 9'b101110110;
      13'h2C4: filaimg <= 9'b101110110;
      13'h2C5: filaimg <= 9'b101110110;
      13'h2C6: filaimg <= 9'b101110110;
      13'h2C7: filaimg <= 9'b101110110;
      13'h2C8: filaimg <= 9'b101110110;
      13'h2C9: filaimg <= 9'b101110110;
      13'h2CA: filaimg <= 9'b101110110;
      13'h2CB: filaimg <= 9'b101110110;
      13'h2CC: filaimg <= 9'b101110110;
      13'h2CD: filaimg <= 9'b101110110;
      13'h2CE: filaimg <= 9'b101110110;
      13'h2CF: filaimg <= 9'b101110110;
      13'h2D0: filaimg <= 9'b101110110;
      13'h2D1: filaimg <= 9'b101110110;
      13'h2D2: filaimg <= 9'b101110110;
      13'h2D3: filaimg <= 9'b101110110;
      13'h2D4: filaimg <= 9'b101110110;
      13'h2D5: filaimg <= 9'b101110110;
      13'h2D6: filaimg <= 9'b101110110;
      13'h2D7: filaimg <= 9'b101110110;
      13'h2D8: filaimg <= 9'b101110110;
      13'h2D9: filaimg <= 9'b101110110;
      13'h2DA: filaimg <= 9'b101110110;
      13'h2DB: filaimg <= 9'b101110110;
      13'h2DC: filaimg <= 9'b101110110;
      13'h2DD: filaimg <= 9'b101110110;
      13'h2DE: filaimg <= 9'b101110110;
      13'h2DF: filaimg <= 9'b101110110;
      13'h2E0: filaimg <= 9'b101110110;
      13'h2E1: filaimg <= 9'b101110110;
      13'h2E2: filaimg <= 9'b101110110;
      13'h2E3: filaimg <= 9'b101110110;
      13'h2E4: filaimg <= 9'b101110110;
      13'h2E5: filaimg <= 9'b101110110;
      13'h2E6: filaimg <= 9'b101110110;
      13'h2E7: filaimg <= 9'b101110110;
      13'h2E8: filaimg <= 9'b101110110;
      13'h2E9: filaimg <= 9'b101110110;
      13'h2EA: filaimg <= 9'b101110110;
      13'h2EB: filaimg <= 9'b101110110;
      13'h2EC: filaimg <= 9'b101110110;
      13'h2ED: filaimg <= 9'b101110110;
      13'h2EE: filaimg <= 9'b101110110;
      13'h2EF: filaimg <= 9'b101110110;
      13'h2F0: filaimg <= 9'b101110110;
      13'h2F1: filaimg <= 9'b101110110;
      13'h2F2: filaimg <= 9'b101110110;
      13'h2F3: filaimg <= 9'b101110110;
      13'h2F4: filaimg <= 9'b101110110;
      13'h2F5: filaimg <= 9'b101110110;
      13'h2F6: filaimg <= 9'b101110110;
      13'h2F7: filaimg <= 9'b101110110;
      13'h2F8: filaimg <= 9'b101110110;
      13'h2F9: filaimg <= 9'b101110110;
      13'h2FA: filaimg <= 9'b101110110;
      13'h2FB: filaimg <= 9'b101110110;
      13'h2FC: filaimg <= 9'b101110110;
      13'h2FD: filaimg <= 9'b101110110;
      13'h2FE: filaimg <= 9'b101110110;
      13'h2FF: filaimg <= 9'b101110110;
      13'h300: filaimg <= 9'b101110110;
      13'h301: filaimg <= 9'b101110110;
      13'h302: filaimg <= 9'b101110110;
      13'h303: filaimg <= 9'b101110110;
      13'h304: filaimg <= 9'b101110110;
      13'h305: filaimg <= 9'b101110110;
      13'h306: filaimg <= 9'b101110110;
      13'h307: filaimg <= 9'b101110110;
      13'h308: filaimg <= 9'b101110110;
      13'h309: filaimg <= 9'b101110110;
      13'h30A: filaimg <= 9'b101110110;
      13'h30B: filaimg <= 9'b101110110;
      13'h30C: filaimg <= 9'b101110110;
      13'h30D: filaimg <= 9'b101110110;
      13'h30E: filaimg <= 9'b101110110;
      13'h30F: filaimg <= 9'b101110110;
      13'h310: filaimg <= 9'b101110110;
      13'h311: filaimg <= 9'b101110110;
      13'h312: filaimg <= 9'b101110110;
      13'h313: filaimg <= 9'b101110110;
      13'h314: filaimg <= 9'b101110110;
      13'h315: filaimg <= 9'b101110110;
      13'h316: filaimg <= 9'b101110110;
      13'h317: filaimg <= 9'b101110110;
      13'h318: filaimg <= 9'b101110110;
      13'h319: filaimg <= 9'b101110110;
      13'h31A: filaimg <= 9'b101110110;
      13'h31B: filaimg <= 9'b101110110;
      13'h31C: filaimg <= 9'b101110110;
      13'h31D: filaimg <= 9'b101110110;
      13'h31E: filaimg <= 9'b101110110;
      13'h31F: filaimg <= 9'b101110110;
      13'h320: filaimg <= 9'b101110110;
      13'h321: filaimg <= 9'b101110110;
      13'h322: filaimg <= 9'b101110110;
      13'h323: filaimg <= 9'b101110110;
      13'h324: filaimg <= 9'b101110110;
      13'h325: filaimg <= 9'b101110110;
      13'h326: filaimg <= 9'b101110110;
      13'h327: filaimg <= 9'b101110110;
      13'h328: filaimg <= 9'b101110110;
      13'h329: filaimg <= 9'b101110110;
      13'h32A: filaimg <= 9'b101110110;
      13'h32B: filaimg <= 9'b101110110;
      13'h32C: filaimg <= 9'b101110110;
      13'h32D: filaimg <= 9'b101110110;
      13'h32E: filaimg <= 9'b101110110;
      13'h32F: filaimg <= 9'b101110110;
      13'h330: filaimg <= 9'b101110110;
      13'h331: filaimg <= 9'b101110110;
      13'h332: filaimg <= 9'b101110110;
      13'h333: filaimg <= 9'b101110110;
      13'h334: filaimg <= 9'b101110110;
      13'h335: filaimg <= 9'b101110110;
      13'h336: filaimg <= 9'b101110110;
      13'h337: filaimg <= 9'b101110110;
      13'h338: filaimg <= 9'b101110110;
      13'h339: filaimg <= 9'b101110110;
      13'h33A: filaimg <= 9'b101110110;
      13'h33B: filaimg <= 9'b101110110;
      13'h33C: filaimg <= 9'b101110110;
      13'h33D: filaimg <= 9'b101110110;
      13'h33E: filaimg <= 9'b101110110;
      13'h33F: filaimg <= 9'b101110110;
      13'h340: filaimg <= 9'b101110110;
      13'h341: filaimg <= 9'b101110110;
      13'h342: filaimg <= 9'b101110110;
      13'h343: filaimg <= 9'b101110110;
      13'h344: filaimg <= 9'b101110110;
      13'h345: filaimg <= 9'b101110110;
      13'h346: filaimg <= 9'b101110110;
      13'h347: filaimg <= 9'b101110110;
      13'h348: filaimg <= 9'b101110110;
      13'h349: filaimg <= 9'b101110110;
      13'h34A: filaimg <= 9'b101110110;
      13'h34B: filaimg <= 9'b101110110;
      13'h34C: filaimg <= 9'b101110110;
      13'h34D: filaimg <= 9'b101110110;
      13'h34E: filaimg <= 9'b101110110;
      13'h34F: filaimg <= 9'b101110110;
      13'h350: filaimg <= 9'b101110110;
      13'h351: filaimg <= 9'b101110110;
      13'h352: filaimg <= 9'b101110110;
      13'h353: filaimg <= 9'b101110110;
      13'h354: filaimg <= 9'b101110110;
      13'h355: filaimg <= 9'b101110110;
      13'h356: filaimg <= 9'b101110110;
      13'h357: filaimg <= 9'b101110110;
      13'h358: filaimg <= 9'b101110110;
      13'h359: filaimg <= 9'b101110110;
      13'h35A: filaimg <= 9'b101110110;
      13'h35B: filaimg <= 9'b101110110;
      13'h35C: filaimg <= 9'b101110110;
      13'h35D: filaimg <= 9'b101110110;
      13'h35E: filaimg <= 9'b101110110;
      13'h35F: filaimg <= 9'b101110110;
      13'h360: filaimg <= 9'b101110110;
      13'h361: filaimg <= 9'b101110110;
      13'h362: filaimg <= 9'b101110110;
      13'h363: filaimg <= 9'b101110110;
      13'h364: filaimg <= 9'b101110110;
      13'h365: filaimg <= 9'b101110110;
      13'h366: filaimg <= 9'b101110110;
      13'h367: filaimg <= 9'b101110110;
      13'h368: filaimg <= 9'b101110110;
      13'h369: filaimg <= 9'b101110110;
      13'h36A: filaimg <= 9'b101110110;
      13'h36B: filaimg <= 9'b101110110;
      13'h36C: filaimg <= 9'b101110110;
      13'h36D: filaimg <= 9'b101110110;
      13'h36E: filaimg <= 9'b101110110;
      13'h36F: filaimg <= 9'b101110110;
      13'h370: filaimg <= 9'b101110110;
      13'h371: filaimg <= 9'b101110110;
      13'h372: filaimg <= 9'b101110110;
      13'h373: filaimg <= 9'b101110110;
      13'h374: filaimg <= 9'b101110110;
      13'h375: filaimg <= 9'b101110110;
      13'h376: filaimg <= 9'b101110110;
      13'h377: filaimg <= 9'b101110110;
      13'h378: filaimg <= 9'b101110110;
      13'h379: filaimg <= 9'b101110110;
      13'h37A: filaimg <= 9'b101110110;
      13'h37B: filaimg <= 9'b101110110;
      13'h37C: filaimg <= 9'b101110110;
      13'h37D: filaimg <= 9'b101110110;
      13'h37E: filaimg <= 9'b101110110;
      13'h37F: filaimg <= 9'b101110110;
      13'h380: filaimg <= 9'b101110110;
      13'h381: filaimg <= 9'b101110110;
      13'h382: filaimg <= 9'b101110110;
      13'h383: filaimg <= 9'b101110110;
      13'h384: filaimg <= 9'b101110110;
      13'h385: filaimg <= 9'b101110110;
      13'h386: filaimg <= 9'b101110110;
      13'h387: filaimg <= 9'b101110110;
      13'h388: filaimg <= 9'b101110110;
      13'h389: filaimg <= 9'b101110110;
      13'h38A: filaimg <= 9'b101110110;
      13'h38B: filaimg <= 9'b101110110;
      13'h38C: filaimg <= 9'b101110110;
      13'h38D: filaimg <= 9'b101110110;
      13'h38E: filaimg <= 9'b101110110;
      13'h38F: filaimg <= 9'b101110110;
      13'h390: filaimg <= 9'b101110110;
      13'h391: filaimg <= 9'b101110110;
      13'h392: filaimg <= 9'b101110110;
      13'h393: filaimg <= 9'b101110110;
      13'h394: filaimg <= 9'b101110110;
      13'h395: filaimg <= 9'b101110110;
      13'h396: filaimg <= 9'b101110110;
      13'h397: filaimg <= 9'b101110110;
      13'h398: filaimg <= 9'b101110110;
      13'h399: filaimg <= 9'b101110110;
      13'h39A: filaimg <= 9'b101110110;
      13'h39B: filaimg <= 9'b101110110;
      13'h39C: filaimg <= 9'b101110110;
      13'h39D: filaimg <= 9'b101110110;
      13'h39E: filaimg <= 9'b101110110;
      13'h39F: filaimg <= 9'b101110110;
      13'h3A0: filaimg <= 9'b101110110;
      13'h3A1: filaimg <= 9'b101110110;
      13'h3A2: filaimg <= 9'b101110110;
      13'h3A3: filaimg <= 9'b101110110;
      13'h3A4: filaimg <= 9'b101110110;
      13'h3A5: filaimg <= 9'b101110110;
      13'h3A6: filaimg <= 9'b101110110;
      13'h3A7: filaimg <= 9'b101110110;
      13'h3A8: filaimg <= 9'b101110110;
      13'h3A9: filaimg <= 9'b101110110;
      13'h3AA: filaimg <= 9'b101110110;
      13'h3AB: filaimg <= 9'b101110110;
      13'h3AC: filaimg <= 9'b101110110;
      13'h3AD: filaimg <= 9'b101110110;
      13'h3AE: filaimg <= 9'b101110110;
      13'h3AF: filaimg <= 9'b101110110;
      13'h3B0: filaimg <= 9'b101110110;
      13'h3B1: filaimg <= 9'b101110110;
      13'h3B2: filaimg <= 9'b101110110;
      13'h3B3: filaimg <= 9'b101110110;
      13'h3B4: filaimg <= 9'b101110110;
      13'h3B5: filaimg <= 9'b101110110;
      13'h3B6: filaimg <= 9'b101110110;
      13'h3B7: filaimg <= 9'b101110110;
      13'h3B8: filaimg <= 9'b101110110;
      13'h3B9: filaimg <= 9'b101110110;
      13'h3BA: filaimg <= 9'b101110110;
      13'h3BB: filaimg <= 9'b101110110;
      13'h3BC: filaimg <= 9'b101110110;
      13'h3BD: filaimg <= 9'b101110110;
      13'h3BE: filaimg <= 9'b101110110;
      13'h3BF: filaimg <= 9'b101110110;
      13'h3C0: filaimg <= 9'b101110110;
      13'h3C1: filaimg <= 9'b101110110;
      13'h3C2: filaimg <= 9'b101110110;
      13'h3C3: filaimg <= 9'b101110110;
      13'h3C4: filaimg <= 9'b101110110;
      13'h3C5: filaimg <= 9'b101110110;
      13'h3C6: filaimg <= 9'b101110110;
      13'h3C7: filaimg <= 9'b101110110;
      13'h3C8: filaimg <= 9'b101110110;
      13'h3C9: filaimg <= 9'b101110110;
      13'h3CA: filaimg <= 9'b101110110;
      13'h3CB: filaimg <= 9'b101110110;
      13'h3CC: filaimg <= 9'b101110110;
      13'h3CD: filaimg <= 9'b101110110;
      13'h3CE: filaimg <= 9'b101110110;
      13'h3CF: filaimg <= 9'b101110110;
      13'h3D0: filaimg <= 9'b101110110;
      13'h3D1: filaimg <= 9'b101110110;
      13'h3D2: filaimg <= 9'b101110110;
      13'h3D3: filaimg <= 9'b101110110;
      13'h3D4: filaimg <= 9'b101110110;
      13'h3D5: filaimg <= 9'b101110110;
      13'h3D6: filaimg <= 9'b101110110;
      13'h3D7: filaimg <= 9'b101110110;
      13'h3D8: filaimg <= 9'b101110110;
      13'h3D9: filaimg <= 9'b101110110;
      13'h3DA: filaimg <= 9'b101110110;
      13'h3DB: filaimg <= 9'b101110110;
      13'h3DC: filaimg <= 9'b101110110;
      13'h3DD: filaimg <= 9'b101110110;
      13'h3DE: filaimg <= 9'b101110110;
      13'h3DF: filaimg <= 9'b101110110;
      13'h3E0: filaimg <= 9'b101110110;
      13'h3E1: filaimg <= 9'b101110110;
      13'h3E2: filaimg <= 9'b101110110;
      13'h3E3: filaimg <= 9'b101110110;
      13'h3E4: filaimg <= 9'b101110110;
      13'h3E5: filaimg <= 9'b101110110;
      13'h3E6: filaimg <= 9'b101110110;
      13'h3E7: filaimg <= 9'b101110110;
      13'h3E8: filaimg <= 9'b101110110;
      13'h3E9: filaimg <= 9'b101110110;
      13'h3EA: filaimg <= 9'b101110110;
      13'h3EB: filaimg <= 9'b101110110;
      13'h3EC: filaimg <= 9'b101110110;
      13'h3ED: filaimg <= 9'b101110110;
      13'h3EE: filaimg <= 9'b101110110;
      13'h3EF: filaimg <= 9'b101110110;
      13'h3F0: filaimg <= 9'b101110110;
      13'h3F1: filaimg <= 9'b101110110;
      13'h3F2: filaimg <= 9'b101110110;
      13'h3F3: filaimg <= 9'b101110110;
      13'h3F4: filaimg <= 9'b101110110;
      13'h3F5: filaimg <= 9'b101110110;
      13'h3F6: filaimg <= 9'b101110110;
      13'h3F7: filaimg <= 9'b101110110;
      13'h3F8: filaimg <= 9'b101110110;
      13'h3F9: filaimg <= 9'b101110110;
      13'h3FA: filaimg <= 9'b101110110;
      13'h3FB: filaimg <= 9'b101110110;
      13'h3FC: filaimg <= 9'b101110110;
      13'h3FD: filaimg <= 9'b101110110;
      13'h3FE: filaimg <= 9'b101110110;
      13'h3FF: filaimg <= 9'b101110110;
      13'h400: filaimg <= 9'b101110110;
      13'h401: filaimg <= 9'b101110110;
      13'h402: filaimg <= 9'b101110110;
      13'h403: filaimg <= 9'b101110110;
      13'h404: filaimg <= 9'b101110110;
      13'h405: filaimg <= 9'b101110110;
      13'h406: filaimg <= 9'b101110110;
      13'h407: filaimg <= 9'b101110110;
      13'h408: filaimg <= 9'b101110110;
      13'h409: filaimg <= 9'b101110110;
      13'h40A: filaimg <= 9'b101110110;
      13'h40B: filaimg <= 9'b101110110;
      13'h40C: filaimg <= 9'b101110110;
      13'h40D: filaimg <= 9'b101110110;
      13'h40E: filaimg <= 9'b101110110;
      13'h40F: filaimg <= 9'b101110110;
      13'h410: filaimg <= 9'b101110110;
      13'h411: filaimg <= 9'b101110110;
      13'h412: filaimg <= 9'b101110110;
      13'h413: filaimg <= 9'b101110110;
      13'h414: filaimg <= 9'b101110110;
      13'h415: filaimg <= 9'b101110110;
      13'h416: filaimg <= 9'b101110110;
      13'h417: filaimg <= 9'b101110110;
      13'h418: filaimg <= 9'b101110110;
      13'h419: filaimg <= 9'b101110110;
      13'h41A: filaimg <= 9'b101110110;
      13'h41B: filaimg <= 9'b101110110;
      13'h41C: filaimg <= 9'b101110110;
      13'h41D: filaimg <= 9'b101110110;
      13'h41E: filaimg <= 9'b101110110;
      13'h41F: filaimg <= 9'b101110110;
      13'h420: filaimg <= 9'b101110110;
      13'h421: filaimg <= 9'b101110110;
      13'h422: filaimg <= 9'b101110110;
      13'h423: filaimg <= 9'b101110110;
      13'h424: filaimg <= 9'b101110110;
      13'h425: filaimg <= 9'b101110110;
      13'h426: filaimg <= 9'b101110110;
      13'h427: filaimg <= 9'b101110110;
      13'h428: filaimg <= 9'b101110110;
      13'h429: filaimg <= 9'b101110110;
      13'h42A: filaimg <= 9'b101110110;
      13'h42B: filaimg <= 9'b101110110;
      13'h42C: filaimg <= 9'b101110110;
      13'h42D: filaimg <= 9'b101110110;
      13'h42E: filaimg <= 9'b101110110;
      13'h42F: filaimg <= 9'b101110110;
      13'h430: filaimg <= 9'b101110110;
      13'h431: filaimg <= 9'b101110110;
      13'h432: filaimg <= 9'b101110110;
      13'h433: filaimg <= 9'b101110110;
      13'h434: filaimg <= 9'b101110110;
      13'h435: filaimg <= 9'b101110110;
      13'h436: filaimg <= 9'b101110110;
      13'h437: filaimg <= 9'b101110110;
      13'h438: filaimg <= 9'b101110110;
      13'h439: filaimg <= 9'b101110110;
      13'h43A: filaimg <= 9'b101110110;
      13'h43B: filaimg <= 9'b101110110;
      13'h43C: filaimg <= 9'b101110110;
      13'h43D: filaimg <= 9'b101110110;
      13'h43E: filaimg <= 9'b101110110;
      13'h43F: filaimg <= 9'b101110110;
      13'h440: filaimg <= 9'b101110110;
      13'h441: filaimg <= 9'b101110110;
      13'h442: filaimg <= 9'b101110110;
      13'h443: filaimg <= 9'b101110110;
      13'h444: filaimg <= 9'b101110110;
      13'h445: filaimg <= 9'b101110110;
      13'h446: filaimg <= 9'b101110110;
      13'h447: filaimg <= 9'b101110110;
      13'h448: filaimg <= 9'b101110110;
      13'h449: filaimg <= 9'b101110110;
      13'h44A: filaimg <= 9'b101110110;
      13'h44B: filaimg <= 9'b101110110;
      13'h44C: filaimg <= 9'b101110110;
      13'h44D: filaimg <= 9'b101110110;
      13'h44E: filaimg <= 9'b101110110;
      13'h44F: filaimg <= 9'b101110110;
      13'h450: filaimg <= 9'b101110110;
      13'h451: filaimg <= 9'b101110110;
      13'h452: filaimg <= 9'b101110110;
      13'h453: filaimg <= 9'b101110110;
      13'h454: filaimg <= 9'b101110110;
      13'h455: filaimg <= 9'b101110110;
      13'h456: filaimg <= 9'b101110110;
      13'h457: filaimg <= 9'b101110110;
      13'h458: filaimg <= 9'b101110110;
      13'h459: filaimg <= 9'b101110110;
      13'h45A: filaimg <= 9'b101110110;
      13'h45B: filaimg <= 9'b101110110;
      13'h45C: filaimg <= 9'b101110110;
      13'h45D: filaimg <= 9'b101110110;
      13'h45E: filaimg <= 9'b101110110;
      13'h45F: filaimg <= 9'b101110110;
      13'h460: filaimg <= 9'b101110110;
      13'h461: filaimg <= 9'b101110110;
      13'h462: filaimg <= 9'b101110110;
      13'h463: filaimg <= 9'b101110110;
      13'h464: filaimg <= 9'b101110110;
      13'h465: filaimg <= 9'b101110110;
      13'h466: filaimg <= 9'b101110110;
      13'h467: filaimg <= 9'b101110110;
      13'h468: filaimg <= 9'b101110110;
      13'h469: filaimg <= 9'b101110110;
      13'h46A: filaimg <= 9'b101110110;
      13'h46B: filaimg <= 9'b101110110;
      13'h46C: filaimg <= 9'b101110110;
      13'h46D: filaimg <= 9'b101110110;
      13'h46E: filaimg <= 9'b101110110;
      13'h46F: filaimg <= 9'b101110110;
      13'h470: filaimg <= 9'b101110110;
      13'h471: filaimg <= 9'b101110110;
      13'h472: filaimg <= 9'b101110110;
      13'h473: filaimg <= 9'b101110110;
      13'h474: filaimg <= 9'b101110110;
      13'h475: filaimg <= 9'b101110110;
      13'h476: filaimg <= 9'b101110110;
      13'h477: filaimg <= 9'b101110110;
      13'h478: filaimg <= 9'b101110110;
      13'h479: filaimg <= 9'b101110110;
      13'h47A: filaimg <= 9'b101110110;
      13'h47B: filaimg <= 9'b101110110;
      13'h47C: filaimg <= 9'b101110110;
      13'h47D: filaimg <= 9'b101110110;
      13'h47E: filaimg <= 9'b101110110;
      13'h47F: filaimg <= 9'b101110110;
      13'h480: filaimg <= 9'b101110110;
      13'h481: filaimg <= 9'b101110110;
      13'h482: filaimg <= 9'b101110110;
      13'h483: filaimg <= 9'b101110110;
      13'h484: filaimg <= 9'b101110110;
      13'h485: filaimg <= 9'b101110110;
      13'h486: filaimg <= 9'b101110110;
      13'h487: filaimg <= 9'b101110110;
      13'h488: filaimg <= 9'b101110110;
      13'h489: filaimg <= 9'b101110110;
      13'h48A: filaimg <= 9'b101110110;
      13'h48B: filaimg <= 9'b101110110;
      13'h48C: filaimg <= 9'b101110110;
      13'h48D: filaimg <= 9'b101110110;
      13'h48E: filaimg <= 9'b101110110;
      13'h48F: filaimg <= 9'b101110110;
      13'h490: filaimg <= 9'b101110110;
      13'h491: filaimg <= 9'b101110110;
      13'h492: filaimg <= 9'b101110110;
      13'h493: filaimg <= 9'b101110110;
      13'h494: filaimg <= 9'b101110110;
      13'h495: filaimg <= 9'b101110110;
      13'h496: filaimg <= 9'b101110110;
      13'h497: filaimg <= 9'b101110110;
      13'h498: filaimg <= 9'b101110110;
      13'h499: filaimg <= 9'b101110110;
      13'h49A: filaimg <= 9'b101110110;
      13'h49B: filaimg <= 9'b101110110;
      13'h49C: filaimg <= 9'b101110110;
      13'h49D: filaimg <= 9'b101110110;
      13'h49E: filaimg <= 9'b101110110;
      13'h49F: filaimg <= 9'b101110110;
      13'h4A0: filaimg <= 9'b101110110;
      13'h4A1: filaimg <= 9'b101110110;
      13'h4A2: filaimg <= 9'b101110110;
      13'h4A3: filaimg <= 9'b101110110;
      13'h4A4: filaimg <= 9'b101110110;
      13'h4A5: filaimg <= 9'b101110110;
      13'h4A6: filaimg <= 9'b101110110;
      13'h4A7: filaimg <= 9'b101110110;
      13'h4A8: filaimg <= 9'b101110110;
      13'h4A9: filaimg <= 9'b101110110;
      13'h4AA: filaimg <= 9'b101110110;
      13'h4AB: filaimg <= 9'b101110110;
      13'h4AC: filaimg <= 9'b101110110;
      13'h4AD: filaimg <= 9'b101110110;
      13'h4AE: filaimg <= 9'b101110110;
      13'h4AF: filaimg <= 9'b101110110;
      13'h4B0: filaimg <= 9'b101110110;
      13'h4B1: filaimg <= 9'b101110110;
      13'h4B2: filaimg <= 9'b101110110;
      13'h4B3: filaimg <= 9'b101110110;
      13'h4B4: filaimg <= 9'b101110110;
      13'h4B5: filaimg <= 9'b101110110;
      13'h4B6: filaimg <= 9'b101110110;
      13'h4B7: filaimg <= 9'b101110110;
      13'h4B8: filaimg <= 9'b101110110;
      13'h4B9: filaimg <= 9'b101110110;
      13'h4BA: filaimg <= 9'b101110110;
      13'h4BB: filaimg <= 9'b101110110;
      13'h4BC: filaimg <= 9'b101110110;
      13'h4BD: filaimg <= 9'b101110110;
      13'h4BE: filaimg <= 9'b101110110;
      13'h4BF: filaimg <= 9'b101110110;
      13'h4C0: filaimg <= 9'b101110110;
      13'h4C1: filaimg <= 9'b101110110;
      13'h4C2: filaimg <= 9'b101110110;
      13'h4C3: filaimg <= 9'b101110110;
      13'h4C4: filaimg <= 9'b101110110;
      13'h4C5: filaimg <= 9'b101110110;
      13'h4C6: filaimg <= 9'b101110110;
      13'h4C7: filaimg <= 9'b101110110;
      13'h4C8: filaimg <= 9'b101110110;
      13'h4C9: filaimg <= 9'b101110110;
      13'h4CA: filaimg <= 9'b101110110;
      13'h4CB: filaimg <= 9'b101110110;
      13'h4CC: filaimg <= 9'b101110110;
      13'h4CD: filaimg <= 9'b101110110;
      13'h4CE: filaimg <= 9'b101110110;
      13'h4CF: filaimg <= 9'b101110110;
      13'h4D0: filaimg <= 9'b101110110;
      13'h4D1: filaimg <= 9'b101110110;
      13'h4D2: filaimg <= 9'b101110110;
      13'h4D3: filaimg <= 9'b101110110;
      13'h4D4: filaimg <= 9'b101110110;
      13'h4D5: filaimg <= 9'b101110110;
      13'h4D6: filaimg <= 9'b101110110;
      13'h4D7: filaimg <= 9'b101110110;
      13'h4D8: filaimg <= 9'b101110110;
      13'h4D9: filaimg <= 9'b101110110;
      13'h4DA: filaimg <= 9'b101110110;
      13'h4DB: filaimg <= 9'b101110110;
      13'h4DC: filaimg <= 9'b101110110;
      13'h4DD: filaimg <= 9'b101110110;
      13'h4DE: filaimg <= 9'b101110110;
      13'h4DF: filaimg <= 9'b101110110;
      13'h4E0: filaimg <= 9'b101110110;
      13'h4E1: filaimg <= 9'b101110110;
      13'h4E2: filaimg <= 9'b101110110;
      13'h4E3: filaimg <= 9'b101110110;
      13'h4E4: filaimg <= 9'b101110110;
      13'h4E5: filaimg <= 9'b101110110;
      13'h4E6: filaimg <= 9'b101110110;
      13'h4E7: filaimg <= 9'b101110110;
      13'h4E8: filaimg <= 9'b101110110;
      13'h4E9: filaimg <= 9'b101110110;
      13'h4EA: filaimg <= 9'b101110110;
      13'h4EB: filaimg <= 9'b101110110;
      13'h4EC: filaimg <= 9'b101110110;
      13'h4ED: filaimg <= 9'b101110110;
      13'h4EE: filaimg <= 9'b101110110;
      13'h4EF: filaimg <= 9'b101110110;
      13'h4F0: filaimg <= 9'b101110110;
      13'h4F1: filaimg <= 9'b101110110;
      13'h4F2: filaimg <= 9'b101110110;
      13'h4F3: filaimg <= 9'b101110110;
      13'h4F4: filaimg <= 9'b101110110;
      13'h4F5: filaimg <= 9'b101110110;
      13'h4F6: filaimg <= 9'b101110110;
      13'h4F7: filaimg <= 9'b101110110;
      13'h4F8: filaimg <= 9'b101110110;
      13'h4F9: filaimg <= 9'b101110110;
      13'h4FA: filaimg <= 9'b101110110;
      13'h4FB: filaimg <= 9'b101110110;
      13'h4FC: filaimg <= 9'b101110110;
      13'h4FD: filaimg <= 9'b101110110;
      13'h4FE: filaimg <= 9'b101110110;
      13'h4FF: filaimg <= 9'b101110110;
      13'h500: filaimg <= 9'b101110110;
      13'h501: filaimg <= 9'b101110110;
      13'h502: filaimg <= 9'b101110110;
      13'h503: filaimg <= 9'b101110110;
      13'h504: filaimg <= 9'b101110110;
      13'h505: filaimg <= 9'b101110110;
      13'h506: filaimg <= 9'b101110110;
      13'h507: filaimg <= 9'b101110110;
      13'h508: filaimg <= 9'b101110110;
      13'h509: filaimg <= 9'b101110110;
      13'h50A: filaimg <= 9'b101110110;
      13'h50B: filaimg <= 9'b101110110;
      13'h50C: filaimg <= 9'b101110110;
      13'h50D: filaimg <= 9'b101110110;
      13'h50E: filaimg <= 9'b101110110;
      13'h50F: filaimg <= 9'b101110110;
      13'h510: filaimg <= 9'b101110110;
      13'h511: filaimg <= 9'b101110110;
      13'h512: filaimg <= 9'b101110110;
      13'h513: filaimg <= 9'b101110110;
      13'h514: filaimg <= 9'b101110110;
      13'h515: filaimg <= 9'b101110110;
      13'h516: filaimg <= 9'b101110110;
      13'h517: filaimg <= 9'b101110110;
      13'h518: filaimg <= 9'b101110110;
      13'h519: filaimg <= 9'b101110110;
      13'h51A: filaimg <= 9'b101110110;
      13'h51B: filaimg <= 9'b101110110;
      13'h51C: filaimg <= 9'b101110110;
      13'h51D: filaimg <= 9'b101110110;
      13'h51E: filaimg <= 9'b101110110;
      13'h51F: filaimg <= 9'b101110110;
      13'h520: filaimg <= 9'b101110110;
      13'h521: filaimg <= 9'b101110110;
      13'h522: filaimg <= 9'b101110110;
      13'h523: filaimg <= 9'b101110110;
      13'h524: filaimg <= 9'b101110110;
      13'h525: filaimg <= 9'b101110110;
      13'h526: filaimg <= 9'b101110110;
      13'h527: filaimg <= 9'b101110110;
      13'h528: filaimg <= 9'b101110110;
      13'h529: filaimg <= 9'b101110110;
      13'h52A: filaimg <= 9'b101110110;
      13'h52B: filaimg <= 9'b101110110;
      13'h52C: filaimg <= 9'b101110110;
      13'h52D: filaimg <= 9'b101110110;
      13'h52E: filaimg <= 9'b101110110;
      13'h52F: filaimg <= 9'b101110110;
      13'h530: filaimg <= 9'b101110110;
      13'h531: filaimg <= 9'b101110110;
      13'h532: filaimg <= 9'b101110110;
      13'h533: filaimg <= 9'b101110110;
      13'h534: filaimg <= 9'b101110110;
      13'h535: filaimg <= 9'b101110110;
      13'h536: filaimg <= 9'b101110110;
      13'h537: filaimg <= 9'b101110110;
      13'h538: filaimg <= 9'b101110110;
      13'h539: filaimg <= 9'b101110110;
      13'h53A: filaimg <= 9'b101110110;
      13'h53B: filaimg <= 9'b101110110;
      13'h53C: filaimg <= 9'b101110110;
      13'h53D: filaimg <= 9'b101110110;
      13'h53E: filaimg <= 9'b101110110;
      13'h53F: filaimg <= 9'b101110110;
      13'h540: filaimg <= 9'b101110110;
      13'h541: filaimg <= 9'b101110110;
      13'h542: filaimg <= 9'b101110110;
      13'h543: filaimg <= 9'b101110110;
      13'h544: filaimg <= 9'b101110110;
      13'h545: filaimg <= 9'b101110110;
      13'h546: filaimg <= 9'b101110110;
      13'h547: filaimg <= 9'b101110110;
      13'h548: filaimg <= 9'b101110110;
      13'h549: filaimg <= 9'b101110110;
      13'h54A: filaimg <= 9'b101110110;
      13'h54B: filaimg <= 9'b101110110;
      13'h54C: filaimg <= 9'b101110110;
      13'h54D: filaimg <= 9'b101110110;
      13'h54E: filaimg <= 9'b101110110;
      13'h54F: filaimg <= 9'b101110110;
      13'h550: filaimg <= 9'b101110110;
      13'h551: filaimg <= 9'b101110110;
      13'h552: filaimg <= 9'b101110110;
      13'h553: filaimg <= 9'b101110110;
      13'h554: filaimg <= 9'b101110110;
      13'h555: filaimg <= 9'b101110110;
      13'h556: filaimg <= 9'b101110110;
      13'h557: filaimg <= 9'b101110110;
      13'h558: filaimg <= 9'b101110110;
      13'h559: filaimg <= 9'b101110110;
      13'h55A: filaimg <= 9'b101110110;
      13'h55B: filaimg <= 9'b101110110;
      13'h55C: filaimg <= 9'b101110110;
      13'h55D: filaimg <= 9'b101110110;
      13'h55E: filaimg <= 9'b101110110;
      13'h55F: filaimg <= 9'b101110110;
      13'h560: filaimg <= 9'b101110110;
      13'h561: filaimg <= 9'b101110110;
      13'h562: filaimg <= 9'b101110110;
      13'h563: filaimg <= 9'b101110110;
      13'h564: filaimg <= 9'b101110110;
      13'h565: filaimg <= 9'b101110110;
      13'h566: filaimg <= 9'b101110110;
      13'h567: filaimg <= 9'b101110110;
      13'h568: filaimg <= 9'b101110110;
      13'h569: filaimg <= 9'b101110110;
      13'h56A: filaimg <= 9'b101110110;
      13'h56B: filaimg <= 9'b101110110;
      13'h56C: filaimg <= 9'b101110110;
      13'h56D: filaimg <= 9'b101110110;
      13'h56E: filaimg <= 9'b101110110;
      13'h56F: filaimg <= 9'b101110110;
      13'h570: filaimg <= 9'b101110110;
      13'h571: filaimg <= 9'b101110110;
      13'h572: filaimg <= 9'b101110110;
      13'h573: filaimg <= 9'b101110110;
      13'h574: filaimg <= 9'b101110110;
      13'h575: filaimg <= 9'b101110110;
      13'h576: filaimg <= 9'b101110110;
      13'h577: filaimg <= 9'b101110110;
      13'h578: filaimg <= 9'b101110110;
      13'h579: filaimg <= 9'b101110110;
      13'h57A: filaimg <= 9'b101110110;
      13'h57B: filaimg <= 9'b101110110;
      13'h57C: filaimg <= 9'b101110110;
      13'h57D: filaimg <= 9'b101110110;
      13'h57E: filaimg <= 9'b101110110;
      13'h57F: filaimg <= 9'b101110110;
      13'h580: filaimg <= 9'b101110110;
      13'h581: filaimg <= 9'b101110110;
      13'h582: filaimg <= 9'b101110110;
      13'h583: filaimg <= 9'b101110110;
      13'h584: filaimg <= 9'b101110110;
      13'h585: filaimg <= 9'b101110110;
      13'h586: filaimg <= 9'b101110110;
      13'h587: filaimg <= 9'b101110110;
      13'h588: filaimg <= 9'b101110110;
      13'h589: filaimg <= 9'b101110110;
      13'h58A: filaimg <= 9'b101110110;
      13'h58B: filaimg <= 9'b101110110;
      13'h58C: filaimg <= 9'b101110110;
      13'h58D: filaimg <= 9'b101110110;
      13'h58E: filaimg <= 9'b101110110;
      13'h58F: filaimg <= 9'b101110110;
      13'h590: filaimg <= 9'b101110110;
      13'h591: filaimg <= 9'b101110110;
      13'h592: filaimg <= 9'b101110110;
      13'h593: filaimg <= 9'b101110110;
      13'h594: filaimg <= 9'b101110110;
      13'h595: filaimg <= 9'b101110110;
      13'h596: filaimg <= 9'b101110110;
      13'h597: filaimg <= 9'b101110110;
      13'h598: filaimg <= 9'b101110110;
      13'h599: filaimg <= 9'b101110110;
      13'h59A: filaimg <= 9'b101110110;
      13'h59B: filaimg <= 9'b101110110;
      13'h59C: filaimg <= 9'b101110110;
      13'h59D: filaimg <= 9'b101110110;
      13'h59E: filaimg <= 9'b101110110;
      13'h59F: filaimg <= 9'b101110110;
      13'h5A0: filaimg <= 9'b101110110;
      13'h5A1: filaimg <= 9'b101110110;
      13'h5A2: filaimg <= 9'b101110110;
      13'h5A3: filaimg <= 9'b101110110;
      13'h5A4: filaimg <= 9'b101110110;
      13'h5A5: filaimg <= 9'b101110110;
      13'h5A6: filaimg <= 9'b101110110;
      13'h5A7: filaimg <= 9'b101110110;
      13'h5A8: filaimg <= 9'b101110110;
      13'h5A9: filaimg <= 9'b101110110;
      13'h5AA: filaimg <= 9'b101110110;
      13'h5AB: filaimg <= 9'b101110110;
      13'h5AC: filaimg <= 9'b101110110;
      13'h5AD: filaimg <= 9'b101110110;
      13'h5AE: filaimg <= 9'b101110110;
      13'h5AF: filaimg <= 9'b101110110;
      13'h5B0: filaimg <= 9'b101110110;
      13'h5B1: filaimg <= 9'b101110110;
      13'h5B2: filaimg <= 9'b101110110;
      13'h5B3: filaimg <= 9'b101110110;
      13'h5B4: filaimg <= 9'b101110110;
      13'h5B5: filaimg <= 9'b101110110;
      13'h5B6: filaimg <= 9'b101110110;
      13'h5B7: filaimg <= 9'b101110110;
      13'h5B8: filaimg <= 9'b101110110;
      13'h5B9: filaimg <= 9'b101110110;
      13'h5BA: filaimg <= 9'b101110110;
      13'h5BB: filaimg <= 9'b101110110;
      13'h5BC: filaimg <= 9'b101110110;
      13'h5BD: filaimg <= 9'b101110110;
      13'h5BE: filaimg <= 9'b101110110;
      13'h5BF: filaimg <= 9'b101110110;
      13'h5C0: filaimg <= 9'b101110110;
      13'h5C1: filaimg <= 9'b101110110;
      13'h5C2: filaimg <= 9'b101110110;
      13'h5C3: filaimg <= 9'b101110110;
      13'h5C4: filaimg <= 9'b101110110;
      13'h5C5: filaimg <= 9'b101110110;
      13'h5C6: filaimg <= 9'b101110110;
      13'h5C7: filaimg <= 9'b101110110;
      13'h5C8: filaimg <= 9'b101110110;
      13'h5C9: filaimg <= 9'b101110110;
      13'h5CA: filaimg <= 9'b101110110;
      13'h5CB: filaimg <= 9'b101110110;
      13'h5CC: filaimg <= 9'b101110110;
      13'h5CD: filaimg <= 9'b101110110;
      13'h5CE: filaimg <= 9'b101110110;
      13'h5CF: filaimg <= 9'b101110110;
      13'h5D0: filaimg <= 9'b101110110;
      13'h5D1: filaimg <= 9'b101110110;
      13'h5D2: filaimg <= 9'b101110110;
      13'h5D3: filaimg <= 9'b101110110;
      13'h5D4: filaimg <= 9'b101110110;
      13'h5D5: filaimg <= 9'b101110110;
      13'h5D6: filaimg <= 9'b101110110;
      13'h5D7: filaimg <= 9'b101110110;
      13'h5D8: filaimg <= 9'b101110110;
      13'h5D9: filaimg <= 9'b101110110;
      13'h5DA: filaimg <= 9'b101110110;
      13'h5DB: filaimg <= 9'b101110110;
      13'h5DC: filaimg <= 9'b101110110;
      13'h5DD: filaimg <= 9'b101110110;
      13'h5DE: filaimg <= 9'b101110110;
      13'h5DF: filaimg <= 9'b101110110;
      13'h5E0: filaimg <= 9'b101110110;
      13'h5E1: filaimg <= 9'b101110110;
      13'h5E2: filaimg <= 9'b101110110;
      13'h5E3: filaimg <= 9'b101110110;
      13'h5E4: filaimg <= 9'b101110110;
      13'h5E5: filaimg <= 9'b101110110;
      13'h5E6: filaimg <= 9'b101110110;
      13'h5E7: filaimg <= 9'b101110110;
      13'h5E8: filaimg <= 9'b101110110;
      13'h5E9: filaimg <= 9'b101110110;
      13'h5EA: filaimg <= 9'b101110110;
      13'h5EB: filaimg <= 9'b101110110;
      13'h5EC: filaimg <= 9'b101110110;
      13'h5ED: filaimg <= 9'b101110110;
      13'h5EE: filaimg <= 9'b101110110;
      13'h5EF: filaimg <= 9'b101110110;
      13'h5F0: filaimg <= 9'b101110110;
      13'h5F1: filaimg <= 9'b101110110;
      13'h5F2: filaimg <= 9'b101110110;
      13'h5F3: filaimg <= 9'b101110110;
      13'h5F4: filaimg <= 9'b101110110;
      13'h5F5: filaimg <= 9'b101110110;
      13'h5F6: filaimg <= 9'b101110110;
      13'h5F7: filaimg <= 9'b101110110;
      13'h5F8: filaimg <= 9'b101110110;
      13'h5F9: filaimg <= 9'b101110110;
      13'h5FA: filaimg <= 9'b101110110;
      13'h5FB: filaimg <= 9'b101110110;
      13'h5FC: filaimg <= 9'b101110110;
      13'h5FD: filaimg <= 9'b101110110;
      13'h5FE: filaimg <= 9'b101110110;
      13'h5FF: filaimg <= 9'b101110110;
      13'h600: filaimg <= 9'b101110110;
      13'h601: filaimg <= 9'b101110110;
      13'h602: filaimg <= 9'b101110110;
      13'h603: filaimg <= 9'b101110110;
      13'h604: filaimg <= 9'b101110110;
      13'h605: filaimg <= 9'b101110110;
      13'h606: filaimg <= 9'b101110110;
      13'h607: filaimg <= 9'b101110110;
      13'h608: filaimg <= 9'b101110110;
      13'h609: filaimg <= 9'b101110110;
      13'h60A: filaimg <= 9'b101110110;
      13'h60B: filaimg <= 9'b101110110;
      13'h60C: filaimg <= 9'b101110110;
      13'h60D: filaimg <= 9'b101110110;
      13'h60E: filaimg <= 9'b101110110;
      13'h60F: filaimg <= 9'b101110110;
      13'h610: filaimg <= 9'b101110110;
      13'h611: filaimg <= 9'b101110110;
      13'h612: filaimg <= 9'b101110110;
      13'h613: filaimg <= 9'b101110110;
      13'h614: filaimg <= 9'b101110110;
      13'h615: filaimg <= 9'b101110110;
      13'h616: filaimg <= 9'b101110110;
      13'h617: filaimg <= 9'b101110110;
      13'h618: filaimg <= 9'b101110110;
      13'h619: filaimg <= 9'b101110110;
      13'h61A: filaimg <= 9'b101110110;
      13'h61B: filaimg <= 9'b101110110;
      13'h61C: filaimg <= 9'b101110110;
      13'h61D: filaimg <= 9'b101110110;
      13'h61E: filaimg <= 9'b101110110;
      13'h61F: filaimg <= 9'b101110110;
      13'h620: filaimg <= 9'b101110110;
      13'h621: filaimg <= 9'b101110110;
      13'h622: filaimg <= 9'b101110110;
      13'h623: filaimg <= 9'b101110110;
      13'h624: filaimg <= 9'b101110110;
      13'h625: filaimg <= 9'b101110110;
      13'h626: filaimg <= 9'b101110110;
      13'h627: filaimg <= 9'b101110110;
      13'h628: filaimg <= 9'b101110110;
      13'h629: filaimg <= 9'b101110110;
      13'h62A: filaimg <= 9'b101110110;
      13'h62B: filaimg <= 9'b101110110;
      13'h62C: filaimg <= 9'b101110110;
      13'h62D: filaimg <= 9'b101110110;
      13'h62E: filaimg <= 9'b101110110;
      13'h62F: filaimg <= 9'b101110110;
      13'h630: filaimg <= 9'b101110110;
      13'h631: filaimg <= 9'b101110110;
      13'h632: filaimg <= 9'b101110110;
      13'h633: filaimg <= 9'b101110110;
      13'h634: filaimg <= 9'b101110110;
      13'h635: filaimg <= 9'b101110110;
      13'h636: filaimg <= 9'b101110110;
      13'h637: filaimg <= 9'b101110110;
      13'h638: filaimg <= 9'b101110110;
      13'h639: filaimg <= 9'b101110110;
      13'h63A: filaimg <= 9'b101110110;
      13'h63B: filaimg <= 9'b101110110;
      13'h63C: filaimg <= 9'b101110110;
      13'h63D: filaimg <= 9'b101110110;
      13'h63E: filaimg <= 9'b101110110;
      13'h63F: filaimg <= 9'b101110110;
      13'h640: filaimg <= 9'b101110110;
      13'h641: filaimg <= 9'b101110110;
      13'h642: filaimg <= 9'b101110110;
      13'h643: filaimg <= 9'b101110110;
      13'h644: filaimg <= 9'b101110110;
      13'h645: filaimg <= 9'b101110110;
      13'h646: filaimg <= 9'b101110110;
      13'h647: filaimg <= 9'b101110110;
      13'h648: filaimg <= 9'b101110110;
      13'h649: filaimg <= 9'b101110110;
      13'h64A: filaimg <= 9'b101110110;
      13'h64B: filaimg <= 9'b101110110;
      13'h64C: filaimg <= 9'b101110110;
      13'h64D: filaimg <= 9'b101110110;
      13'h64E: filaimg <= 9'b101110110;
      13'h64F: filaimg <= 9'b101110110;
      13'h650: filaimg <= 9'b101110110;
      13'h651: filaimg <= 9'b101110110;
      13'h652: filaimg <= 9'b101110110;
      13'h653: filaimg <= 9'b101110110;
      13'h654: filaimg <= 9'b101110110;
      13'h655: filaimg <= 9'b101110110;
      13'h656: filaimg <= 9'b101110110;
      13'h657: filaimg <= 9'b101110110;
      13'h658: filaimg <= 9'b101110110;
      13'h659: filaimg <= 9'b101110110;
      13'h65A: filaimg <= 9'b101110110;
      13'h65B: filaimg <= 9'b101110110;
      13'h65C: filaimg <= 9'b101110110;
      13'h65D: filaimg <= 9'b101110110;
      13'h65E: filaimg <= 9'b101110110;
      13'h65F: filaimg <= 9'b101110110;
      13'h660: filaimg <= 9'b101110110;
      13'h661: filaimg <= 9'b101110110;
      13'h662: filaimg <= 9'b101110110;
      13'h663: filaimg <= 9'b101110110;
      13'h664: filaimg <= 9'b101110110;
      13'h665: filaimg <= 9'b101110110;
      13'h666: filaimg <= 9'b101110110;
      13'h667: filaimg <= 9'b101110110;
      13'h668: filaimg <= 9'b101110110;
      13'h669: filaimg <= 9'b101110110;
      13'h66A: filaimg <= 9'b101110110;
      13'h66B: filaimg <= 9'b101110110;
      13'h66C: filaimg <= 9'b101110110;
      13'h66D: filaimg <= 9'b101110110;
      13'h66E: filaimg <= 9'b101110110;
      13'h66F: filaimg <= 9'b101110110;
      13'h670: filaimg <= 9'b101110110;
      13'h671: filaimg <= 9'b101110110;
      13'h672: filaimg <= 9'b101110110;
      13'h673: filaimg <= 9'b101110110;
      13'h674: filaimg <= 9'b101110110;
      13'h675: filaimg <= 9'b101110110;
      13'h676: filaimg <= 9'b101110110;
      13'h677: filaimg <= 9'b101110110;
      13'h678: filaimg <= 9'b101110110;
      13'h679: filaimg <= 9'b101110110;
      13'h67A: filaimg <= 9'b101110110;
      13'h67B: filaimg <= 9'b101110110;
      13'h67C: filaimg <= 9'b101110110;
      13'h67D: filaimg <= 9'b101110110;
      13'h67E: filaimg <= 9'b101110110;
      13'h67F: filaimg <= 9'b101110110;
      13'h680: filaimg <= 9'b101110110;
      13'h681: filaimg <= 9'b101110110;
      13'h682: filaimg <= 9'b101110110;
      13'h683: filaimg <= 9'b101110110;
      13'h684: filaimg <= 9'b101110110;
      13'h685: filaimg <= 9'b101110110;
      13'h686: filaimg <= 9'b101110110;
      13'h687: filaimg <= 9'b101110110;
      13'h688: filaimg <= 9'b101110110;
      13'h689: filaimg <= 9'b101110110;
      13'h68A: filaimg <= 9'b101110110;
      13'h68B: filaimg <= 9'b101110110;
      13'h68C: filaimg <= 9'b101110110;
      13'h68D: filaimg <= 9'b101110110;
      13'h68E: filaimg <= 9'b101110110;
      13'h68F: filaimg <= 9'b101110110;
      13'h690: filaimg <= 9'b101110110;
      13'h691: filaimg <= 9'b101110110;
      13'h692: filaimg <= 9'b101110110;
      13'h693: filaimg <= 9'b101110110;
      13'h694: filaimg <= 9'b101110110;
      13'h695: filaimg <= 9'b101110110;
      13'h696: filaimg <= 9'b101110110;
      13'h697: filaimg <= 9'b101110110;
      13'h698: filaimg <= 9'b101110110;
      13'h699: filaimg <= 9'b101110110;
      13'h69A: filaimg <= 9'b101110110;
      13'h69B: filaimg <= 9'b101110110;
      13'h69C: filaimg <= 9'b101110110;
      13'h69D: filaimg <= 9'b101110110;
      13'h69E: filaimg <= 9'b101110110;
      13'h69F: filaimg <= 9'b101110110;
      13'h6A0: filaimg <= 9'b101110110;
      13'h6A1: filaimg <= 9'b101110110;
      13'h6A2: filaimg <= 9'b101110110;
      13'h6A3: filaimg <= 9'b101110110;
      13'h6A4: filaimg <= 9'b101110110;
      13'h6A5: filaimg <= 9'b101110110;
      13'h6A6: filaimg <= 9'b101110110;
      13'h6A7: filaimg <= 9'b101110110;
      13'h6A8: filaimg <= 9'b101110110;
      13'h6A9: filaimg <= 9'b101110110;
      13'h6AA: filaimg <= 9'b101110110;
      13'h6AB: filaimg <= 9'b101110110;
      13'h6AC: filaimg <= 9'b101110110;
      13'h6AD: filaimg <= 9'b101110110;
      13'h6AE: filaimg <= 9'b101110110;
      13'h6AF: filaimg <= 9'b101110110;
      13'h6B0: filaimg <= 9'b101110110;
      13'h6B1: filaimg <= 9'b101110110;
      13'h6B2: filaimg <= 9'b101110110;
      13'h6B3: filaimg <= 9'b101110110;
      13'h6B4: filaimg <= 9'b101110110;
      13'h6B5: filaimg <= 9'b101110110;
      13'h6B6: filaimg <= 9'b101110110;
      13'h6B7: filaimg <= 9'b101110110;
      13'h6B8: filaimg <= 9'b101110110;
      13'h6B9: filaimg <= 9'b101110110;
      13'h6BA: filaimg <= 9'b101110110;
      13'h6BB: filaimg <= 9'b101110110;
      13'h6BC: filaimg <= 9'b101110110;
      13'h6BD: filaimg <= 9'b101110110;
      13'h6BE: filaimg <= 9'b101110110;
      13'h6BF: filaimg <= 9'b101110110;
      13'h6C0: filaimg <= 9'b101110110;
      13'h6C1: filaimg <= 9'b101110110;
      13'h6C2: filaimg <= 9'b101110110;
      13'h6C3: filaimg <= 9'b101110110;
      13'h6C4: filaimg <= 9'b101110110;
      13'h6C5: filaimg <= 9'b101110110;
      13'h6C6: filaimg <= 9'b101110110;
      13'h6C7: filaimg <= 9'b101110110;
      13'h6C8: filaimg <= 9'b101110110;
      13'h6C9: filaimg <= 9'b101110110;
      13'h6CA: filaimg <= 9'b101110110;
      13'h6CB: filaimg <= 9'b101110110;
      13'h6CC: filaimg <= 9'b101110110;
      13'h6CD: filaimg <= 9'b101110110;
      13'h6CE: filaimg <= 9'b101110110;
      13'h6CF: filaimg <= 9'b101110110;
      13'h6D0: filaimg <= 9'b101110110;
      13'h6D1: filaimg <= 9'b101110110;
      13'h6D2: filaimg <= 9'b101110110;
      13'h6D3: filaimg <= 9'b101110110;
      13'h6D4: filaimg <= 9'b101110110;
      13'h6D5: filaimg <= 9'b101110110;
      13'h6D6: filaimg <= 9'b101110110;
      13'h6D7: filaimg <= 9'b101110110;
      13'h6D8: filaimg <= 9'b101110110;
      13'h6D9: filaimg <= 9'b101110110;
      13'h6DA: filaimg <= 9'b101110110;
      13'h6DB: filaimg <= 9'b101110110;
      13'h6DC: filaimg <= 9'b101110110;
      13'h6DD: filaimg <= 9'b101110110;
      13'h6DE: filaimg <= 9'b101110110;
      13'h6DF: filaimg <= 9'b101110110;
      13'h6E0: filaimg <= 9'b101110110;
      13'h6E1: filaimg <= 9'b101110110;
      13'h6E2: filaimg <= 9'b101110110;
      13'h6E3: filaimg <= 9'b101110110;
      13'h6E4: filaimg <= 9'b101110110;
      13'h6E5: filaimg <= 9'b101110110;
      13'h6E6: filaimg <= 9'b101110110;
      13'h6E7: filaimg <= 9'b101110110;
      13'h6E8: filaimg <= 9'b101110110;
      13'h6E9: filaimg <= 9'b101110110;
      13'h6EA: filaimg <= 9'b101110110;
      13'h6EB: filaimg <= 9'b101110110;
      13'h6EC: filaimg <= 9'b101110110;
      13'h6ED: filaimg <= 9'b101110110;
      13'h6EE: filaimg <= 9'b101110110;
      13'h6EF: filaimg <= 9'b101110110;
      13'h6F0: filaimg <= 9'b101110110;
      13'h6F1: filaimg <= 9'b101110110;
      13'h6F2: filaimg <= 9'b101110110;
      13'h6F3: filaimg <= 9'b101110110;
      13'h6F4: filaimg <= 9'b101110110;
      13'h6F5: filaimg <= 9'b111000000;
      13'h6F6: filaimg <= 9'b111000000;
      13'h6F7: filaimg <= 9'b111000000;
      13'h6F8: filaimg <= 9'b111000000;
      13'h6F9: filaimg <= 9'b111000000;
      13'h6FA: filaimg <= 9'b111000000;
      13'h6FB: filaimg <= 9'b111000000;
      13'h6FC: filaimg <= 9'b111000000;
      13'h6FD: filaimg <= 9'b111000000;
      13'h6FE: filaimg <= 9'b111000000;
      13'h6FF: filaimg <= 9'b111000000;
      13'h700: filaimg <= 9'b111000000;
      13'h701: filaimg <= 9'b111000000;
      13'h702: filaimg <= 9'b111000000;
      13'h703: filaimg <= 9'b111000000;
      13'h704: filaimg <= 9'b111000000;
      13'h705: filaimg <= 9'b111000000;
      13'h706: filaimg <= 9'b111000000;
      13'h707: filaimg <= 9'b111000000;
      13'h708: filaimg <= 9'b111000000;
      13'h709: filaimg <= 9'b111000000;
      13'h70A: filaimg <= 9'b111000000;
      13'h70B: filaimg <= 9'b101110110;
      13'h70C: filaimg <= 9'b101110110;
      13'h70D: filaimg <= 9'b101110110;
      13'h70E: filaimg <= 9'b101110110;
      13'h70F: filaimg <= 9'b101110110;
      13'h710: filaimg <= 9'b101110110;
      13'h711: filaimg <= 9'b101110110;
      13'h712: filaimg <= 9'b101110110;
      13'h713: filaimg <= 9'b101110110;
      13'h714: filaimg <= 9'b101110110;
      13'h715: filaimg <= 9'b101110110;
      13'h716: filaimg <= 9'b101110110;
      13'h717: filaimg <= 9'b101110110;
      13'h718: filaimg <= 9'b101110110;
      13'h719: filaimg <= 9'b101110110;
      13'h71A: filaimg <= 9'b101110110;
      13'h71B: filaimg <= 9'b101110110;
      13'h71C: filaimg <= 9'b101110110;
      13'h71D: filaimg <= 9'b101110110;
      13'h71E: filaimg <= 9'b101110110;
      13'h71F: filaimg <= 9'b101110110;
      13'h720: filaimg <= 9'b101110110;
      13'h721: filaimg <= 9'b101110110;
      13'h722: filaimg <= 9'b101110110;
      13'h723: filaimg <= 9'b101110110;
      13'h724: filaimg <= 9'b101110110;
      13'h725: filaimg <= 9'b101110110;
      13'h726: filaimg <= 9'b101110110;
      13'h727: filaimg <= 9'b101110110;
      13'h728: filaimg <= 9'b101110110;
      13'h729: filaimg <= 9'b101110110;
      13'h72A: filaimg <= 9'b101110110;
      13'h72B: filaimg <= 9'b101110110;
      13'h72C: filaimg <= 9'b101110110;
      13'h72D: filaimg <= 9'b101110110;
      13'h72E: filaimg <= 9'b101110110;
      13'h72F: filaimg <= 9'b101110110;
      13'h730: filaimg <= 9'b101110110;
      13'h731: filaimg <= 9'b101110110;
      13'h732: filaimg <= 9'b101110110;
      13'h733: filaimg <= 9'b101110110;
      13'h734: filaimg <= 9'b101110110;
      13'h735: filaimg <= 9'b101110110;
      13'h736: filaimg <= 9'b101110110;
      13'h737: filaimg <= 9'b101110110;
      13'h738: filaimg <= 9'b101110110;
      13'h739: filaimg <= 9'b101110110;
      13'h73A: filaimg <= 9'b101110110;
      13'h73B: filaimg <= 9'b101110110;
      13'h73C: filaimg <= 9'b101110110;
      13'h73D: filaimg <= 9'b101110110;
      13'h73E: filaimg <= 9'b101110110;
      13'h73F: filaimg <= 9'b101110110;
      13'h740: filaimg <= 9'b101110110;
      13'h741: filaimg <= 9'b101110110;
      13'h742: filaimg <= 9'b101110110;
      13'h743: filaimg <= 9'b101110110;
      13'h744: filaimg <= 9'b101110110;
      13'h745: filaimg <= 9'b111000000;
      13'h746: filaimg <= 9'b111000000;
      13'h747: filaimg <= 9'b111000000;
      13'h748: filaimg <= 9'b111000000;
      13'h749: filaimg <= 9'b111000000;
      13'h74A: filaimg <= 9'b111000000;
      13'h74B: filaimg <= 9'b111000000;
      13'h74C: filaimg <= 9'b111000000;
      13'h74D: filaimg <= 9'b111000000;
      13'h74E: filaimg <= 9'b111000000;
      13'h74F: filaimg <= 9'b111000000;
      13'h750: filaimg <= 9'b111000000;
      13'h751: filaimg <= 9'b111000000;
      13'h752: filaimg <= 9'b111000000;
      13'h753: filaimg <= 9'b111000000;
      13'h754: filaimg <= 9'b111000000;
      13'h755: filaimg <= 9'b111000000;
      13'h756: filaimg <= 9'b111000000;
      13'h757: filaimg <= 9'b111000000;
      13'h758: filaimg <= 9'b111000000;
      13'h759: filaimg <= 9'b111000000;
      13'h75A: filaimg <= 9'b111000000;
      13'h75B: filaimg <= 9'b101110110;
      13'h75C: filaimg <= 9'b101110110;
      13'h75D: filaimg <= 9'b101110110;
      13'h75E: filaimg <= 9'b101110110;
      13'h75F: filaimg <= 9'b101110110;
      13'h760: filaimg <= 9'b101110110;
      13'h761: filaimg <= 9'b101110110;
      13'h762: filaimg <= 9'b101110110;
      13'h763: filaimg <= 9'b101110110;
      13'h764: filaimg <= 9'b101110110;
      13'h765: filaimg <= 9'b101110110;
      13'h766: filaimg <= 9'b101110110;
      13'h767: filaimg <= 9'b101110110;
      13'h768: filaimg <= 9'b101110110;
      13'h769: filaimg <= 9'b101110110;
      13'h76A: filaimg <= 9'b101110110;
      13'h76B: filaimg <= 9'b101110110;
      13'h76C: filaimg <= 9'b101110110;
      13'h76D: filaimg <= 9'b101110110;
      13'h76E: filaimg <= 9'b101110110;
      13'h76F: filaimg <= 9'b101110110;
      13'h770: filaimg <= 9'b101110110;
      13'h771: filaimg <= 9'b101110110;
      13'h772: filaimg <= 9'b101110110;
      13'h773: filaimg <= 9'b101110110;
      13'h774: filaimg <= 9'b101110110;
      13'h775: filaimg <= 9'b101110110;
      13'h776: filaimg <= 9'b101110110;
      13'h777: filaimg <= 9'b101110110;
      13'h778: filaimg <= 9'b101110110;
      13'h779: filaimg <= 9'b101110110;
      13'h77A: filaimg <= 9'b101110110;
      13'h77B: filaimg <= 9'b101110110;
      13'h77C: filaimg <= 9'b101110110;
      13'h77D: filaimg <= 9'b101110110;
      13'h77E: filaimg <= 9'b101110110;
      13'h77F: filaimg <= 9'b101110110;
      13'h780: filaimg <= 9'b101110110;
      13'h781: filaimg <= 9'b101110110;
      13'h782: filaimg <= 9'b101110110;
      13'h783: filaimg <= 9'b101110110;
      13'h784: filaimg <= 9'b101110110;
      13'h785: filaimg <= 9'b101110110;
      13'h786: filaimg <= 9'b101110110;
      13'h787: filaimg <= 9'b101110110;
      13'h788: filaimg <= 9'b101110110;
      13'h789: filaimg <= 9'b101110110;
      13'h78A: filaimg <= 9'b101110110;
      13'h78B: filaimg <= 9'b101110110;
      13'h78C: filaimg <= 9'b101110110;
      13'h78D: filaimg <= 9'b101110110;
      13'h78E: filaimg <= 9'b101110110;
      13'h78F: filaimg <= 9'b101110110;
      13'h790: filaimg <= 9'b101110110;
      13'h791: filaimg <= 9'b101110110;
      13'h792: filaimg <= 9'b101110110;
      13'h793: filaimg <= 9'b101110110;
      13'h794: filaimg <= 9'b101110110;
      13'h795: filaimg <= 9'b111000000;
      13'h796: filaimg <= 9'b111000000;
      13'h797: filaimg <= 9'b111000000;
      13'h798: filaimg <= 9'b111000000;
      13'h799: filaimg <= 9'b111000000;
      13'h79A: filaimg <= 9'b111000000;
      13'h79B: filaimg <= 9'b111000000;
      13'h79C: filaimg <= 9'b111000000;
      13'h79D: filaimg <= 9'b111000000;
      13'h79E: filaimg <= 9'b111000000;
      13'h79F: filaimg <= 9'b111000000;
      13'h7A0: filaimg <= 9'b111000000;
      13'h7A1: filaimg <= 9'b111000000;
      13'h7A2: filaimg <= 9'b111000000;
      13'h7A3: filaimg <= 9'b111000000;
      13'h7A4: filaimg <= 9'b111000000;
      13'h7A5: filaimg <= 9'b111000000;
      13'h7A6: filaimg <= 9'b111000000;
      13'h7A7: filaimg <= 9'b111000000;
      13'h7A8: filaimg <= 9'b111000000;
      13'h7A9: filaimg <= 9'b111000000;
      13'h7AA: filaimg <= 9'b111000000;
      13'h7AB: filaimg <= 9'b101110110;
      13'h7AC: filaimg <= 9'b101110110;
      13'h7AD: filaimg <= 9'b101110110;
      13'h7AE: filaimg <= 9'b101110110;
      13'h7AF: filaimg <= 9'b101110110;
      13'h7B0: filaimg <= 9'b101110110;
      13'h7B1: filaimg <= 9'b101110110;
      13'h7B2: filaimg <= 9'b101110110;
      13'h7B3: filaimg <= 9'b101110110;
      13'h7B4: filaimg <= 9'b101110110;
      13'h7B5: filaimg <= 9'b101110110;
      13'h7B6: filaimg <= 9'b101110110;
      13'h7B7: filaimg <= 9'b101110110;
      13'h7B8: filaimg <= 9'b101110110;
      13'h7B9: filaimg <= 9'b101110110;
      13'h7BA: filaimg <= 9'b101110110;
      13'h7BB: filaimg <= 9'b101110110;
      13'h7BC: filaimg <= 9'b101110110;
      13'h7BD: filaimg <= 9'b101110110;
      13'h7BE: filaimg <= 9'b101110110;
      13'h7BF: filaimg <= 9'b101110110;
      13'h7C0: filaimg <= 9'b101110110;
      13'h7C1: filaimg <= 9'b101110110;
      13'h7C2: filaimg <= 9'b101110110;
      13'h7C3: filaimg <= 9'b101110110;
      13'h7C4: filaimg <= 9'b101110110;
      13'h7C5: filaimg <= 9'b101110110;
      13'h7C6: filaimg <= 9'b101110110;
      13'h7C7: filaimg <= 9'b101110110;
      13'h7C8: filaimg <= 9'b101110110;
      13'h7C9: filaimg <= 9'b101110110;
      13'h7CA: filaimg <= 9'b101110110;
      13'h7CB: filaimg <= 9'b101110110;
      13'h7CC: filaimg <= 9'b101110110;
      13'h7CD: filaimg <= 9'b101110110;
      13'h7CE: filaimg <= 9'b101110110;
      13'h7CF: filaimg <= 9'b101110110;
      13'h7D0: filaimg <= 9'b101110110;
      13'h7D1: filaimg <= 9'b101110110;
      13'h7D2: filaimg <= 9'b101110110;
      13'h7D3: filaimg <= 9'b101110110;
      13'h7D4: filaimg <= 9'b101110110;
      13'h7D5: filaimg <= 9'b101110110;
      13'h7D6: filaimg <= 9'b101110110;
      13'h7D7: filaimg <= 9'b101110110;
      13'h7D8: filaimg <= 9'b101110110;
      13'h7D9: filaimg <= 9'b101110110;
      13'h7DA: filaimg <= 9'b101110110;
      13'h7DB: filaimg <= 9'b101110110;
      13'h7DC: filaimg <= 9'b101110110;
      13'h7DD: filaimg <= 9'b101110110;
      13'h7DE: filaimg <= 9'b101110110;
      13'h7DF: filaimg <= 9'b101110110;
      13'h7E0: filaimg <= 9'b101110110;
      13'h7E1: filaimg <= 9'b101110110;
      13'h7E2: filaimg <= 9'b101110110;
      13'h7E3: filaimg <= 9'b101110110;
      13'h7E4: filaimg <= 9'b101110110;
      13'h7E5: filaimg <= 9'b111000000;
      13'h7E6: filaimg <= 9'b111000000;
      13'h7E7: filaimg <= 9'b111000000;
      13'h7E8: filaimg <= 9'b111000000;
      13'h7E9: filaimg <= 9'b111000000;
      13'h7EA: filaimg <= 9'b111000000;
      13'h7EB: filaimg <= 9'b111000000;
      13'h7EC: filaimg <= 9'b111000000;
      13'h7ED: filaimg <= 9'b111000000;
      13'h7EE: filaimg <= 9'b111000000;
      13'h7EF: filaimg <= 9'b111000000;
      13'h7F0: filaimg <= 9'b111000000;
      13'h7F1: filaimg <= 9'b111000000;
      13'h7F2: filaimg <= 9'b111000000;
      13'h7F3: filaimg <= 9'b111000000;
      13'h7F4: filaimg <= 9'b111000000;
      13'h7F5: filaimg <= 9'b111000000;
      13'h7F6: filaimg <= 9'b111000000;
      13'h7F7: filaimg <= 9'b111000000;
      13'h7F8: filaimg <= 9'b111000000;
      13'h7F9: filaimg <= 9'b111000000;
      13'h7FA: filaimg <= 9'b111000000;
      13'h7FB: filaimg <= 9'b101110110;
      13'h7FC: filaimg <= 9'b101110110;
      13'h7FD: filaimg <= 9'b101110110;
      13'h7FE: filaimg <= 9'b101110110;
      13'h7FF: filaimg <= 9'b101110110;
      13'h800: filaimg <= 9'b101110110;
      13'h801: filaimg <= 9'b101110110;
      13'h802: filaimg <= 9'b101110110;
      13'h803: filaimg <= 9'b101110110;
      13'h804: filaimg <= 9'b101110110;
      13'h805: filaimg <= 9'b101110110;
      13'h806: filaimg <= 9'b101110110;
      13'h807: filaimg <= 9'b101110110;
      13'h808: filaimg <= 9'b101110110;
      13'h809: filaimg <= 9'b101110110;
      13'h80A: filaimg <= 9'b101110110;
      13'h80B: filaimg <= 9'b101110110;
      13'h80C: filaimg <= 9'b101110110;
      13'h80D: filaimg <= 9'b101110110;
      13'h80E: filaimg <= 9'b101110110;
      13'h80F: filaimg <= 9'b101110110;
      13'h810: filaimg <= 9'b101110110;
      13'h811: filaimg <= 9'b101110110;
      13'h812: filaimg <= 9'b101110110;
      13'h813: filaimg <= 9'b101110110;
      13'h814: filaimg <= 9'b101110110;
      13'h815: filaimg <= 9'b101110110;
      13'h816: filaimg <= 9'b101110110;
      13'h817: filaimg <= 9'b101110110;
      13'h818: filaimg <= 9'b101110110;
      13'h819: filaimg <= 9'b101110110;
      13'h81A: filaimg <= 9'b101110110;
      13'h81B: filaimg <= 9'b101110110;
      13'h81C: filaimg <= 9'b101110110;
      13'h81D: filaimg <= 9'b101110110;
      13'h81E: filaimg <= 9'b101110110;
      13'h81F: filaimg <= 9'b101110110;
      13'h820: filaimg <= 9'b101110110;
      13'h821: filaimg <= 9'b101110110;
      13'h822: filaimg <= 9'b101110110;
      13'h823: filaimg <= 9'b101110110;
      13'h824: filaimg <= 9'b101110110;
      13'h825: filaimg <= 9'b101110110;
      13'h826: filaimg <= 9'b101110110;
      13'h827: filaimg <= 9'b101110110;
      13'h828: filaimg <= 9'b101110110;
      13'h829: filaimg <= 9'b101110110;
      13'h82A: filaimg <= 9'b101110110;
      13'h82B: filaimg <= 9'b101110110;
      13'h82C: filaimg <= 9'b101110110;
      13'h82D: filaimg <= 9'b101110110;
      13'h82E: filaimg <= 9'b101110110;
      13'h82F: filaimg <= 9'b101110110;
      13'h830: filaimg <= 9'b101110110;
      13'h831: filaimg <= 9'b101110110;
      13'h832: filaimg <= 9'b101110110;
      13'h833: filaimg <= 9'b101110110;
      13'h834: filaimg <= 9'b101110110;
      13'h835: filaimg <= 9'b111000000;
      13'h836: filaimg <= 9'b111000000;
      13'h837: filaimg <= 9'b111000000;
      13'h838: filaimg <= 9'b111000000;
      13'h839: filaimg <= 9'b111000000;
      13'h83A: filaimg <= 9'b111000000;
      13'h83B: filaimg <= 9'b111000000;
      13'h83C: filaimg <= 9'b111000000;
      13'h83D: filaimg <= 9'b111000000;
      13'h83E: filaimg <= 9'b111000000;
      13'h83F: filaimg <= 9'b111000000;
      13'h840: filaimg <= 9'b111000000;
      13'h841: filaimg <= 9'b111000000;
      13'h842: filaimg <= 9'b111000000;
      13'h843: filaimg <= 9'b111000000;
      13'h844: filaimg <= 9'b111000000;
      13'h845: filaimg <= 9'b111000000;
      13'h846: filaimg <= 9'b111000000;
      13'h847: filaimg <= 9'b111000000;
      13'h848: filaimg <= 9'b111000000;
      13'h849: filaimg <= 9'b111000000;
      13'h84A: filaimg <= 9'b111000000;
      13'h84B: filaimg <= 9'b101110110;
      13'h84C: filaimg <= 9'b101110110;
      13'h84D: filaimg <= 9'b101110110;
      13'h84E: filaimg <= 9'b101110110;
      13'h84F: filaimg <= 9'b101110110;
      13'h850: filaimg <= 9'b101110110;
      13'h851: filaimg <= 9'b101110110;
      13'h852: filaimg <= 9'b101110110;
      13'h853: filaimg <= 9'b101110110;
      13'h854: filaimg <= 9'b101110110;
      13'h855: filaimg <= 9'b101110110;
      13'h856: filaimg <= 9'b101110110;
      13'h857: filaimg <= 9'b101110110;
      13'h858: filaimg <= 9'b101110110;
      13'h859: filaimg <= 9'b101110110;
      13'h85A: filaimg <= 9'b101110110;
      13'h85B: filaimg <= 9'b101110110;
      13'h85C: filaimg <= 9'b101110110;
      13'h85D: filaimg <= 9'b101110110;
      13'h85E: filaimg <= 9'b101110110;
      13'h85F: filaimg <= 9'b101110110;
      13'h860: filaimg <= 9'b101110110;
      13'h861: filaimg <= 9'b101110110;
      13'h862: filaimg <= 9'b101110110;
      13'h863: filaimg <= 9'b101110110;
      13'h864: filaimg <= 9'b101110110;
      13'h865: filaimg <= 9'b101110110;
      13'h866: filaimg <= 9'b101110110;
      13'h867: filaimg <= 9'b101110110;
      13'h868: filaimg <= 9'b101110110;
      13'h869: filaimg <= 9'b101110110;
      13'h86A: filaimg <= 9'b101110110;
      13'h86B: filaimg <= 9'b101110110;
      13'h86C: filaimg <= 9'b101110110;
      13'h86D: filaimg <= 9'b101110110;
      13'h86E: filaimg <= 9'b101110110;
      13'h86F: filaimg <= 9'b101110110;
      13'h870: filaimg <= 9'b101110110;
      13'h871: filaimg <= 9'b101110110;
      13'h872: filaimg <= 9'b101110110;
      13'h873: filaimg <= 9'b101110110;
      13'h874: filaimg <= 9'b101110110;
      13'h875: filaimg <= 9'b101110110;
      13'h876: filaimg <= 9'b101110110;
      13'h877: filaimg <= 9'b101110110;
      13'h878: filaimg <= 9'b101110110;
      13'h879: filaimg <= 9'b101110110;
      13'h87A: filaimg <= 9'b101110110;
      13'h87B: filaimg <= 9'b101110110;
      13'h87C: filaimg <= 9'b101110110;
      13'h87D: filaimg <= 9'b101110110;
      13'h87E: filaimg <= 9'b101110110;
      13'h87F: filaimg <= 9'b101110110;
      13'h880: filaimg <= 9'b101110110;
      13'h881: filaimg <= 9'b101110110;
      13'h882: filaimg <= 9'b101110110;
      13'h883: filaimg <= 9'b101110110;
      13'h884: filaimg <= 9'b101110110;
      13'h885: filaimg <= 9'b111000000;
      13'h886: filaimg <= 9'b111000000;
      13'h887: filaimg <= 9'b111000000;
      13'h888: filaimg <= 9'b111000000;
      13'h889: filaimg <= 9'b111000000;
      13'h88A: filaimg <= 9'b111000000;
      13'h88B: filaimg <= 9'b111000000;
      13'h88C: filaimg <= 9'b111000000;
      13'h88D: filaimg <= 9'b111000000;
      13'h88E: filaimg <= 9'b111000000;
      13'h88F: filaimg <= 9'b111000000;
      13'h890: filaimg <= 9'b111000000;
      13'h891: filaimg <= 9'b111000000;
      13'h892: filaimg <= 9'b111000000;
      13'h893: filaimg <= 9'b111000000;
      13'h894: filaimg <= 9'b111000000;
      13'h895: filaimg <= 9'b111000000;
      13'h896: filaimg <= 9'b111000000;
      13'h897: filaimg <= 9'b111000000;
      13'h898: filaimg <= 9'b111000000;
      13'h899: filaimg <= 9'b111000000;
      13'h89A: filaimg <= 9'b111000000;
      13'h89B: filaimg <= 9'b101110110;
      13'h89C: filaimg <= 9'b101110110;
      13'h89D: filaimg <= 9'b101110110;
      13'h89E: filaimg <= 9'b101110110;
      13'h89F: filaimg <= 9'b101110110;
      13'h8A0: filaimg <= 9'b101110110;
      13'h8A1: filaimg <= 9'b101110110;
      13'h8A2: filaimg <= 9'b101110110;
      13'h8A3: filaimg <= 9'b101110110;
      13'h8A4: filaimg <= 9'b101110110;
      13'h8A5: filaimg <= 9'b101110110;
      13'h8A6: filaimg <= 9'b101110110;
      13'h8A7: filaimg <= 9'b101110110;
      13'h8A8: filaimg <= 9'b101110110;
      13'h8A9: filaimg <= 9'b101110110;
      13'h8AA: filaimg <= 9'b101110110;
      13'h8AB: filaimg <= 9'b101110110;
      13'h8AC: filaimg <= 9'b101110110;
      13'h8AD: filaimg <= 9'b101110110;
      13'h8AE: filaimg <= 9'b101110110;
      13'h8AF: filaimg <= 9'b101110110;
      13'h8B0: filaimg <= 9'b101110110;
      13'h8B1: filaimg <= 9'b101110110;
      13'h8B2: filaimg <= 9'b101110110;
      13'h8B3: filaimg <= 9'b101110110;
      13'h8B4: filaimg <= 9'b101110110;
      13'h8B5: filaimg <= 9'b101110110;
      13'h8B6: filaimg <= 9'b101110110;
      13'h8B7: filaimg <= 9'b101110110;
      13'h8B8: filaimg <= 9'b101110110;
      13'h8B9: filaimg <= 9'b101110110;
      13'h8BA: filaimg <= 9'b101110110;
      13'h8BB: filaimg <= 9'b101110110;
      13'h8BC: filaimg <= 9'b101110110;
      13'h8BD: filaimg <= 9'b101110110;
      13'h8BE: filaimg <= 9'b101110110;
      13'h8BF: filaimg <= 9'b101110110;
      13'h8C0: filaimg <= 9'b101110110;
      13'h8C1: filaimg <= 9'b101110110;
      13'h8C2: filaimg <= 9'b101110110;
      13'h8C3: filaimg <= 9'b101110110;
      13'h8C4: filaimg <= 9'b101110110;
      13'h8C5: filaimg <= 9'b101110110;
      13'h8C6: filaimg <= 9'b101110110;
      13'h8C7: filaimg <= 9'b101110110;
      13'h8C8: filaimg <= 9'b101110110;
      13'h8C9: filaimg <= 9'b101110110;
      13'h8CA: filaimg <= 9'b101110110;
      13'h8CB: filaimg <= 9'b101110110;
      13'h8CC: filaimg <= 9'b101110110;
      13'h8CD: filaimg <= 9'b101110110;
      13'h8CE: filaimg <= 9'b101110110;
      13'h8CF: filaimg <= 9'b101110110;
      13'h8D0: filaimg <= 9'b101110110;
      13'h8D1: filaimg <= 9'b101110110;
      13'h8D2: filaimg <= 9'b101110110;
      13'h8D3: filaimg <= 9'b101110110;
      13'h8D4: filaimg <= 9'b101110110;
      13'h8D5: filaimg <= 9'b111000000;
      13'h8D6: filaimg <= 9'b111000000;
      13'h8D7: filaimg <= 9'b111000000;
      13'h8D8: filaimg <= 9'b111000000;
      13'h8D9: filaimg <= 9'b111000000;
      13'h8DA: filaimg <= 9'b111000000;
      13'h8DB: filaimg <= 9'b111000000;
      13'h8DC: filaimg <= 9'b111000000;
      13'h8DD: filaimg <= 9'b111000000;
      13'h8DE: filaimg <= 9'b111000000;
      13'h8DF: filaimg <= 9'b111000000;
      13'h8E0: filaimg <= 9'b111000000;
      13'h8E1: filaimg <= 9'b111000000;
      13'h8E2: filaimg <= 9'b111000000;
      13'h8E3: filaimg <= 9'b111000000;
      13'h8E4: filaimg <= 9'b111000000;
      13'h8E5: filaimg <= 9'b111000000;
      13'h8E6: filaimg <= 9'b111000000;
      13'h8E7: filaimg <= 9'b111000000;
      13'h8E8: filaimg <= 9'b111000000;
      13'h8E9: filaimg <= 9'b111000000;
      13'h8EA: filaimg <= 9'b111000000;
      13'h8EB: filaimg <= 9'b101110110;
      13'h8EC: filaimg <= 9'b101110110;
      13'h8ED: filaimg <= 9'b101110110;
      13'h8EE: filaimg <= 9'b101110110;
      13'h8EF: filaimg <= 9'b101110110;
      13'h8F0: filaimg <= 9'b101110110;
      13'h8F1: filaimg <= 9'b101110110;
      13'h8F2: filaimg <= 9'b101110110;
      13'h8F3: filaimg <= 9'b101110110;
      13'h8F4: filaimg <= 9'b101110110;
      13'h8F5: filaimg <= 9'b101110110;
      13'h8F6: filaimg <= 9'b101110110;
      13'h8F7: filaimg <= 9'b101110110;
      13'h8F8: filaimg <= 9'b101110110;
      13'h8F9: filaimg <= 9'b101110110;
      13'h8FA: filaimg <= 9'b101110110;
      13'h8FB: filaimg <= 9'b101110110;
      13'h8FC: filaimg <= 9'b101110110;
      13'h8FD: filaimg <= 9'b101110110;
      13'h8FE: filaimg <= 9'b101110110;
      13'h8FF: filaimg <= 9'b101110110;
      13'h900: filaimg <= 9'b101110110;
      13'h901: filaimg <= 9'b101110110;
      13'h902: filaimg <= 9'b101110110;
      13'h903: filaimg <= 9'b101110110;
      13'h904: filaimg <= 9'b101110110;
      13'h905: filaimg <= 9'b101110110;
      13'h906: filaimg <= 9'b101110110;
      13'h907: filaimg <= 9'b101110110;
      13'h908: filaimg <= 9'b101110110;
      13'h909: filaimg <= 9'b101110110;
      13'h90A: filaimg <= 9'b101110110;
      13'h90B: filaimg <= 9'b101110110;
      13'h90C: filaimg <= 9'b101110110;
      13'h90D: filaimg <= 9'b101110110;
      13'h90E: filaimg <= 9'b101110110;
      13'h90F: filaimg <= 9'b101110110;
      13'h910: filaimg <= 9'b101110110;
      13'h911: filaimg <= 9'b101110110;
      13'h912: filaimg <= 9'b101110110;
      13'h913: filaimg <= 9'b101110110;
      13'h914: filaimg <= 9'b101110110;
      13'h915: filaimg <= 9'b101110110;
      13'h916: filaimg <= 9'b101110110;
      13'h917: filaimg <= 9'b101110110;
      13'h918: filaimg <= 9'b101110110;
      13'h919: filaimg <= 9'b101110110;
      13'h91A: filaimg <= 9'b101110110;
      13'h91B: filaimg <= 9'b101110110;
      13'h91C: filaimg <= 9'b101110110;
      13'h91D: filaimg <= 9'b101110110;
      13'h91E: filaimg <= 9'b101110110;
      13'h91F: filaimg <= 9'b101110110;
      13'h920: filaimg <= 9'b101110110;
      13'h921: filaimg <= 9'b101110110;
      13'h922: filaimg <= 9'b101110110;
      13'h923: filaimg <= 9'b101110110;
      13'h924: filaimg <= 9'b101110110;
      13'h925: filaimg <= 9'b111000000;
      13'h926: filaimg <= 9'b111000000;
      13'h927: filaimg <= 9'b111000000;
      13'h928: filaimg <= 9'b111000000;
      13'h929: filaimg <= 9'b111000000;
      13'h92A: filaimg <= 9'b111000000;
      13'h92B: filaimg <= 9'b111000000;
      13'h92C: filaimg <= 9'b111000000;
      13'h92D: filaimg <= 9'b111000000;
      13'h92E: filaimg <= 9'b111000000;
      13'h92F: filaimg <= 9'b111000000;
      13'h930: filaimg <= 9'b111000000;
      13'h931: filaimg <= 9'b111000000;
      13'h932: filaimg <= 9'b111000000;
      13'h933: filaimg <= 9'b111000000;
      13'h934: filaimg <= 9'b111000000;
      13'h935: filaimg <= 9'b111000000;
      13'h936: filaimg <= 9'b111000000;
      13'h937: filaimg <= 9'b111000000;
      13'h938: filaimg <= 9'b111000000;
      13'h939: filaimg <= 9'b111000000;
      13'h93A: filaimg <= 9'b111000000;
      13'h93B: filaimg <= 9'b101110110;
      13'h93C: filaimg <= 9'b101110110;
      13'h93D: filaimg <= 9'b101110110;
      13'h93E: filaimg <= 9'b101110110;
      13'h93F: filaimg <= 9'b101110110;
      13'h940: filaimg <= 9'b101110110;
      13'h941: filaimg <= 9'b101110110;
      13'h942: filaimg <= 9'b101110110;
      13'h943: filaimg <= 9'b101110110;
      13'h944: filaimg <= 9'b101110110;
      13'h945: filaimg <= 9'b101110110;
      13'h946: filaimg <= 9'b101110110;
      13'h947: filaimg <= 9'b101110110;
      13'h948: filaimg <= 9'b101110110;
      13'h949: filaimg <= 9'b101110110;
      13'h94A: filaimg <= 9'b101110110;
      13'h94B: filaimg <= 9'b101110110;
      13'h94C: filaimg <= 9'b101110110;
      13'h94D: filaimg <= 9'b101110110;
      13'h94E: filaimg <= 9'b101110110;
      13'h94F: filaimg <= 9'b101110110;
      13'h950: filaimg <= 9'b101110110;
      13'h951: filaimg <= 9'b101110110;
      13'h952: filaimg <= 9'b101110110;
      13'h953: filaimg <= 9'b101110110;
      13'h954: filaimg <= 9'b101110110;
      13'h955: filaimg <= 9'b101110110;
      13'h956: filaimg <= 9'b101110110;
      13'h957: filaimg <= 9'b101110110;
      13'h958: filaimg <= 9'b101110110;
      13'h959: filaimg <= 9'b101110110;
      13'h95A: filaimg <= 9'b101110110;
      13'h95B: filaimg <= 9'b101110110;
      13'h95C: filaimg <= 9'b101110110;
      13'h95D: filaimg <= 9'b101110110;
      13'h95E: filaimg <= 9'b101110110;
      13'h95F: filaimg <= 9'b101110110;
      13'h960: filaimg <= 9'b101110110;
      13'h961: filaimg <= 9'b101110110;
      13'h962: filaimg <= 9'b101110110;
      13'h963: filaimg <= 9'b101110110;
      13'h964: filaimg <= 9'b101110110;
      13'h965: filaimg <= 9'b101110110;
      13'h966: filaimg <= 9'b101110110;
      13'h967: filaimg <= 9'b101110110;
      13'h968: filaimg <= 9'b101110110;
      13'h969: filaimg <= 9'b101110110;
      13'h96A: filaimg <= 9'b101110110;
      13'h96B: filaimg <= 9'b101110110;
      13'h96C: filaimg <= 9'b101110110;
      13'h96D: filaimg <= 9'b101110110;
      13'h96E: filaimg <= 9'b101110110;
      13'h96F: filaimg <= 9'b101110110;
      13'h970: filaimg <= 9'b101110110;
      13'h971: filaimg <= 9'b101110110;
      13'h972: filaimg <= 9'b101110110;
      13'h973: filaimg <= 9'b101110110;
      13'h974: filaimg <= 9'b101110110;
      13'h975: filaimg <= 9'b111000000;
      13'h976: filaimg <= 9'b111000000;
      13'h977: filaimg <= 9'b111000000;
      13'h978: filaimg <= 9'b111000000;
      13'h979: filaimg <= 9'b111000000;
      13'h97A: filaimg <= 9'b111000000;
      13'h97B: filaimg <= 9'b111000000;
      13'h97C: filaimg <= 9'b111000000;
      13'h97D: filaimg <= 9'b111000000;
      13'h97E: filaimg <= 9'b111000000;
      13'h97F: filaimg <= 9'b111000000;
      13'h980: filaimg <= 9'b111000000;
      13'h981: filaimg <= 9'b111000000;
      13'h982: filaimg <= 9'b111000000;
      13'h983: filaimg <= 9'b111000000;
      13'h984: filaimg <= 9'b111000000;
      13'h985: filaimg <= 9'b111000000;
      13'h986: filaimg <= 9'b111000000;
      13'h987: filaimg <= 9'b111000000;
      13'h988: filaimg <= 9'b111000000;
      13'h989: filaimg <= 9'b111000000;
      13'h98A: filaimg <= 9'b111000000;
      13'h98B: filaimg <= 9'b101110110;
      13'h98C: filaimg <= 9'b101110110;
      13'h98D: filaimg <= 9'b101110110;
      13'h98E: filaimg <= 9'b101110110;
      13'h98F: filaimg <= 9'b101110110;
      13'h990: filaimg <= 9'b101110110;
      13'h991: filaimg <= 9'b101110110;
      13'h992: filaimg <= 9'b101110110;
      13'h993: filaimg <= 9'b101110110;
      13'h994: filaimg <= 9'b101110110;
      13'h995: filaimg <= 9'b101110110;
      13'h996: filaimg <= 9'b101110110;
      13'h997: filaimg <= 9'b101110110;
      13'h998: filaimg <= 9'b101110110;
      13'h999: filaimg <= 9'b101110110;
      13'h99A: filaimg <= 9'b101110110;
      13'h99B: filaimg <= 9'b101110110;
      13'h99C: filaimg <= 9'b101110110;
      13'h99D: filaimg <= 9'b101110110;
      13'h99E: filaimg <= 9'b101110110;
      13'h99F: filaimg <= 9'b101110110;
      13'h9A0: filaimg <= 9'b101110110;
      13'h9A1: filaimg <= 9'b101110110;
      13'h9A2: filaimg <= 9'b101110110;
      13'h9A3: filaimg <= 9'b101110110;
      13'h9A4: filaimg <= 9'b101110110;
      13'h9A5: filaimg <= 9'b101110110;
      13'h9A6: filaimg <= 9'b101110110;
      13'h9A7: filaimg <= 9'b101110110;
      13'h9A8: filaimg <= 9'b101110110;
      13'h9A9: filaimg <= 9'b101110110;
      13'h9AA: filaimg <= 9'b101110110;
      13'h9AB: filaimg <= 9'b101110110;
      13'h9AC: filaimg <= 9'b101110110;
      13'h9AD: filaimg <= 9'b101110110;
      13'h9AE: filaimg <= 9'b101110110;
      13'h9AF: filaimg <= 9'b101110110;
      13'h9B0: filaimg <= 9'b101110110;
      13'h9B1: filaimg <= 9'b101110110;
      13'h9B2: filaimg <= 9'b101110110;
      13'h9B3: filaimg <= 9'b101110110;
      13'h9B4: filaimg <= 9'b101110110;
      13'h9B5: filaimg <= 9'b101110110;
      13'h9B6: filaimg <= 9'b101110110;
      13'h9B7: filaimg <= 9'b101110110;
      13'h9B8: filaimg <= 9'b101110110;
      13'h9B9: filaimg <= 9'b101110110;
      13'h9BA: filaimg <= 9'b101110110;
      13'h9BB: filaimg <= 9'b101110110;
      13'h9BC: filaimg <= 9'b101110110;
      13'h9BD: filaimg <= 9'b101110110;
      13'h9BE: filaimg <= 9'b101110110;
      13'h9BF: filaimg <= 9'b101110110;
      13'h9C0: filaimg <= 9'b101110110;
      13'h9C1: filaimg <= 9'b101110110;
      13'h9C2: filaimg <= 9'b101110110;
      13'h9C3: filaimg <= 9'b101110110;
      13'h9C4: filaimg <= 9'b101110110;
      13'h9C5: filaimg <= 9'b111000000;
      13'h9C6: filaimg <= 9'b111000000;
      13'h9C7: filaimg <= 9'b111000000;
      13'h9C8: filaimg <= 9'b111000000;
      13'h9C9: filaimg <= 9'b111000000;
      13'h9CA: filaimg <= 9'b111000000;
      13'h9CB: filaimg <= 9'b111000000;
      13'h9CC: filaimg <= 9'b111000000;
      13'h9CD: filaimg <= 9'b111000000;
      13'h9CE: filaimg <= 9'b111000000;
      13'h9CF: filaimg <= 9'b111000000;
      13'h9D0: filaimg <= 9'b111000000;
      13'h9D1: filaimg <= 9'b111000000;
      13'h9D2: filaimg <= 9'b111000000;
      13'h9D3: filaimg <= 9'b111000000;
      13'h9D4: filaimg <= 9'b111000000;
      13'h9D5: filaimg <= 9'b111000000;
      13'h9D6: filaimg <= 9'b111000000;
      13'h9D7: filaimg <= 9'b111000000;
      13'h9D8: filaimg <= 9'b111000000;
      13'h9D9: filaimg <= 9'b111000000;
      13'h9DA: filaimg <= 9'b111000000;
      13'h9DB: filaimg <= 9'b101110110;
      13'h9DC: filaimg <= 9'b101110110;
      13'h9DD: filaimg <= 9'b101110110;
      13'h9DE: filaimg <= 9'b101110110;
      13'h9DF: filaimg <= 9'b101110110;
      13'h9E0: filaimg <= 9'b101110110;
      13'h9E1: filaimg <= 9'b101110110;
      13'h9E2: filaimg <= 9'b101110110;
      13'h9E3: filaimg <= 9'b101110110;
      13'h9E4: filaimg <= 9'b101110110;
      13'h9E5: filaimg <= 9'b101110110;
      13'h9E6: filaimg <= 9'b101110110;
      13'h9E7: filaimg <= 9'b101110110;
      13'h9E8: filaimg <= 9'b101110110;
      13'h9E9: filaimg <= 9'b101110110;
      13'h9EA: filaimg <= 9'b101110110;
      13'h9EB: filaimg <= 9'b101110110;
      13'h9EC: filaimg <= 9'b101110110;
      13'h9ED: filaimg <= 9'b101110110;
      13'h9EE: filaimg <= 9'b101110110;
      13'h9EF: filaimg <= 9'b101110110;
      13'h9F0: filaimg <= 9'b101110110;
      13'h9F1: filaimg <= 9'b101110110;
      13'h9F2: filaimg <= 9'b101110110;
      13'h9F3: filaimg <= 9'b101110110;
      13'h9F4: filaimg <= 9'b101110110;
      13'h9F5: filaimg <= 9'b101110110;
      13'h9F6: filaimg <= 9'b101110110;
      13'h9F7: filaimg <= 9'b101110110;
      13'h9F8: filaimg <= 9'b101110110;
      13'h9F9: filaimg <= 9'b101110110;
      13'h9FA: filaimg <= 9'b101110110;
      13'h9FB: filaimg <= 9'b101110110;
      13'h9FC: filaimg <= 9'b101110110;
      13'h9FD: filaimg <= 9'b101110110;
      13'h9FE: filaimg <= 9'b101110110;
      13'h9FF: filaimg <= 9'b101110110;
      13'hA00: filaimg <= 9'b101110110;
      13'hA01: filaimg <= 9'b101110110;
      13'hA02: filaimg <= 9'b101110110;
      13'hA03: filaimg <= 9'b101110110;
      13'hA04: filaimg <= 9'b101110110;
      13'hA05: filaimg <= 9'b101110110;
      13'hA06: filaimg <= 9'b101110110;
      13'hA07: filaimg <= 9'b101110110;
      13'hA08: filaimg <= 9'b101110110;
      13'hA09: filaimg <= 9'b101110110;
      13'hA0A: filaimg <= 9'b101110110;
      13'hA0B: filaimg <= 9'b101110110;
      13'hA0C: filaimg <= 9'b101110110;
      13'hA0D: filaimg <= 9'b101110110;
      13'hA0E: filaimg <= 9'b101110110;
      13'hA0F: filaimg <= 9'b101110110;
      13'hA10: filaimg <= 9'b101110110;
      13'hA11: filaimg <= 9'b101110110;
      13'hA12: filaimg <= 9'b101110110;
      13'hA13: filaimg <= 9'b101110110;
      13'hA14: filaimg <= 9'b101110110;
      13'hA15: filaimg <= 9'b111000000;
      13'hA16: filaimg <= 9'b111000000;
      13'hA17: filaimg <= 9'b111000000;
      13'hA18: filaimg <= 9'b111000000;
      13'hA19: filaimg <= 9'b111000000;
      13'hA1A: filaimg <= 9'b111000000;
      13'hA1B: filaimg <= 9'b111000000;
      13'hA1C: filaimg <= 9'b111000000;
      13'hA1D: filaimg <= 9'b111000000;
      13'hA1E: filaimg <= 9'b111000000;
      13'hA1F: filaimg <= 9'b111000000;
      13'hA20: filaimg <= 9'b111000000;
      13'hA21: filaimg <= 9'b111000000;
      13'hA22: filaimg <= 9'b111000000;
      13'hA23: filaimg <= 9'b111000000;
      13'hA24: filaimg <= 9'b111000000;
      13'hA25: filaimg <= 9'b111000000;
      13'hA26: filaimg <= 9'b111000000;
      13'hA27: filaimg <= 9'b111000000;
      13'hA28: filaimg <= 9'b111000000;
      13'hA29: filaimg <= 9'b111000000;
      13'hA2A: filaimg <= 9'b111000000;
      13'hA2B: filaimg <= 9'b101110110;
      13'hA2C: filaimg <= 9'b101110110;
      13'hA2D: filaimg <= 9'b101110110;
      13'hA2E: filaimg <= 9'b101110110;
      13'hA2F: filaimg <= 9'b101110110;
      13'hA30: filaimg <= 9'b101110110;
      13'hA31: filaimg <= 9'b101110110;
      13'hA32: filaimg <= 9'b101110110;
      13'hA33: filaimg <= 9'b101110110;
      13'hA34: filaimg <= 9'b101110110;
      13'hA35: filaimg <= 9'b101110110;
      13'hA36: filaimg <= 9'b101110110;
      13'hA37: filaimg <= 9'b101110110;
      13'hA38: filaimg <= 9'b101110110;
      13'hA39: filaimg <= 9'b101110110;
      13'hA3A: filaimg <= 9'b101110110;
      13'hA3B: filaimg <= 9'b101110110;
      13'hA3C: filaimg <= 9'b101110110;
      13'hA3D: filaimg <= 9'b101110110;
      13'hA3E: filaimg <= 9'b101110110;
      13'hA3F: filaimg <= 9'b101110110;
      13'hA40: filaimg <= 9'b101110110;
      13'hA41: filaimg <= 9'b101110110;
      13'hA42: filaimg <= 9'b101110110;
      13'hA43: filaimg <= 9'b101110110;
      13'hA44: filaimg <= 9'b101110110;
      13'hA45: filaimg <= 9'b101110110;
      13'hA46: filaimg <= 9'b101110110;
      13'hA47: filaimg <= 9'b101110110;
      13'hA48: filaimg <= 9'b101110110;
      13'hA49: filaimg <= 9'b101110110;
      13'hA4A: filaimg <= 9'b101110110;
      13'hA4B: filaimg <= 9'b101110110;
      13'hA4C: filaimg <= 9'b101110110;
      13'hA4D: filaimg <= 9'b101110110;
      13'hA4E: filaimg <= 9'b101110110;
      13'hA4F: filaimg <= 9'b101110110;
      13'hA50: filaimg <= 9'b101110110;
      13'hA51: filaimg <= 9'b101110110;
      13'hA52: filaimg <= 9'b101110110;
      13'hA53: filaimg <= 9'b101110110;
      13'hA54: filaimg <= 9'b101110110;
      13'hA55: filaimg <= 9'b101110110;
      13'hA56: filaimg <= 9'b101110110;
      13'hA57: filaimg <= 9'b101110110;
      13'hA58: filaimg <= 9'b101110110;
      13'hA59: filaimg <= 9'b101110110;
      13'hA5A: filaimg <= 9'b101110110;
      13'hA5B: filaimg <= 9'b101110110;
      13'hA5C: filaimg <= 9'b101110110;
      13'hA5D: filaimg <= 9'b101110110;
      13'hA5E: filaimg <= 9'b101110110;
      13'hA5F: filaimg <= 9'b101110110;
      13'hA60: filaimg <= 9'b101110110;
      13'hA61: filaimg <= 9'b101110110;
      13'hA62: filaimg <= 9'b101110110;
      13'hA63: filaimg <= 9'b101110110;
      13'hA64: filaimg <= 9'b101110110;
      13'hA65: filaimg <= 9'b111000000;
      13'hA66: filaimg <= 9'b111000000;
      13'hA67: filaimg <= 9'b111000000;
      13'hA68: filaimg <= 9'b111000000;
      13'hA69: filaimg <= 9'b111000000;
      13'hA6A: filaimg <= 9'b111000000;
      13'hA6B: filaimg <= 9'b111000000;
      13'hA6C: filaimg <= 9'b111000000;
      13'hA6D: filaimg <= 9'b111000000;
      13'hA6E: filaimg <= 9'b111000000;
      13'hA6F: filaimg <= 9'b111000000;
      13'hA70: filaimg <= 9'b111000000;
      13'hA71: filaimg <= 9'b111000000;
      13'hA72: filaimg <= 9'b111000000;
      13'hA73: filaimg <= 9'b111000000;
      13'hA74: filaimg <= 9'b111000000;
      13'hA75: filaimg <= 9'b111000000;
      13'hA76: filaimg <= 9'b111000000;
      13'hA77: filaimg <= 9'b111000000;
      13'hA78: filaimg <= 9'b111000000;
      13'hA79: filaimg <= 9'b111000000;
      13'hA7A: filaimg <= 9'b111000000;
      13'hA7B: filaimg <= 9'b101110110;
      13'hA7C: filaimg <= 9'b101110110;
      13'hA7D: filaimg <= 9'b101110110;
      13'hA7E: filaimg <= 9'b101110110;
      13'hA7F: filaimg <= 9'b101110110;
      13'hA80: filaimg <= 9'b101110110;
      13'hA81: filaimg <= 9'b101110110;
      13'hA82: filaimg <= 9'b101110110;
      13'hA83: filaimg <= 9'b101110110;
      13'hA84: filaimg <= 9'b101110110;
      13'hA85: filaimg <= 9'b101110110;
      13'hA86: filaimg <= 9'b101110110;
      13'hA87: filaimg <= 9'b101110110;
      13'hA88: filaimg <= 9'b101110110;
      13'hA89: filaimg <= 9'b101110110;
      13'hA8A: filaimg <= 9'b101110110;
      13'hA8B: filaimg <= 9'b101110110;
      13'hA8C: filaimg <= 9'b101110110;
      13'hA8D: filaimg <= 9'b101110110;
      13'hA8E: filaimg <= 9'b101110110;
      13'hA8F: filaimg <= 9'b101110110;
      13'hA90: filaimg <= 9'b101110110;
      13'hA91: filaimg <= 9'b101110110;
      13'hA92: filaimg <= 9'b101110110;
      13'hA93: filaimg <= 9'b101110110;
      13'hA94: filaimg <= 9'b101110110;
      13'hA95: filaimg <= 9'b101110110;
      13'hA96: filaimg <= 9'b101110110;
      13'hA97: filaimg <= 9'b101110110;
      13'hA98: filaimg <= 9'b101110110;
      13'hA99: filaimg <= 9'b101110110;
      13'hA9A: filaimg <= 9'b101110110;
      13'hA9B: filaimg <= 9'b101110110;
      13'hA9C: filaimg <= 9'b101110110;
      13'hA9D: filaimg <= 9'b101110110;
      13'hA9E: filaimg <= 9'b101110110;
      13'hA9F: filaimg <= 9'b101110110;
      13'hAA0: filaimg <= 9'b101110110;
      13'hAA1: filaimg <= 9'b101110110;
      13'hAA2: filaimg <= 9'b101110110;
      13'hAA3: filaimg <= 9'b101110110;
      13'hAA4: filaimg <= 9'b101110110;
      13'hAA5: filaimg <= 9'b101110110;
      13'hAA6: filaimg <= 9'b101110110;
      13'hAA7: filaimg <= 9'b101110110;
      13'hAA8: filaimg <= 9'b101110110;
      13'hAA9: filaimg <= 9'b101110110;
      13'hAAA: filaimg <= 9'b101110110;
      13'hAAB: filaimg <= 9'b101110110;
      13'hAAC: filaimg <= 9'b101110110;
      13'hAAD: filaimg <= 9'b101110110;
      13'hAAE: filaimg <= 9'b101110110;
      13'hAAF: filaimg <= 9'b101110110;
      13'hAB0: filaimg <= 9'b101110110;
      13'hAB1: filaimg <= 9'b101110110;
      13'hAB2: filaimg <= 9'b101110110;
      13'hAB3: filaimg <= 9'b101110110;
      13'hAB4: filaimg <= 9'b101110110;
      13'hAB5: filaimg <= 9'b111000000;
      13'hAB6: filaimg <= 9'b111000000;
      13'hAB7: filaimg <= 9'b111000000;
      13'hAB8: filaimg <= 9'b111000000;
      13'hAB9: filaimg <= 9'b111000000;
      13'hABA: filaimg <= 9'b111000000;
      13'hABB: filaimg <= 9'b111000000;
      13'hABC: filaimg <= 9'b111000000;
      13'hABD: filaimg <= 9'b111000000;
      13'hABE: filaimg <= 9'b111000000;
      13'hABF: filaimg <= 9'b111000000;
      13'hAC0: filaimg <= 9'b111000000;
      13'hAC1: filaimg <= 9'b111000000;
      13'hAC2: filaimg <= 9'b111000000;
      13'hAC3: filaimg <= 9'b111000000;
      13'hAC4: filaimg <= 9'b111000000;
      13'hAC5: filaimg <= 9'b111000000;
      13'hAC6: filaimg <= 9'b111000000;
      13'hAC7: filaimg <= 9'b111000000;
      13'hAC8: filaimg <= 9'b111000000;
      13'hAC9: filaimg <= 9'b111000000;
      13'hACA: filaimg <= 9'b111000000;
      13'hACB: filaimg <= 9'b101110110;
      13'hACC: filaimg <= 9'b101110110;
      13'hACD: filaimg <= 9'b101110110;
      13'hACE: filaimg <= 9'b101110110;
      13'hACF: filaimg <= 9'b101110110;
      13'hAD0: filaimg <= 9'b101110110;
      13'hAD1: filaimg <= 9'b101110110;
      13'hAD2: filaimg <= 9'b101110110;
      13'hAD3: filaimg <= 9'b101110110;
      13'hAD4: filaimg <= 9'b101110110;
      13'hAD5: filaimg <= 9'b101110110;
      13'hAD6: filaimg <= 9'b101110110;
      13'hAD7: filaimg <= 9'b101110110;
      13'hAD8: filaimg <= 9'b101110110;
      13'hAD9: filaimg <= 9'b101110110;
      13'hADA: filaimg <= 9'b101110110;
      13'hADB: filaimg <= 9'b101110110;
      13'hADC: filaimg <= 9'b101110110;
      13'hADD: filaimg <= 9'b101110110;
      13'hADE: filaimg <= 9'b101110110;
      13'hADF: filaimg <= 9'b101110110;
      13'hAE0: filaimg <= 9'b101110110;
      13'hAE1: filaimg <= 9'b101110110;
      13'hAE2: filaimg <= 9'b101110110;
      13'hAE3: filaimg <= 9'b101110110;
      13'hAE4: filaimg <= 9'b101110110;
      13'hAE5: filaimg <= 9'b101110110;
      13'hAE6: filaimg <= 9'b101110110;
      13'hAE7: filaimg <= 9'b101110110;
      13'hAE8: filaimg <= 9'b101110110;
      13'hAE9: filaimg <= 9'b101110110;
      13'hAEA: filaimg <= 9'b101110110;
      13'hAEB: filaimg <= 9'b101110110;
      13'hAEC: filaimg <= 9'b101110110;
      13'hAED: filaimg <= 9'b101110110;
      13'hAEE: filaimg <= 9'b101110110;
      13'hAEF: filaimg <= 9'b101110110;
      13'hAF0: filaimg <= 9'b101110110;
      13'hAF1: filaimg <= 9'b101110110;
      13'hAF2: filaimg <= 9'b101110110;
      13'hAF3: filaimg <= 9'b101110110;
      13'hAF4: filaimg <= 9'b101110110;
      13'hAF5: filaimg <= 9'b101110110;
      13'hAF6: filaimg <= 9'b101110110;
      13'hAF7: filaimg <= 9'b101110110;
      13'hAF8: filaimg <= 9'b101110110;
      13'hAF9: filaimg <= 9'b101110110;
      13'hAFA: filaimg <= 9'b101110110;
      13'hAFB: filaimg <= 9'b101110110;
      13'hAFC: filaimg <= 9'b101110110;
      13'hAFD: filaimg <= 9'b101110110;
      13'hAFE: filaimg <= 9'b101110110;
      13'hAFF: filaimg <= 9'b101110110;
      13'hB00: filaimg <= 9'b101110110;
      13'hB01: filaimg <= 9'b101110110;
      13'hB02: filaimg <= 9'b101110110;
      13'hB03: filaimg <= 9'b101110110;
      13'hB04: filaimg <= 9'b101110110;
      13'hB05: filaimg <= 9'b111000000;
      13'hB06: filaimg <= 9'b111000000;
      13'hB07: filaimg <= 9'b111000000;
      13'hB08: filaimg <= 9'b111000000;
      13'hB09: filaimg <= 9'b111000000;
      13'hB0A: filaimg <= 9'b111000000;
      13'hB0B: filaimg <= 9'b111000000;
      13'hB0C: filaimg <= 9'b111000000;
      13'hB0D: filaimg <= 9'b111000000;
      13'hB0E: filaimg <= 9'b111000000;
      13'hB0F: filaimg <= 9'b111000000;
      13'hB10: filaimg <= 9'b111000000;
      13'hB11: filaimg <= 9'b111000000;
      13'hB12: filaimg <= 9'b111000000;
      13'hB13: filaimg <= 9'b111000000;
      13'hB14: filaimg <= 9'b111000000;
      13'hB15: filaimg <= 9'b111000000;
      13'hB16: filaimg <= 9'b111000000;
      13'hB17: filaimg <= 9'b111000000;
      13'hB18: filaimg <= 9'b111000000;
      13'hB19: filaimg <= 9'b111000000;
      13'hB1A: filaimg <= 9'b111000000;
      13'hB1B: filaimg <= 9'b101110110;
      13'hB1C: filaimg <= 9'b101110110;
      13'hB1D: filaimg <= 9'b101110110;
      13'hB1E: filaimg <= 9'b101110110;
      13'hB1F: filaimg <= 9'b101110110;
      13'hB20: filaimg <= 9'b101110110;
      13'hB21: filaimg <= 9'b101110110;
      13'hB22: filaimg <= 9'b101110110;
      13'hB23: filaimg <= 9'b101110110;
      13'hB24: filaimg <= 9'b101110110;
      13'hB25: filaimg <= 9'b101110110;
      13'hB26: filaimg <= 9'b101110110;
      13'hB27: filaimg <= 9'b101110110;
      13'hB28: filaimg <= 9'b101110110;
      13'hB29: filaimg <= 9'b101110110;
      13'hB2A: filaimg <= 9'b101110110;
      13'hB2B: filaimg <= 9'b101110110;
      13'hB2C: filaimg <= 9'b101110110;
      13'hB2D: filaimg <= 9'b101110110;
      13'hB2E: filaimg <= 9'b101110110;
      13'hB2F: filaimg <= 9'b101110110;
      13'hB30: filaimg <= 9'b101110110;
      13'hB31: filaimg <= 9'b101110110;
      13'hB32: filaimg <= 9'b101110110;
      13'hB33: filaimg <= 9'b101110110;
      13'hB34: filaimg <= 9'b101110110;
      13'hB35: filaimg <= 9'b101110110;
      13'hB36: filaimg <= 9'b101110110;
      13'hB37: filaimg <= 9'b101110110;
      13'hB38: filaimg <= 9'b101110110;
      13'hB39: filaimg <= 9'b101110110;
      13'hB3A: filaimg <= 9'b101110110;
      13'hB3B: filaimg <= 9'b101110110;
      13'hB3C: filaimg <= 9'b101110110;
      13'hB3D: filaimg <= 9'b101110110;
      13'hB3E: filaimg <= 9'b101110110;
      13'hB3F: filaimg <= 9'b101110110;
      13'hB40: filaimg <= 9'b101110110;
      13'hB41: filaimg <= 9'b101110110;
      13'hB42: filaimg <= 9'b101110110;
      13'hB43: filaimg <= 9'b101110110;
      13'hB44: filaimg <= 9'b101110110;
      13'hB45: filaimg <= 9'b101110110;
      13'hB46: filaimg <= 9'b101110110;
      13'hB47: filaimg <= 9'b101110110;
      13'hB48: filaimg <= 9'b101110110;
      13'hB49: filaimg <= 9'b101110110;
      13'hB4A: filaimg <= 9'b101110110;
      13'hB4B: filaimg <= 9'b101110110;
      13'hB4C: filaimg <= 9'b101110110;
      13'hB4D: filaimg <= 9'b101110110;
      13'hB4E: filaimg <= 9'b101110110;
      13'hB4F: filaimg <= 9'b101110110;
      13'hB50: filaimg <= 9'b101110110;
      13'hB51: filaimg <= 9'b101110110;
      13'hB52: filaimg <= 9'b101110110;
      13'hB53: filaimg <= 9'b101110110;
      13'hB54: filaimg <= 9'b101110110;
      13'hB55: filaimg <= 9'b111000000;
      13'hB56: filaimg <= 9'b111000000;
      13'hB57: filaimg <= 9'b111000000;
      13'hB58: filaimg <= 9'b111000000;
      13'hB59: filaimg <= 9'b111000000;
      13'hB5A: filaimg <= 9'b111000000;
      13'hB5B: filaimg <= 9'b111000000;
      13'hB5C: filaimg <= 9'b111000000;
      13'hB5D: filaimg <= 9'b111000000;
      13'hB5E: filaimg <= 9'b111000000;
      13'hB5F: filaimg <= 9'b111000000;
      13'hB60: filaimg <= 9'b111000000;
      13'hB61: filaimg <= 9'b111000000;
      13'hB62: filaimg <= 9'b111000000;
      13'hB63: filaimg <= 9'b111000000;
      13'hB64: filaimg <= 9'b111000000;
      13'hB65: filaimg <= 9'b111000000;
      13'hB66: filaimg <= 9'b111000000;
      13'hB67: filaimg <= 9'b111000000;
      13'hB68: filaimg <= 9'b111000000;
      13'hB69: filaimg <= 9'b111000000;
      13'hB6A: filaimg <= 9'b111000000;
      13'hB6B: filaimg <= 9'b101110110;
      13'hB6C: filaimg <= 9'b101110110;
      13'hB6D: filaimg <= 9'b101110110;
      13'hB6E: filaimg <= 9'b101110110;
      13'hB6F: filaimg <= 9'b101110110;
      13'hB70: filaimg <= 9'b101110110;
      13'hB71: filaimg <= 9'b101110110;
      13'hB72: filaimg <= 9'b101110110;
      13'hB73: filaimg <= 9'b101110110;
      13'hB74: filaimg <= 9'b101110110;
      13'hB75: filaimg <= 9'b101110110;
      13'hB76: filaimg <= 9'b101110110;
      13'hB77: filaimg <= 9'b101110110;
      13'hB78: filaimg <= 9'b101110110;
      13'hB79: filaimg <= 9'b101110110;
      13'hB7A: filaimg <= 9'b101110110;
      13'hB7B: filaimg <= 9'b101110110;
      13'hB7C: filaimg <= 9'b101110110;
      13'hB7D: filaimg <= 9'b101110110;
      13'hB7E: filaimg <= 9'b101110110;
      13'hB7F: filaimg <= 9'b101110110;
      13'hB80: filaimg <= 9'b101110110;
      13'hB81: filaimg <= 9'b101110110;
      13'hB82: filaimg <= 9'b101110110;
      13'hB83: filaimg <= 9'b101110110;
      13'hB84: filaimg <= 9'b101110110;
      13'hB85: filaimg <= 9'b101110110;
      13'hB86: filaimg <= 9'b101110110;
      13'hB87: filaimg <= 9'b101110110;
      13'hB88: filaimg <= 9'b101110110;
      13'hB89: filaimg <= 9'b101110110;
      13'hB8A: filaimg <= 9'b101110110;
      13'hB8B: filaimg <= 9'b101110110;
      13'hB8C: filaimg <= 9'b101110110;
      13'hB8D: filaimg <= 9'b101110110;
      13'hB8E: filaimg <= 9'b101110110;
      13'hB8F: filaimg <= 9'b101110110;
      13'hB90: filaimg <= 9'b101110110;
      13'hB91: filaimg <= 9'b101110110;
      13'hB92: filaimg <= 9'b101110110;
      13'hB93: filaimg <= 9'b101110110;
      13'hB94: filaimg <= 9'b101110110;
      13'hB95: filaimg <= 9'b101110110;
      13'hB96: filaimg <= 9'b101110110;
      13'hB97: filaimg <= 9'b101110110;
      13'hB98: filaimg <= 9'b101110110;
      13'hB99: filaimg <= 9'b101110110;
      13'hB9A: filaimg <= 9'b101110110;
      13'hB9B: filaimg <= 9'b101110110;
      13'hB9C: filaimg <= 9'b101110110;
      13'hB9D: filaimg <= 9'b101110110;
      13'hB9E: filaimg <= 9'b101110110;
      13'hB9F: filaimg <= 9'b101110110;
      13'hBA0: filaimg <= 9'b101110110;
      13'hBA1: filaimg <= 9'b101110110;
      13'hBA2: filaimg <= 9'b101110110;
      13'hBA3: filaimg <= 9'b101110110;
      13'hBA4: filaimg <= 9'b101110110;
      13'hBA5: filaimg <= 9'b111000000;
      13'hBA6: filaimg <= 9'b111000000;
      13'hBA7: filaimg <= 9'b111000000;
      13'hBA8: filaimg <= 9'b111000000;
      13'hBA9: filaimg <= 9'b111000000;
      13'hBAA: filaimg <= 9'b111000000;
      13'hBAB: filaimg <= 9'b111000000;
      13'hBAC: filaimg <= 9'b111000000;
      13'hBAD: filaimg <= 9'b111000000;
      13'hBAE: filaimg <= 9'b111000000;
      13'hBAF: filaimg <= 9'b111000000;
      13'hBB0: filaimg <= 9'b111000000;
      13'hBB1: filaimg <= 9'b111000000;
      13'hBB2: filaimg <= 9'b111000000;
      13'hBB3: filaimg <= 9'b111000000;
      13'hBB4: filaimg <= 9'b111000000;
      13'hBB5: filaimg <= 9'b111000000;
      13'hBB6: filaimg <= 9'b111000000;
      13'hBB7: filaimg <= 9'b111000000;
      13'hBB8: filaimg <= 9'b111000000;
      13'hBB9: filaimg <= 9'b111000000;
      13'hBBA: filaimg <= 9'b111000000;
      13'hBBB: filaimg <= 9'b101110110;
      13'hBBC: filaimg <= 9'b101110110;
      13'hBBD: filaimg <= 9'b101110110;
      13'hBBE: filaimg <= 9'b101110110;
      13'hBBF: filaimg <= 9'b101110110;
      13'hBC0: filaimg <= 9'b101110110;
      13'hBC1: filaimg <= 9'b101110110;
      13'hBC2: filaimg <= 9'b101110110;
      13'hBC3: filaimg <= 9'b101110110;
      13'hBC4: filaimg <= 9'b101110110;
      13'hBC5: filaimg <= 9'b101110110;
      13'hBC6: filaimg <= 9'b101110110;
      13'hBC7: filaimg <= 9'b101110110;
      13'hBC8: filaimg <= 9'b101110110;
      13'hBC9: filaimg <= 9'b101110110;
      13'hBCA: filaimg <= 9'b101110110;
      13'hBCB: filaimg <= 9'b101110110;
      13'hBCC: filaimg <= 9'b101110110;
      13'hBCD: filaimg <= 9'b101110110;
      13'hBCE: filaimg <= 9'b101110110;
      13'hBCF: filaimg <= 9'b101110110;
      13'hBD0: filaimg <= 9'b101110110;
      13'hBD1: filaimg <= 9'b101110110;
      13'hBD2: filaimg <= 9'b101110110;
      13'hBD3: filaimg <= 9'b101110110;
      13'hBD4: filaimg <= 9'b101110110;
      13'hBD5: filaimg <= 9'b101110110;
      13'hBD6: filaimg <= 9'b101110110;
      13'hBD7: filaimg <= 9'b101110110;
      13'hBD8: filaimg <= 9'b101110110;
      13'hBD9: filaimg <= 9'b101110110;
      13'hBDA: filaimg <= 9'b101110110;
      13'hBDB: filaimg <= 9'b101110110;
      13'hBDC: filaimg <= 9'b101110110;
      13'hBDD: filaimg <= 9'b101110110;
      13'hBDE: filaimg <= 9'b101110110;
      13'hBDF: filaimg <= 9'b101110110;
      13'hBE0: filaimg <= 9'b101110110;
      13'hBE1: filaimg <= 9'b101110110;
      13'hBE2: filaimg <= 9'b101110110;
      13'hBE3: filaimg <= 9'b101110110;
      13'hBE4: filaimg <= 9'b101110110;
      13'hBE5: filaimg <= 9'b101110110;
      13'hBE6: filaimg <= 9'b101110110;
      13'hBE7: filaimg <= 9'b101110110;
      13'hBE8: filaimg <= 9'b101110110;
      13'hBE9: filaimg <= 9'b101110110;
      13'hBEA: filaimg <= 9'b101110110;
      13'hBEB: filaimg <= 9'b101110110;
      13'hBEC: filaimg <= 9'b101110110;
      13'hBED: filaimg <= 9'b101110110;
      13'hBEE: filaimg <= 9'b101110110;
      13'hBEF: filaimg <= 9'b101110110;
      13'hBF0: filaimg <= 9'b101110110;
      13'hBF1: filaimg <= 9'b101110110;
      13'hBF2: filaimg <= 9'b101110110;
      13'hBF3: filaimg <= 9'b101110110;
      13'hBF4: filaimg <= 9'b101110110;
      13'hBF5: filaimg <= 9'b111000000;
      13'hBF6: filaimg <= 9'b111000000;
      13'hBF7: filaimg <= 9'b111000000;
      13'hBF8: filaimg <= 9'b111000000;
      13'hBF9: filaimg <= 9'b111000000;
      13'hBFA: filaimg <= 9'b111000000;
      13'hBFB: filaimg <= 9'b111000000;
      13'hBFC: filaimg <= 9'b111000000;
      13'hBFD: filaimg <= 9'b111000000;
      13'hBFE: filaimg <= 9'b111000000;
      13'hBFF: filaimg <= 9'b111000000;
      13'hC00: filaimg <= 9'b111000000;
      13'hC01: filaimg <= 9'b111000000;
      13'hC02: filaimg <= 9'b111000000;
      13'hC03: filaimg <= 9'b111000000;
      13'hC04: filaimg <= 9'b111000000;
      13'hC05: filaimg <= 9'b111000000;
      13'hC06: filaimg <= 9'b111000000;
      13'hC07: filaimg <= 9'b111000000;
      13'hC08: filaimg <= 9'b111000000;
      13'hC09: filaimg <= 9'b111000000;
      13'hC0A: filaimg <= 9'b111000000;
      13'hC0B: filaimg <= 9'b101110110;
      13'hC0C: filaimg <= 9'b101110110;
      13'hC0D: filaimg <= 9'b101110110;
      13'hC0E: filaimg <= 9'b101110110;
      13'hC0F: filaimg <= 9'b101110110;
      13'hC10: filaimg <= 9'b101110110;
      13'hC11: filaimg <= 9'b101110110;
      13'hC12: filaimg <= 9'b101110110;
      13'hC13: filaimg <= 9'b101110110;
      13'hC14: filaimg <= 9'b101110110;
      13'hC15: filaimg <= 9'b101110110;
      13'hC16: filaimg <= 9'b101110110;
      13'hC17: filaimg <= 9'b101110110;
      13'hC18: filaimg <= 9'b101110110;
      13'hC19: filaimg <= 9'b101110110;
      13'hC1A: filaimg <= 9'b101110110;
      13'hC1B: filaimg <= 9'b101110110;
      13'hC1C: filaimg <= 9'b101110110;
      13'hC1D: filaimg <= 9'b101110110;
      13'hC1E: filaimg <= 9'b101110110;
      13'hC1F: filaimg <= 9'b101110110;
      13'hC20: filaimg <= 9'b101110110;
      13'hC21: filaimg <= 9'b101110110;
      13'hC22: filaimg <= 9'b101110110;
      13'hC23: filaimg <= 9'b101110110;
      13'hC24: filaimg <= 9'b101110110;
      13'hC25: filaimg <= 9'b101110110;
      13'hC26: filaimg <= 9'b101110110;
      13'hC27: filaimg <= 9'b101110110;
      13'hC28: filaimg <= 9'b101110110;
      13'hC29: filaimg <= 9'b101110110;
      13'hC2A: filaimg <= 9'b101110110;
      13'hC2B: filaimg <= 9'b101110110;
      13'hC2C: filaimg <= 9'b101110110;
      13'hC2D: filaimg <= 9'b101110110;
      13'hC2E: filaimg <= 9'b101110110;
      13'hC2F: filaimg <= 9'b101110110;
      13'hC30: filaimg <= 9'b101110110;
      13'hC31: filaimg <= 9'b101110110;
      13'hC32: filaimg <= 9'b101110110;
      13'hC33: filaimg <= 9'b101110110;
      13'hC34: filaimg <= 9'b101110110;
      13'hC35: filaimg <= 9'b101110110;
      13'hC36: filaimg <= 9'b101110110;
      13'hC37: filaimg <= 9'b101110110;
      13'hC38: filaimg <= 9'b101110110;
      13'hC39: filaimg <= 9'b101110110;
      13'hC3A: filaimg <= 9'b101110110;
      13'hC3B: filaimg <= 9'b101110110;
      13'hC3C: filaimg <= 9'b101110110;
      13'hC3D: filaimg <= 9'b101110110;
      13'hC3E: filaimg <= 9'b101110110;
      13'hC3F: filaimg <= 9'b101110110;
      13'hC40: filaimg <= 9'b101110110;
      13'hC41: filaimg <= 9'b101110110;
      13'hC42: filaimg <= 9'b101110110;
      13'hC43: filaimg <= 9'b101110110;
      13'hC44: filaimg <= 9'b101110110;
      13'hC45: filaimg <= 9'b101110110;
      13'hC46: filaimg <= 9'b101110110;
      13'hC47: filaimg <= 9'b101110110;
      13'hC48: filaimg <= 9'b101110110;
      13'hC49: filaimg <= 9'b101110110;
      13'hC4A: filaimg <= 9'b101110110;
      13'hC4B: filaimg <= 9'b101110110;
      13'hC4C: filaimg <= 9'b101110110;
      13'hC4D: filaimg <= 9'b101110110;
      13'hC4E: filaimg <= 9'b101110110;
      13'hC4F: filaimg <= 9'b101110110;
      13'hC50: filaimg <= 9'b101110110;
      13'hC51: filaimg <= 9'b101110110;
      13'hC52: filaimg <= 9'b101110110;
      13'hC53: filaimg <= 9'b101110110;
      13'hC54: filaimg <= 9'b101110110;
      13'hC55: filaimg <= 9'b101110110;
      13'hC56: filaimg <= 9'b101110110;
      13'hC57: filaimg <= 9'b101110110;
      13'hC58: filaimg <= 9'b101110110;
      13'hC59: filaimg <= 9'b101110110;
      13'hC5A: filaimg <= 9'b101110110;
      13'hC5B: filaimg <= 9'b101110110;
      13'hC5C: filaimg <= 9'b101110110;
      13'hC5D: filaimg <= 9'b101110110;
      13'hC5E: filaimg <= 9'b101110110;
      13'hC5F: filaimg <= 9'b101110110;
      13'hC60: filaimg <= 9'b101110110;
      13'hC61: filaimg <= 9'b101110110;
      13'hC62: filaimg <= 9'b101110110;
      13'hC63: filaimg <= 9'b101110110;
      13'hC64: filaimg <= 9'b101110110;
      13'hC65: filaimg <= 9'b101110110;
      13'hC66: filaimg <= 9'b101110110;
      13'hC67: filaimg <= 9'b101110110;
      13'hC68: filaimg <= 9'b101110110;
      13'hC69: filaimg <= 9'b101110110;
      13'hC6A: filaimg <= 9'b101110110;
      13'hC6B: filaimg <= 9'b101110110;
      13'hC6C: filaimg <= 9'b101110110;
      13'hC6D: filaimg <= 9'b101110110;
      13'hC6E: filaimg <= 9'b101110110;
      13'hC6F: filaimg <= 9'b101110110;
      13'hC70: filaimg <= 9'b101110110;
      13'hC71: filaimg <= 9'b101110110;
      13'hC72: filaimg <= 9'b101110110;
      13'hC73: filaimg <= 9'b101110110;
      13'hC74: filaimg <= 9'b101110110;
      13'hC75: filaimg <= 9'b101110110;
      13'hC76: filaimg <= 9'b101110110;
      13'hC77: filaimg <= 9'b101110110;
      13'hC78: filaimg <= 9'b101110110;
      13'hC79: filaimg <= 9'b101110110;
      13'hC7A: filaimg <= 9'b101110110;
      13'hC7B: filaimg <= 9'b101110110;
      13'hC7C: filaimg <= 9'b101110110;
      13'hC7D: filaimg <= 9'b101110110;
      13'hC7E: filaimg <= 9'b101110110;
      13'hC7F: filaimg <= 9'b101110110;
      13'hC80: filaimg <= 9'b101110110;
      13'hC81: filaimg <= 9'b101110110;
      13'hC82: filaimg <= 9'b101110110;
      13'hC83: filaimg <= 9'b101110110;
      13'hC84: filaimg <= 9'b101110110;
      13'hC85: filaimg <= 9'b101110110;
      13'hC86: filaimg <= 9'b101110110;
      13'hC87: filaimg <= 9'b101110110;
      13'hC88: filaimg <= 9'b101110110;
      13'hC89: filaimg <= 9'b101110110;
      13'hC8A: filaimg <= 9'b101110110;
      13'hC8B: filaimg <= 9'b101110110;
      13'hC8C: filaimg <= 9'b101110110;
      13'hC8D: filaimg <= 9'b101110110;
      13'hC8E: filaimg <= 9'b101110110;
      13'hC8F: filaimg <= 9'b101110110;
      13'hC90: filaimg <= 9'b101110110;
      13'hC91: filaimg <= 9'b101110110;
      13'hC92: filaimg <= 9'b101110110;
      13'hC93: filaimg <= 9'b101110110;
      13'hC94: filaimg <= 9'b101110110;
      13'hC95: filaimg <= 9'b101110110;
      13'hC96: filaimg <= 9'b101110110;
      13'hC97: filaimg <= 9'b101110110;
      13'hC98: filaimg <= 9'b101110110;
      13'hC99: filaimg <= 9'b101110110;
      13'hC9A: filaimg <= 9'b101110110;
      13'hC9B: filaimg <= 9'b101110110;
      13'hC9C: filaimg <= 9'b101110110;
      13'hC9D: filaimg <= 9'b101110110;
      13'hC9E: filaimg <= 9'b101110110;
      13'hC9F: filaimg <= 9'b101110110;
      13'hCA0: filaimg <= 9'b101110110;
      13'hCA1: filaimg <= 9'b101110110;
      13'hCA2: filaimg <= 9'b101110110;
      13'hCA3: filaimg <= 9'b101110110;
      13'hCA4: filaimg <= 9'b101110110;
      13'hCA5: filaimg <= 9'b101110110;
      13'hCA6: filaimg <= 9'b101110110;
      13'hCA7: filaimg <= 9'b101110110;
      13'hCA8: filaimg <= 9'b101110110;
      13'hCA9: filaimg <= 9'b101110110;
      13'hCAA: filaimg <= 9'b101110110;
      13'hCAB: filaimg <= 9'b101110110;
      13'hCAC: filaimg <= 9'b101110110;
      13'hCAD: filaimg <= 9'b101110110;
      13'hCAE: filaimg <= 9'b101110110;
      13'hCAF: filaimg <= 9'b101110110;
      13'hCB0: filaimg <= 9'b101110110;
      13'hCB1: filaimg <= 9'b101110110;
      13'hCB2: filaimg <= 9'b101110110;
      13'hCB3: filaimg <= 9'b101110110;
      13'hCB4: filaimg <= 9'b101110110;
      13'hCB5: filaimg <= 9'b101110110;
      13'hCB6: filaimg <= 9'b101110110;
      13'hCB7: filaimg <= 9'b101110110;
      13'hCB8: filaimg <= 9'b101110110;
      13'hCB9: filaimg <= 9'b101110110;
      13'hCBA: filaimg <= 9'b101110110;
      13'hCBB: filaimg <= 9'b101110110;
      13'hCBC: filaimg <= 9'b101110110;
      13'hCBD: filaimg <= 9'b101110110;
      13'hCBE: filaimg <= 9'b101110110;
      13'hCBF: filaimg <= 9'b101110110;
      13'hCC0: filaimg <= 9'b101110110;
      13'hCC1: filaimg <= 9'b101110110;
      13'hCC2: filaimg <= 9'b101110110;
      13'hCC3: filaimg <= 9'b101110110;
      13'hCC4: filaimg <= 9'b101110110;
      13'hCC5: filaimg <= 9'b101110110;
      13'hCC6: filaimg <= 9'b101110110;
      13'hCC7: filaimg <= 9'b101110110;
      13'hCC8: filaimg <= 9'b101110110;
      13'hCC9: filaimg <= 9'b101110110;
      13'hCCA: filaimg <= 9'b101110110;
      13'hCCB: filaimg <= 9'b101110110;
      13'hCCC: filaimg <= 9'b101110110;
      13'hCCD: filaimg <= 9'b101110110;
      13'hCCE: filaimg <= 9'b101110110;
      13'hCCF: filaimg <= 9'b101110110;
      13'hCD0: filaimg <= 9'b101110110;
      13'hCD1: filaimg <= 9'b101110110;
      13'hCD2: filaimg <= 9'b101110110;
      13'hCD3: filaimg <= 9'b101110110;
      13'hCD4: filaimg <= 9'b101110110;
      13'hCD5: filaimg <= 9'b101110110;
      13'hCD6: filaimg <= 9'b101110110;
      13'hCD7: filaimg <= 9'b101110110;
      13'hCD8: filaimg <= 9'b101110110;
      13'hCD9: filaimg <= 9'b101110110;
      13'hCDA: filaimg <= 9'b101110110;
      13'hCDB: filaimg <= 9'b101110110;
      13'hCDC: filaimg <= 9'b101110110;
      13'hCDD: filaimg <= 9'b101110110;
      13'hCDE: filaimg <= 9'b101110110;
      13'hCDF: filaimg <= 9'b101110110;
      13'hCE0: filaimg <= 9'b101110110;
      13'hCE1: filaimg <= 9'b101110110;
      13'hCE2: filaimg <= 9'b101110110;
      13'hCE3: filaimg <= 9'b101110110;
      13'hCE4: filaimg <= 9'b101110110;
      13'hCE5: filaimg <= 9'b101110110;
      13'hCE6: filaimg <= 9'b101110110;
      13'hCE7: filaimg <= 9'b101110110;
      13'hCE8: filaimg <= 9'b101110110;
      13'hCE9: filaimg <= 9'b101110110;
      13'hCEA: filaimg <= 9'b101110110;
      13'hCEB: filaimg <= 9'b101110110;
      13'hCEC: filaimg <= 9'b101110110;
      13'hCED: filaimg <= 9'b101110110;
      13'hCEE: filaimg <= 9'b101110110;
      13'hCEF: filaimg <= 9'b101110110;
      13'hCF0: filaimg <= 9'b101110110;
      13'hCF1: filaimg <= 9'b101110110;
      13'hCF2: filaimg <= 9'b101110110;
      13'hCF3: filaimg <= 9'b101110110;
      13'hCF4: filaimg <= 9'b101110110;
      13'hCF5: filaimg <= 9'b101110110;
      13'hCF6: filaimg <= 9'b101110110;
      13'hCF7: filaimg <= 9'b101110110;
      13'hCF8: filaimg <= 9'b101110110;
      13'hCF9: filaimg <= 9'b101110110;
      13'hCFA: filaimg <= 9'b101110110;
      13'hCFB: filaimg <= 9'b101110110;
      13'hCFC: filaimg <= 9'b101110110;
      13'hCFD: filaimg <= 9'b101110110;
      13'hCFE: filaimg <= 9'b101110110;
      13'hCFF: filaimg <= 9'b101110110;
      13'hD00: filaimg <= 9'b101110110;
      13'hD01: filaimg <= 9'b101110110;
      13'hD02: filaimg <= 9'b101110110;
      13'hD03: filaimg <= 9'b101110110;
      13'hD04: filaimg <= 9'b101110110;
      13'hD05: filaimg <= 9'b101110110;
      13'hD06: filaimg <= 9'b101110110;
      13'hD07: filaimg <= 9'b101110110;
      13'hD08: filaimg <= 9'b101110110;
      13'hD09: filaimg <= 9'b101110110;
      13'hD0A: filaimg <= 9'b101110110;
      13'hD0B: filaimg <= 9'b101110110;
      13'hD0C: filaimg <= 9'b101110110;
      13'hD0D: filaimg <= 9'b101110110;
      13'hD0E: filaimg <= 9'b101110110;
      13'hD0F: filaimg <= 9'b101110110;
      13'hD10: filaimg <= 9'b101110110;
      13'hD11: filaimg <= 9'b101110110;
      13'hD12: filaimg <= 9'b101110110;
      13'hD13: filaimg <= 9'b101110110;
      13'hD14: filaimg <= 9'b101110110;
      13'hD15: filaimg <= 9'b101110110;
      13'hD16: filaimg <= 9'b101110110;
      13'hD17: filaimg <= 9'b101110110;
      13'hD18: filaimg <= 9'b101110110;
      13'hD19: filaimg <= 9'b101110110;
      13'hD1A: filaimg <= 9'b101110110;
      13'hD1B: filaimg <= 9'b101110110;
      13'hD1C: filaimg <= 9'b101110110;
      13'hD1D: filaimg <= 9'b101110110;
      13'hD1E: filaimg <= 9'b101110110;
      13'hD1F: filaimg <= 9'b101110110;
      13'hD20: filaimg <= 9'b101110110;
      13'hD21: filaimg <= 9'b101110110;
      13'hD22: filaimg <= 9'b101110110;
      13'hD23: filaimg <= 9'b101110110;
      13'hD24: filaimg <= 9'b101110110;
      13'hD25: filaimg <= 9'b101110110;
      13'hD26: filaimg <= 9'b101110110;
      13'hD27: filaimg <= 9'b101110110;
      13'hD28: filaimg <= 9'b101110110;
      13'hD29: filaimg <= 9'b101110110;
      13'hD2A: filaimg <= 9'b101110110;
      13'hD2B: filaimg <= 9'b101110110;
      13'hD2C: filaimg <= 9'b101110110;
      13'hD2D: filaimg <= 9'b101110110;
      13'hD2E: filaimg <= 9'b101110110;
      13'hD2F: filaimg <= 9'b101110110;
      13'hD30: filaimg <= 9'b101110110;
      13'hD31: filaimg <= 9'b101110110;
      13'hD32: filaimg <= 9'b101110110;
      13'hD33: filaimg <= 9'b101110110;
      13'hD34: filaimg <= 9'b101110110;
      13'hD35: filaimg <= 9'b101110110;
      13'hD36: filaimg <= 9'b101110110;
      13'hD37: filaimg <= 9'b101110110;
      13'hD38: filaimg <= 9'b101110110;
      13'hD39: filaimg <= 9'b101110110;
      13'hD3A: filaimg <= 9'b101110110;
      13'hD3B: filaimg <= 9'b101110110;
      13'hD3C: filaimg <= 9'b101110110;
      13'hD3D: filaimg <= 9'b101110110;
      13'hD3E: filaimg <= 9'b101110110;
      13'hD3F: filaimg <= 9'b101110110;
      13'hD40: filaimg <= 9'b101110110;
      13'hD41: filaimg <= 9'b101110110;
      13'hD42: filaimg <= 9'b101110110;
      13'hD43: filaimg <= 9'b101110110;
      13'hD44: filaimg <= 9'b101110110;
      13'hD45: filaimg <= 9'b101110110;
      13'hD46: filaimg <= 9'b101110110;
      13'hD47: filaimg <= 9'b101110110;
      13'hD48: filaimg <= 9'b101110110;
      13'hD49: filaimg <= 9'b101110110;
      13'hD4A: filaimg <= 9'b101110110;
      13'hD4B: filaimg <= 9'b101110110;
      13'hD4C: filaimg <= 9'b101110110;
      13'hD4D: filaimg <= 9'b101110110;
      13'hD4E: filaimg <= 9'b101110110;
      13'hD4F: filaimg <= 9'b101110110;
      13'hD50: filaimg <= 9'b101110110;
      13'hD51: filaimg <= 9'b101110110;
      13'hD52: filaimg <= 9'b101110110;
      13'hD53: filaimg <= 9'b101110110;
      13'hD54: filaimg <= 9'b101110110;
      13'hD55: filaimg <= 9'b101110110;
      13'hD56: filaimg <= 9'b101110110;
      13'hD57: filaimg <= 9'b101110110;
      13'hD58: filaimg <= 9'b101110110;
      13'hD59: filaimg <= 9'b101110110;
      13'hD5A: filaimg <= 9'b101110110;
      13'hD5B: filaimg <= 9'b101110110;
      13'hD5C: filaimg <= 9'b101110110;
      13'hD5D: filaimg <= 9'b101110110;
      13'hD5E: filaimg <= 9'b101110110;
      13'hD5F: filaimg <= 9'b101110110;
      13'hD60: filaimg <= 9'b101110110;
      13'hD61: filaimg <= 9'b101110110;
      13'hD62: filaimg <= 9'b101110110;
      13'hD63: filaimg <= 9'b101110110;
      13'hD64: filaimg <= 9'b101110110;
      13'hD65: filaimg <= 9'b101110110;
      13'hD66: filaimg <= 9'b101110110;
      13'hD67: filaimg <= 9'b101110110;
      13'hD68: filaimg <= 9'b101110110;
      13'hD69: filaimg <= 9'b101110110;
      13'hD6A: filaimg <= 9'b101110110;
      13'hD6B: filaimg <= 9'b101110110;
      13'hD6C: filaimg <= 9'b101110110;
      13'hD6D: filaimg <= 9'b101110110;
      13'hD6E: filaimg <= 9'b101110110;
      13'hD6F: filaimg <= 9'b101110110;
      13'hD70: filaimg <= 9'b101110110;
      13'hD71: filaimg <= 9'b101110110;
      13'hD72: filaimg <= 9'b101110110;
      13'hD73: filaimg <= 9'b101110110;
      13'hD74: filaimg <= 9'b101110110;
      13'hD75: filaimg <= 9'b101110110;
      13'hD76: filaimg <= 9'b101110110;
      13'hD77: filaimg <= 9'b101110110;
      13'hD78: filaimg <= 9'b101110110;
      13'hD79: filaimg <= 9'b101110110;
      13'hD7A: filaimg <= 9'b101110110;
      13'hD7B: filaimg <= 9'b101110110;
      13'hD7C: filaimg <= 9'b101110110;
      13'hD7D: filaimg <= 9'b101110110;
      13'hD7E: filaimg <= 9'b101110110;
      13'hD7F: filaimg <= 9'b101110110;
      13'hD80: filaimg <= 9'b101110110;
      13'hD81: filaimg <= 9'b101110110;
      13'hD82: filaimg <= 9'b101110110;
      13'hD83: filaimg <= 9'b101110110;
      13'hD84: filaimg <= 9'b101110110;
      13'hD85: filaimg <= 9'b101110110;
      13'hD86: filaimg <= 9'b101110110;
      13'hD87: filaimg <= 9'b101110110;
      13'hD88: filaimg <= 9'b101110110;
      13'hD89: filaimg <= 9'b101110110;
      13'hD8A: filaimg <= 9'b101110110;
      13'hD8B: filaimg <= 9'b101110110;
      13'hD8C: filaimg <= 9'b101110110;
      13'hD8D: filaimg <= 9'b101110110;
      13'hD8E: filaimg <= 9'b101110110;
      13'hD8F: filaimg <= 9'b101110110;
      13'hD90: filaimg <= 9'b101110110;
      13'hD91: filaimg <= 9'b101110110;
      13'hD92: filaimg <= 9'b101110110;
      13'hD93: filaimg <= 9'b101110110;
      13'hD94: filaimg <= 9'b101110110;
      13'hD95: filaimg <= 9'b101110110;
      13'hD96: filaimg <= 9'b101110110;
      13'hD97: filaimg <= 9'b101110110;
      13'hD98: filaimg <= 9'b101110110;
      13'hD99: filaimg <= 9'b101110110;
      13'hD9A: filaimg <= 9'b101110110;
      13'hD9B: filaimg <= 9'b101110110;
      13'hD9C: filaimg <= 9'b101110110;
      13'hD9D: filaimg <= 9'b101110110;
      13'hD9E: filaimg <= 9'b101110110;
      13'hD9F: filaimg <= 9'b101110110;
      13'hDA0: filaimg <= 9'b101110110;
      13'hDA1: filaimg <= 9'b101110110;
      13'hDA2: filaimg <= 9'b101110110;
      13'hDA3: filaimg <= 9'b101110110;
      13'hDA4: filaimg <= 9'b101110110;
      13'hDA5: filaimg <= 9'b101110110;
      13'hDA6: filaimg <= 9'b101110110;
      13'hDA7: filaimg <= 9'b101110110;
      13'hDA8: filaimg <= 9'b101110110;
      13'hDA9: filaimg <= 9'b101110110;
      13'hDAA: filaimg <= 9'b101110110;
      13'hDAB: filaimg <= 9'b101110110;
      13'hDAC: filaimg <= 9'b101110110;
      13'hDAD: filaimg <= 9'b101110110;
      13'hDAE: filaimg <= 9'b101110110;
      13'hDAF: filaimg <= 9'b101110110;
      13'hDB0: filaimg <= 9'b101110110;
      13'hDB1: filaimg <= 9'b101110110;
      13'hDB2: filaimg <= 9'b101110110;
      13'hDB3: filaimg <= 9'b101110110;
      13'hDB4: filaimg <= 9'b101110110;
      13'hDB5: filaimg <= 9'b101110110;
      13'hDB6: filaimg <= 9'b101110110;
      13'hDB7: filaimg <= 9'b101110110;
      13'hDB8: filaimg <= 9'b101110110;
      13'hDB9: filaimg <= 9'b101110110;
      13'hDBA: filaimg <= 9'b101110110;
      13'hDBB: filaimg <= 9'b101110110;
      13'hDBC: filaimg <= 9'b101110110;
      13'hDBD: filaimg <= 9'b101110110;
      13'hDBE: filaimg <= 9'b101110110;
      13'hDBF: filaimg <= 9'b101110110;
      13'hDC0: filaimg <= 9'b101110110;
      13'hDC1: filaimg <= 9'b101110110;
      13'hDC2: filaimg <= 9'b101110110;
      13'hDC3: filaimg <= 9'b101110110;
      13'hDC4: filaimg <= 9'b101110110;
      13'hDC5: filaimg <= 9'b101110110;
      13'hDC6: filaimg <= 9'b101110110;
      13'hDC7: filaimg <= 9'b101110110;
      13'hDC8: filaimg <= 9'b101110110;
      13'hDC9: filaimg <= 9'b101110110;
      13'hDCA: filaimg <= 9'b101110110;
      13'hDCB: filaimg <= 9'b101110110;
      13'hDCC: filaimg <= 9'b101110110;
      13'hDCD: filaimg <= 9'b101110110;
      13'hDCE: filaimg <= 9'b101110110;
      13'hDCF: filaimg <= 9'b101110110;
      13'hDD0: filaimg <= 9'b101110110;
      13'hDD1: filaimg <= 9'b101110110;
      13'hDD2: filaimg <= 9'b101110110;
      13'hDD3: filaimg <= 9'b101110110;
      13'hDD4: filaimg <= 9'b101110110;
      13'hDD5: filaimg <= 9'b101110110;
      13'hDD6: filaimg <= 9'b101110110;
      13'hDD7: filaimg <= 9'b101110110;
      13'hDD8: filaimg <= 9'b101110110;
      13'hDD9: filaimg <= 9'b101110110;
      13'hDDA: filaimg <= 9'b101110110;
      13'hDDB: filaimg <= 9'b101110110;
      13'hDDC: filaimg <= 9'b101110110;
      13'hDDD: filaimg <= 9'b101110110;
      13'hDDE: filaimg <= 9'b101110110;
      13'hDDF: filaimg <= 9'b101110110;
      13'hDE0: filaimg <= 9'b101110110;
      13'hDE1: filaimg <= 9'b101110110;
      13'hDE2: filaimg <= 9'b101110110;
      13'hDE3: filaimg <= 9'b101110110;
      13'hDE4: filaimg <= 9'b101110110;
      13'hDE5: filaimg <= 9'b101110110;
      13'hDE6: filaimg <= 9'b101110110;
      13'hDE7: filaimg <= 9'b101110110;
      13'hDE8: filaimg <= 9'b101110110;
      13'hDE9: filaimg <= 9'b101110110;
      13'hDEA: filaimg <= 9'b101110110;
      13'hDEB: filaimg <= 9'b101110110;
      13'hDEC: filaimg <= 9'b101110110;
      13'hDED: filaimg <= 9'b101110110;
      13'hDEE: filaimg <= 9'b101110110;
      13'hDEF: filaimg <= 9'b101110110;
      13'hDF0: filaimg <= 9'b101110110;
      13'hDF1: filaimg <= 9'b101110110;
      13'hDF2: filaimg <= 9'b101110110;
      13'hDF3: filaimg <= 9'b101110110;
      13'hDF4: filaimg <= 9'b101110110;
      13'hDF5: filaimg <= 9'b101110110;
      13'hDF6: filaimg <= 9'b101110110;
      13'hDF7: filaimg <= 9'b101110110;
      13'hDF8: filaimg <= 9'b101110110;
      13'hDF9: filaimg <= 9'b101110110;
      13'hDFA: filaimg <= 9'b101110110;
      13'hDFB: filaimg <= 9'b101110110;
      13'hDFC: filaimg <= 9'b101110110;
      13'hDFD: filaimg <= 9'b101110110;
      13'hDFE: filaimg <= 9'b101110110;
      13'hDFF: filaimg <= 9'b101110110;
      13'hE00: filaimg <= 9'b101110110;
      13'hE01: filaimg <= 9'b101110110;
      13'hE02: filaimg <= 9'b101110110;
      13'hE03: filaimg <= 9'b101110110;
      13'hE04: filaimg <= 9'b101110110;
      13'hE05: filaimg <= 9'b101110110;
      13'hE06: filaimg <= 9'b101110110;
      13'hE07: filaimg <= 9'b101110110;
      13'hE08: filaimg <= 9'b101110110;
      13'hE09: filaimg <= 9'b101110110;
      13'hE0A: filaimg <= 9'b101110110;
      13'hE0B: filaimg <= 9'b101110110;
      13'hE0C: filaimg <= 9'b101110110;
      13'hE0D: filaimg <= 9'b101110110;
      13'hE0E: filaimg <= 9'b101110110;
      13'hE0F: filaimg <= 9'b101110110;
      13'hE10: filaimg <= 9'b101110110;
      13'hE11: filaimg <= 9'b101110110;
      13'hE12: filaimg <= 9'b101110110;
      13'hE13: filaimg <= 9'b101110110;
      13'hE14: filaimg <= 9'b101110110;
      13'hE15: filaimg <= 9'b101110110;
      13'hE16: filaimg <= 9'b101110110;
      13'hE17: filaimg <= 9'b101110110;
      13'hE18: filaimg <= 9'b101110110;
      13'hE19: filaimg <= 9'b101110110;
      13'hE1A: filaimg <= 9'b101110110;
      13'hE1B: filaimg <= 9'b101110110;
      13'hE1C: filaimg <= 9'b101110110;
      13'hE1D: filaimg <= 9'b101110110;
      13'hE1E: filaimg <= 9'b101110110;
      13'hE1F: filaimg <= 9'b101110110;
      13'hE20: filaimg <= 9'b101110110;
      13'hE21: filaimg <= 9'b101110110;
      13'hE22: filaimg <= 9'b101110110;
      13'hE23: filaimg <= 9'b101110110;
      13'hE24: filaimg <= 9'b101110110;
      13'hE25: filaimg <= 9'b101110110;
      13'hE26: filaimg <= 9'b101110110;
      13'hE27: filaimg <= 9'b101110110;
      13'hE28: filaimg <= 9'b101110110;
      13'hE29: filaimg <= 9'b101110110;
      13'hE2A: filaimg <= 9'b101110110;
      13'hE2B: filaimg <= 9'b101110110;
      13'hE2C: filaimg <= 9'b101110110;
      13'hE2D: filaimg <= 9'b101110110;
      13'hE2E: filaimg <= 9'b101110110;
      13'hE2F: filaimg <= 9'b101110110;
      13'hE30: filaimg <= 9'b101110110;
      13'hE31: filaimg <= 9'b101110110;
      13'hE32: filaimg <= 9'b101110110;
      13'hE33: filaimg <= 9'b101110110;
      13'hE34: filaimg <= 9'b101110110;
      13'hE35: filaimg <= 9'b101110110;
      13'hE36: filaimg <= 9'b101110110;
      13'hE37: filaimg <= 9'b101110110;
      13'hE38: filaimg <= 9'b101110110;
      13'hE39: filaimg <= 9'b101110110;
      13'hE3A: filaimg <= 9'b101110110;
      13'hE3B: filaimg <= 9'b101110110;
      13'hE3C: filaimg <= 9'b101110110;
      13'hE3D: filaimg <= 9'b101110110;
      13'hE3E: filaimg <= 9'b101110110;
      13'hE3F: filaimg <= 9'b101110110;
      13'hE40: filaimg <= 9'b101110110;
      13'hE41: filaimg <= 9'b101110110;
      13'hE42: filaimg <= 9'b101110110;
      13'hE43: filaimg <= 9'b101110110;
      13'hE44: filaimg <= 9'b101110110;
      13'hE45: filaimg <= 9'b101110110;
      13'hE46: filaimg <= 9'b101110110;
      13'hE47: filaimg <= 9'b101110110;
      13'hE48: filaimg <= 9'b101110110;
      13'hE49: filaimg <= 9'b101110110;
      13'hE4A: filaimg <= 9'b101110110;
      13'hE4B: filaimg <= 9'b101110110;
      13'hE4C: filaimg <= 9'b101110110;
      13'hE4D: filaimg <= 9'b101110110;
      13'hE4E: filaimg <= 9'b101110110;
      13'hE4F: filaimg <= 9'b101110110;
      13'hE50: filaimg <= 9'b101110110;
      13'hE51: filaimg <= 9'b101110110;
      13'hE52: filaimg <= 9'b101110110;
      13'hE53: filaimg <= 9'b101110110;
      13'hE54: filaimg <= 9'b101110110;
      13'hE55: filaimg <= 9'b101110110;
      13'hE56: filaimg <= 9'b101110110;
      13'hE57: filaimg <= 9'b101110110;
      13'hE58: filaimg <= 9'b101110110;
      13'hE59: filaimg <= 9'b101110110;
      13'hE5A: filaimg <= 9'b101110110;
      13'hE5B: filaimg <= 9'b101110110;
      13'hE5C: filaimg <= 9'b101110110;
      13'hE5D: filaimg <= 9'b101110110;
      13'hE5E: filaimg <= 9'b101110110;
      13'hE5F: filaimg <= 9'b101110110;
      13'hE60: filaimg <= 9'b101110110;
      13'hE61: filaimg <= 9'b101110110;
      13'hE62: filaimg <= 9'b101110110;
      13'hE63: filaimg <= 9'b101110110;
      13'hE64: filaimg <= 9'b101110110;
      13'hE65: filaimg <= 9'b101110110;
      13'hE66: filaimg <= 9'b101110110;
      13'hE67: filaimg <= 9'b101110110;
      13'hE68: filaimg <= 9'b101110110;
      13'hE69: filaimg <= 9'b101110110;
      13'hE6A: filaimg <= 9'b101110110;
      13'hE6B: filaimg <= 9'b101110110;
      13'hE6C: filaimg <= 9'b101110110;
      13'hE6D: filaimg <= 9'b101110110;
      13'hE6E: filaimg <= 9'b101110110;
      13'hE6F: filaimg <= 9'b101110110;
      13'hE70: filaimg <= 9'b101110110;
      13'hE71: filaimg <= 9'b101110110;
      13'hE72: filaimg <= 9'b101110110;
      13'hE73: filaimg <= 9'b101110110;
      13'hE74: filaimg <= 9'b101110110;
      13'hE75: filaimg <= 9'b101110110;
      13'hE76: filaimg <= 9'b101110110;
      13'hE77: filaimg <= 9'b101110110;
      13'hE78: filaimg <= 9'b101110110;
      13'hE79: filaimg <= 9'b101110110;
      13'hE7A: filaimg <= 9'b101110110;
      13'hE7B: filaimg <= 9'b101110110;
      13'hE7C: filaimg <= 9'b101110110;
      13'hE7D: filaimg <= 9'b101110110;
      13'hE7E: filaimg <= 9'b101110110;
      13'hE7F: filaimg <= 9'b101110110;
      13'hE80: filaimg <= 9'b101110110;
      13'hE81: filaimg <= 9'b101110110;
      13'hE82: filaimg <= 9'b101110110;
      13'hE83: filaimg <= 9'b101110110;
      13'hE84: filaimg <= 9'b101110110;
      13'hE85: filaimg <= 9'b101110110;
      13'hE86: filaimg <= 9'b101110110;
      13'hE87: filaimg <= 9'b101110110;
      13'hE88: filaimg <= 9'b101110110;
      13'hE89: filaimg <= 9'b101110110;
      13'hE8A: filaimg <= 9'b101110110;
      13'hE8B: filaimg <= 9'b101110110;
      13'hE8C: filaimg <= 9'b101110110;
      13'hE8D: filaimg <= 9'b101110110;
      13'hE8E: filaimg <= 9'b101110110;
      13'hE8F: filaimg <= 9'b101110110;
      13'hE90: filaimg <= 9'b101110110;
      13'hE91: filaimg <= 9'b101110110;
      13'hE92: filaimg <= 9'b101110110;
      13'hE93: filaimg <= 9'b101110110;
      13'hE94: filaimg <= 9'b101110110;
      13'hE95: filaimg <= 9'b101110110;
      13'hE96: filaimg <= 9'b101110110;
      13'hE97: filaimg <= 9'b101110110;
      13'hE98: filaimg <= 9'b101110110;
      13'hE99: filaimg <= 9'b101110110;
      13'hE9A: filaimg <= 9'b101110110;
      13'hE9B: filaimg <= 9'b101110110;
      13'hE9C: filaimg <= 9'b101110110;
      13'hE9D: filaimg <= 9'b101110110;
      13'hE9E: filaimg <= 9'b101110110;
      13'hE9F: filaimg <= 9'b101110110;
      13'hEA0: filaimg <= 9'b101110110;
      13'hEA1: filaimg <= 9'b101110110;
      13'hEA2: filaimg <= 9'b101110110;
      13'hEA3: filaimg <= 9'b101110110;
      13'hEA4: filaimg <= 9'b101110110;
      13'hEA5: filaimg <= 9'b101110110;
      13'hEA6: filaimg <= 9'b101110110;
      13'hEA7: filaimg <= 9'b101110110;
      13'hEA8: filaimg <= 9'b101110110;
      13'hEA9: filaimg <= 9'b101110110;
      13'hEAA: filaimg <= 9'b101110110;
      13'hEAB: filaimg <= 9'b101110110;
      13'hEAC: filaimg <= 9'b101110110;
      13'hEAD: filaimg <= 9'b101110110;
      13'hEAE: filaimg <= 9'b101110110;
      13'hEAF: filaimg <= 9'b101110110;
      13'hEB0: filaimg <= 9'b101110110;
      13'hEB1: filaimg <= 9'b101110110;
      13'hEB2: filaimg <= 9'b101110110;
      13'hEB3: filaimg <= 9'b101110110;
      13'hEB4: filaimg <= 9'b101110110;
      13'hEB5: filaimg <= 9'b101110110;
      13'hEB6: filaimg <= 9'b101110110;
      13'hEB7: filaimg <= 9'b101110110;
      13'hEB8: filaimg <= 9'b101110110;
      13'hEB9: filaimg <= 9'b101110110;
      13'hEBA: filaimg <= 9'b101110110;
      13'hEBB: filaimg <= 9'b101110110;
      13'hEBC: filaimg <= 9'b101110110;
      13'hEBD: filaimg <= 9'b101110110;
      13'hEBE: filaimg <= 9'b101110110;
      13'hEBF: filaimg <= 9'b101110110;
      13'hEC0: filaimg <= 9'b101110110;
      13'hEC1: filaimg <= 9'b101110110;
      13'hEC2: filaimg <= 9'b101110110;
      13'hEC3: filaimg <= 9'b101110110;
      13'hEC4: filaimg <= 9'b101110110;
      13'hEC5: filaimg <= 9'b101110110;
      13'hEC6: filaimg <= 9'b101110110;
      13'hEC7: filaimg <= 9'b101110110;
      13'hEC8: filaimg <= 9'b101110110;
      13'hEC9: filaimg <= 9'b101110110;
      13'hECA: filaimg <= 9'b101110110;
      13'hECB: filaimg <= 9'b101110110;
      13'hECC: filaimg <= 9'b101110110;
      13'hECD: filaimg <= 9'b101110110;
      13'hECE: filaimg <= 9'b101110110;
      13'hECF: filaimg <= 9'b101110110;
      13'hED0: filaimg <= 9'b101110110;
      13'hED1: filaimg <= 9'b101110110;
      13'hED2: filaimg <= 9'b101110110;
      13'hED3: filaimg <= 9'b101110110;
      13'hED4: filaimg <= 9'b101110110;
      13'hED5: filaimg <= 9'b101110110;
      13'hED6: filaimg <= 9'b101110110;
      13'hED7: filaimg <= 9'b101110110;
      13'hED8: filaimg <= 9'b101110110;
      13'hED9: filaimg <= 9'b101110110;
      13'hEDA: filaimg <= 9'b101110110;
      13'hEDB: filaimg <= 9'b101110110;
      13'hEDC: filaimg <= 9'b101110110;
      13'hEDD: filaimg <= 9'b101110110;
      13'hEDE: filaimg <= 9'b101110110;
      13'hEDF: filaimg <= 9'b101110110;
      13'hEE0: filaimg <= 9'b101110110;
      13'hEE1: filaimg <= 9'b101110110;
      13'hEE2: filaimg <= 9'b101110110;
      13'hEE3: filaimg <= 9'b101110110;
      13'hEE4: filaimg <= 9'b101110110;
      13'hEE5: filaimg <= 9'b101110110;
      13'hEE6: filaimg <= 9'b101110110;
      13'hEE7: filaimg <= 9'b101110110;
      13'hEE8: filaimg <= 9'b101110110;
      13'hEE9: filaimg <= 9'b101110110;
      13'hEEA: filaimg <= 9'b101110110;
      13'hEEB: filaimg <= 9'b101110110;
      13'hEEC: filaimg <= 9'b101110110;
      13'hEED: filaimg <= 9'b101110110;
      13'hEEE: filaimg <= 9'b101110110;
      13'hEEF: filaimg <= 9'b101110110;
      13'hEF0: filaimg <= 9'b101110110;
      13'hEF1: filaimg <= 9'b101110110;
      13'hEF2: filaimg <= 9'b101110110;
      13'hEF3: filaimg <= 9'b101110110;
      13'hEF4: filaimg <= 9'b101110110;
      13'hEF5: filaimg <= 9'b101110110;
      13'hEF6: filaimg <= 9'b101110110;
      13'hEF7: filaimg <= 9'b101110110;
      13'hEF8: filaimg <= 9'b101110110;
      13'hEF9: filaimg <= 9'b101110110;
      13'hEFA: filaimg <= 9'b101110110;
      13'hEFB: filaimg <= 9'b101110110;
      13'hEFC: filaimg <= 9'b101110110;
      13'hEFD: filaimg <= 9'b101110110;
      13'hEFE: filaimg <= 9'b101110110;
      13'hEFF: filaimg <= 9'b101110110;
      13'hF00: filaimg <= 9'b101110110;
      13'hF01: filaimg <= 9'b101110110;
      13'hF02: filaimg <= 9'b101110110;
      13'hF03: filaimg <= 9'b101110110;
      13'hF04: filaimg <= 9'b101110110;
      13'hF05: filaimg <= 9'b101110110;
      13'hF06: filaimg <= 9'b101110110;
      13'hF07: filaimg <= 9'b101110110;
      13'hF08: filaimg <= 9'b101110110;
      13'hF09: filaimg <= 9'b101110110;
      13'hF0A: filaimg <= 9'b101110110;
      13'hF0B: filaimg <= 9'b101110110;
      13'hF0C: filaimg <= 9'b101110110;
      13'hF0D: filaimg <= 9'b101110110;
      13'hF0E: filaimg <= 9'b101110110;
      13'hF0F: filaimg <= 9'b101110110;
      13'hF10: filaimg <= 9'b101110110;
      13'hF11: filaimg <= 9'b101110110;
      13'hF12: filaimg <= 9'b101110110;
      13'hF13: filaimg <= 9'b101110110;
      13'hF14: filaimg <= 9'b101110110;
      13'hF15: filaimg <= 9'b101110110;
      13'hF16: filaimg <= 9'b101110110;
      13'hF17: filaimg <= 9'b101110110;
      13'hF18: filaimg <= 9'b101110110;
      13'hF19: filaimg <= 9'b101110110;
      13'hF1A: filaimg <= 9'b101110110;
      13'hF1B: filaimg <= 9'b101110110;
      13'hF1C: filaimg <= 9'b101110110;
      13'hF1D: filaimg <= 9'b101110110;
      13'hF1E: filaimg <= 9'b101110110;
      13'hF1F: filaimg <= 9'b101110110;
      13'hF20: filaimg <= 9'b101110110;
      13'hF21: filaimg <= 9'b101110110;
      13'hF22: filaimg <= 9'b101110110;
      13'hF23: filaimg <= 9'b101110110;
      13'hF24: filaimg <= 9'b101110110;
      13'hF25: filaimg <= 9'b101110110;
      13'hF26: filaimg <= 9'b101110110;
      13'hF27: filaimg <= 9'b101110110;
      13'hF28: filaimg <= 9'b101110110;
      13'hF29: filaimg <= 9'b101110110;
      13'hF2A: filaimg <= 9'b101110110;
      13'hF2B: filaimg <= 9'b101110110;
      13'hF2C: filaimg <= 9'b101110110;
      13'hF2D: filaimg <= 9'b101110110;
      13'hF2E: filaimg <= 9'b101110110;
      13'hF2F: filaimg <= 9'b101110110;
      13'hF30: filaimg <= 9'b101110110;
      13'hF31: filaimg <= 9'b101110110;
      13'hF32: filaimg <= 9'b101110110;
      13'hF33: filaimg <= 9'b101110110;
      13'hF34: filaimg <= 9'b101110110;
      13'hF35: filaimg <= 9'b101110110;
      13'hF36: filaimg <= 9'b101110110;
      13'hF37: filaimg <= 9'b101110110;
      13'hF38: filaimg <= 9'b101110110;
      13'hF39: filaimg <= 9'b101110110;
      13'hF3A: filaimg <= 9'b101110110;
      13'hF3B: filaimg <= 9'b101110110;
      13'hF3C: filaimg <= 9'b101110110;
      13'hF3D: filaimg <= 9'b101110110;
      13'hF3E: filaimg <= 9'b101110110;
      13'hF3F: filaimg <= 9'b101110110;
      13'hF40: filaimg <= 9'b101110110;
      13'hF41: filaimg <= 9'b101110110;
      13'hF42: filaimg <= 9'b101110110;
      13'hF43: filaimg <= 9'b101110110;
      13'hF44: filaimg <= 9'b101110110;
      13'hF45: filaimg <= 9'b101110110;
      13'hF46: filaimg <= 9'b101110110;
      13'hF47: filaimg <= 9'b101110110;
      13'hF48: filaimg <= 9'b101110110;
      13'hF49: filaimg <= 9'b101110110;
      13'hF4A: filaimg <= 9'b101110110;
      13'hF4B: filaimg <= 9'b101110110;
      13'hF4C: filaimg <= 9'b101110110;
      13'hF4D: filaimg <= 9'b101110110;
      13'hF4E: filaimg <= 9'b101110110;
      13'hF4F: filaimg <= 9'b101110110;
      13'hF50: filaimg <= 9'b101110110;
      13'hF51: filaimg <= 9'b101110110;
      13'hF52: filaimg <= 9'b101110110;
      13'hF53: filaimg <= 9'b101110110;
      13'hF54: filaimg <= 9'b101110110;
      13'hF55: filaimg <= 9'b101110110;
      13'hF56: filaimg <= 9'b101110110;
      13'hF57: filaimg <= 9'b101110110;
      13'hF58: filaimg <= 9'b101110110;
      13'hF59: filaimg <= 9'b101110110;
      13'hF5A: filaimg <= 9'b101110110;
      13'hF5B: filaimg <= 9'b101110110;
      13'hF5C: filaimg <= 9'b101110110;
      13'hF5D: filaimg <= 9'b101110110;
      13'hF5E: filaimg <= 9'b101110110;
      13'hF5F: filaimg <= 9'b101110110;
      13'hF60: filaimg <= 9'b101110110;
      13'hF61: filaimg <= 9'b101110110;
      13'hF62: filaimg <= 9'b101110110;
      13'hF63: filaimg <= 9'b101110110;
      13'hF64: filaimg <= 9'b101110110;
      13'hF65: filaimg <= 9'b101110110;
      13'hF66: filaimg <= 9'b101110110;
      13'hF67: filaimg <= 9'b101110110;
      13'hF68: filaimg <= 9'b101110110;
      13'hF69: filaimg <= 9'b101110110;
      13'hF6A: filaimg <= 9'b101110110;
      13'hF6B: filaimg <= 9'b101110110;
      13'hF6C: filaimg <= 9'b101110110;
      13'hF6D: filaimg <= 9'b101110110;
      13'hF6E: filaimg <= 9'b101110110;
      13'hF6F: filaimg <= 9'b101110110;
      13'hF70: filaimg <= 9'b101110110;
      13'hF71: filaimg <= 9'b101110110;
      13'hF72: filaimg <= 9'b101110110;
      13'hF73: filaimg <= 9'b101110110;
      13'hF74: filaimg <= 9'b101110110;
      13'hF75: filaimg <= 9'b101110110;
      13'hF76: filaimg <= 9'b101110110;
      13'hF77: filaimg <= 9'b101110110;
      13'hF78: filaimg <= 9'b101110110;
      13'hF79: filaimg <= 9'b101110110;
      13'hF7A: filaimg <= 9'b101110110;
      13'hF7B: filaimg <= 9'b101110110;
      13'hF7C: filaimg <= 9'b101110110;
      13'hF7D: filaimg <= 9'b101110110;
      13'hF7E: filaimg <= 9'b101110110;
      13'hF7F: filaimg <= 9'b101110110;
      13'hF80: filaimg <= 9'b101110110;
      13'hF81: filaimg <= 9'b101110110;
      13'hF82: filaimg <= 9'b101110110;
      13'hF83: filaimg <= 9'b101110110;
      13'hF84: filaimg <= 9'b101110110;
      13'hF85: filaimg <= 9'b101110110;
      13'hF86: filaimg <= 9'b101110110;
      13'hF87: filaimg <= 9'b101110110;
      13'hF88: filaimg <= 9'b101110110;
      13'hF89: filaimg <= 9'b101110110;
      13'hF8A: filaimg <= 9'b101110110;
      13'hF8B: filaimg <= 9'b101110110;
      13'hF8C: filaimg <= 9'b101110110;
      13'hF8D: filaimg <= 9'b101110110;
      13'hF8E: filaimg <= 9'b101110110;
      13'hF8F: filaimg <= 9'b101110110;
      13'hF90: filaimg <= 9'b101110110;
      13'hF91: filaimg <= 9'b101110110;
      13'hF92: filaimg <= 9'b101110110;
      13'hF93: filaimg <= 9'b101110110;
      13'hF94: filaimg <= 9'b101110110;
      13'hF95: filaimg <= 9'b101110110;
      13'hF96: filaimg <= 9'b101110110;
      13'hF97: filaimg <= 9'b101110110;
      13'hF98: filaimg <= 9'b101110110;
      13'hF99: filaimg <= 9'b101110110;
      13'hF9A: filaimg <= 9'b101110110;
      13'hF9B: filaimg <= 9'b101110110;
      13'hF9C: filaimg <= 9'b101110110;
      13'hF9D: filaimg <= 9'b101110110;
      13'hF9E: filaimg <= 9'b101110110;
      13'hF9F: filaimg <= 9'b101110110;
      13'hFA0: filaimg <= 9'b101110110;
      13'hFA1: filaimg <= 9'b101110110;
      13'hFA2: filaimg <= 9'b101110110;
      13'hFA3: filaimg <= 9'b101110110;
      13'hFA4: filaimg <= 9'b101110110;
      13'hFA5: filaimg <= 9'b101110110;
      13'hFA6: filaimg <= 9'b101110110;
      13'hFA7: filaimg <= 9'b101110110;
      13'hFA8: filaimg <= 9'b101110110;
      13'hFA9: filaimg <= 9'b101110110;
      13'hFAA: filaimg <= 9'b101110110;
      13'hFAB: filaimg <= 9'b101110110;
      13'hFAC: filaimg <= 9'b101110110;
      13'hFAD: filaimg <= 9'b101110110;
      13'hFAE: filaimg <= 9'b101110110;
      13'hFAF: filaimg <= 9'b101110110;
      13'hFB0: filaimg <= 9'b101110110;
      13'hFB1: filaimg <= 9'b101110110;
      13'hFB2: filaimg <= 9'b101110110;
      13'hFB3: filaimg <= 9'b101110110;
      13'hFB4: filaimg <= 9'b101110110;
      13'hFB5: filaimg <= 9'b101110110;
      13'hFB6: filaimg <= 9'b101110110;
      13'hFB7: filaimg <= 9'b101110110;
      13'hFB8: filaimg <= 9'b101110110;
      13'hFB9: filaimg <= 9'b101110110;
      13'hFBA: filaimg <= 9'b101110110;
      13'hFBB: filaimg <= 9'b101110110;
      13'hFBC: filaimg <= 9'b101110110;
      13'hFBD: filaimg <= 9'b101110110;
      13'hFBE: filaimg <= 9'b101110110;
      13'hFBF: filaimg <= 9'b101110110;
      13'hFC0: filaimg <= 9'b101110110;
      13'hFC1: filaimg <= 9'b101110110;
      13'hFC2: filaimg <= 9'b101110110;
      13'hFC3: filaimg <= 9'b101110110;
      13'hFC4: filaimg <= 9'b101110110;
      13'hFC5: filaimg <= 9'b101110110;
      13'hFC6: filaimg <= 9'b101110110;
      13'hFC7: filaimg <= 9'b101110110;
      13'hFC8: filaimg <= 9'b101110110;
      13'hFC9: filaimg <= 9'b101110110;
      13'hFCA: filaimg <= 9'b101110110;
      13'hFCB: filaimg <= 9'b101110110;
      13'hFCC: filaimg <= 9'b101110110;
      13'hFCD: filaimg <= 9'b101110110;
      13'hFCE: filaimg <= 9'b101110110;
      13'hFCF: filaimg <= 9'b101110110;
      13'hFD0: filaimg <= 9'b101110110;
      13'hFD1: filaimg <= 9'b101110110;
      13'hFD2: filaimg <= 9'b101110110;
      13'hFD3: filaimg <= 9'b101110110;
      13'hFD4: filaimg <= 9'b101110110;
      13'hFD5: filaimg <= 9'b101110110;
      13'hFD6: filaimg <= 9'b101110110;
      13'hFD7: filaimg <= 9'b101110110;
      13'hFD8: filaimg <= 9'b101110110;
      13'hFD9: filaimg <= 9'b101110110;
      13'hFDA: filaimg <= 9'b101110110;
      13'hFDB: filaimg <= 9'b101110110;
      13'hFDC: filaimg <= 9'b101110110;
      13'hFDD: filaimg <= 9'b101110110;
      13'hFDE: filaimg <= 9'b101110110;
      13'hFDF: filaimg <= 9'b101110110;
      13'hFE0: filaimg <= 9'b101110110;
      13'hFE1: filaimg <= 9'b101110110;
      13'hFE2: filaimg <= 9'b101110110;
      13'hFE3: filaimg <= 9'b101110110;
      13'hFE4: filaimg <= 9'b101110110;
      13'hFE5: filaimg <= 9'b101110110;
      13'hFE6: filaimg <= 9'b101110110;
      13'hFE7: filaimg <= 9'b101110110;
      13'hFE8: filaimg <= 9'b101110110;
      13'hFE9: filaimg <= 9'b101110110;
      13'hFEA: filaimg <= 9'b101110110;
      13'hFEB: filaimg <= 9'b101110110;
      13'hFEC: filaimg <= 9'b101110110;
      13'hFED: filaimg <= 9'b101110110;
      13'hFEE: filaimg <= 9'b101110110;
      13'hFEF: filaimg <= 9'b101110110;
      13'hFF0: filaimg <= 9'b101110110;
      13'hFF1: filaimg <= 9'b101110110;
      13'hFF2: filaimg <= 9'b101110110;
      13'hFF3: filaimg <= 9'b101110110;
      13'hFF4: filaimg <= 9'b101110110;
      13'hFF5: filaimg <= 9'b101110110;
      13'hFF6: filaimg <= 9'b101110110;
      13'hFF7: filaimg <= 9'b101110110;
      13'hFF8: filaimg <= 9'b101110110;
      13'hFF9: filaimg <= 9'b101110110;
      13'hFFA: filaimg <= 9'b101110110;
      13'hFFB: filaimg <= 9'b101110110;
      13'hFFC: filaimg <= 9'b101110110;
      13'hFFD: filaimg <= 9'b101110110;
      13'hFFE: filaimg <= 9'b101110110;
      13'hFFF: filaimg <= 9'b101110110;
      13'h1000: filaimg <= 9'b101110110;
      13'h1001: filaimg <= 9'b101110110;
      13'h1002: filaimg <= 9'b101110110;
      13'h1003: filaimg <= 9'b101110110;
      13'h1004: filaimg <= 9'b101110110;
      13'h1005: filaimg <= 9'b101110110;
      13'h1006: filaimg <= 9'b101110110;
      13'h1007: filaimg <= 9'b101110110;
      13'h1008: filaimg <= 9'b101110110;
      13'h1009: filaimg <= 9'b101110110;
      13'h100A: filaimg <= 9'b101110110;
      13'h100B: filaimg <= 9'b101110110;
      13'h100C: filaimg <= 9'b101110110;
      13'h100D: filaimg <= 9'b101110110;
      13'h100E: filaimg <= 9'b101110110;
      13'h100F: filaimg <= 9'b101110110;
      13'h1010: filaimg <= 9'b101110110;
      13'h1011: filaimg <= 9'b101110110;
      13'h1012: filaimg <= 9'b101110110;
      13'h1013: filaimg <= 9'b101110110;
      13'h1014: filaimg <= 9'b101110110;
      13'h1015: filaimg <= 9'b101110110;
      13'h1016: filaimg <= 9'b101110110;
      13'h1017: filaimg <= 9'b101110110;
      13'h1018: filaimg <= 9'b101110110;
      13'h1019: filaimg <= 9'b101110110;
      13'h101A: filaimg <= 9'b101110110;
      13'h101B: filaimg <= 9'b101110110;
      13'h101C: filaimg <= 9'b101110110;
      13'h101D: filaimg <= 9'b101110110;
      13'h101E: filaimg <= 9'b101110110;
      13'h101F: filaimg <= 9'b101110110;
      13'h1020: filaimg <= 9'b101110110;
      13'h1021: filaimg <= 9'b101110110;
      13'h1022: filaimg <= 9'b101110110;
      13'h1023: filaimg <= 9'b101110110;
      13'h1024: filaimg <= 9'b101110110;
      13'h1025: filaimg <= 9'b101110110;
      13'h1026: filaimg <= 9'b101110110;
      13'h1027: filaimg <= 9'b101110110;
      13'h1028: filaimg <= 9'b101110110;
      13'h1029: filaimg <= 9'b101110110;
      13'h102A: filaimg <= 9'b101110110;
      13'h102B: filaimg <= 9'b101110110;
      13'h102C: filaimg <= 9'b101110110;
      13'h102D: filaimg <= 9'b101110110;
      13'h102E: filaimg <= 9'b101110110;
      13'h102F: filaimg <= 9'b101110110;
      13'h1030: filaimg <= 9'b101110110;
      13'h1031: filaimg <= 9'b101110110;
      13'h1032: filaimg <= 9'b101110110;
      13'h1033: filaimg <= 9'b101110110;
      13'h1034: filaimg <= 9'b101110110;
      13'h1035: filaimg <= 9'b101110110;
      13'h1036: filaimg <= 9'b101110110;
      13'h1037: filaimg <= 9'b101110110;
      13'h1038: filaimg <= 9'b101110110;
      13'h1039: filaimg <= 9'b101110110;
      13'h103A: filaimg <= 9'b101110110;
      13'h103B: filaimg <= 9'b101110110;
      13'h103C: filaimg <= 9'b101110110;
      13'h103D: filaimg <= 9'b101110110;
      13'h103E: filaimg <= 9'b101110110;
      13'h103F: filaimg <= 9'b101110110;
      13'h1040: filaimg <= 9'b101110110;
      13'h1041: filaimg <= 9'b101110110;
      13'h1042: filaimg <= 9'b101110110;
      13'h1043: filaimg <= 9'b101110110;
      13'h1044: filaimg <= 9'b101110110;
      13'h1045: filaimg <= 9'b101110110;
      13'h1046: filaimg <= 9'b101110110;
      13'h1047: filaimg <= 9'b101110110;
      13'h1048: filaimg <= 9'b101110110;
      13'h1049: filaimg <= 9'b101110110;
      13'h104A: filaimg <= 9'b101110110;
      13'h104B: filaimg <= 9'b101110110;
      13'h104C: filaimg <= 9'b101110110;
      13'h104D: filaimg <= 9'b101110110;
      13'h104E: filaimg <= 9'b101110110;
      13'h104F: filaimg <= 9'b101110110;
      13'h1050: filaimg <= 9'b101110110;
      13'h1051: filaimg <= 9'b101110110;
      13'h1052: filaimg <= 9'b101110110;
      13'h1053: filaimg <= 9'b101110110;
      13'h1054: filaimg <= 9'b101110110;
      13'h1055: filaimg <= 9'b101110110;
      13'h1056: filaimg <= 9'b101110110;
      13'h1057: filaimg <= 9'b101110110;
      13'h1058: filaimg <= 9'b101110110;
      13'h1059: filaimg <= 9'b101110110;
      13'h105A: filaimg <= 9'b101110110;
      13'h105B: filaimg <= 9'b101110110;
      13'h105C: filaimg <= 9'b101110110;
      13'h105D: filaimg <= 9'b101110110;
      13'h105E: filaimg <= 9'b101110110;
      13'h105F: filaimg <= 9'b101110110;
      13'h1060: filaimg <= 9'b101110110;
      13'h1061: filaimg <= 9'b101110110;
      13'h1062: filaimg <= 9'b101110110;
      13'h1063: filaimg <= 9'b101110110;
      13'h1064: filaimg <= 9'b101110110;
      13'h1065: filaimg <= 9'b101110110;
      13'h1066: filaimg <= 9'b101110110;
      13'h1067: filaimg <= 9'b101110110;
      13'h1068: filaimg <= 9'b101110110;
      13'h1069: filaimg <= 9'b101110110;
      13'h106A: filaimg <= 9'b101110110;
      13'h106B: filaimg <= 9'b101110110;
      13'h106C: filaimg <= 9'b101110110;
      13'h106D: filaimg <= 9'b101110110;
      13'h106E: filaimg <= 9'b101110110;
      13'h106F: filaimg <= 9'b101110110;
      13'h1070: filaimg <= 9'b101110110;
      13'h1071: filaimg <= 9'b101110110;
      13'h1072: filaimg <= 9'b101110110;
      13'h1073: filaimg <= 9'b101110110;
      13'h1074: filaimg <= 9'b101110110;
      13'h1075: filaimg <= 9'b101110110;
      13'h1076: filaimg <= 9'b101110110;
      13'h1077: filaimg <= 9'b101110110;
      13'h1078: filaimg <= 9'b101110110;
      13'h1079: filaimg <= 9'b101110110;
      13'h107A: filaimg <= 9'b101110110;
      13'h107B: filaimg <= 9'b101110110;
      13'h107C: filaimg <= 9'b101110110;
      13'h107D: filaimg <= 9'b101110110;
      13'h107E: filaimg <= 9'b101110110;
      13'h107F: filaimg <= 9'b101110110;
      13'h1080: filaimg <= 9'b101110110;
      13'h1081: filaimg <= 9'b101110110;
      13'h1082: filaimg <= 9'b101110110;
      13'h1083: filaimg <= 9'b101110110;
      13'h1084: filaimg <= 9'b101110110;
      13'h1085: filaimg <= 9'b101110110;
      13'h1086: filaimg <= 9'b101110110;
      13'h1087: filaimg <= 9'b101110110;
      13'h1088: filaimg <= 9'b101110110;
      13'h1089: filaimg <= 9'b101110110;
      13'h108A: filaimg <= 9'b101110110;
      13'h108B: filaimg <= 9'b101110110;
      13'h108C: filaimg <= 9'b101110110;
      13'h108D: filaimg <= 9'b101110110;
      13'h108E: filaimg <= 9'b101110110;
      13'h108F: filaimg <= 9'b101110110;
      13'h1090: filaimg <= 9'b101110110;
      13'h1091: filaimg <= 9'b101110110;
      13'h1092: filaimg <= 9'b101110110;
      13'h1093: filaimg <= 9'b101110110;
      13'h1094: filaimg <= 9'b101110110;
      13'h1095: filaimg <= 9'b101110110;
      13'h1096: filaimg <= 9'b101110110;
      13'h1097: filaimg <= 9'b101110110;
      13'h1098: filaimg <= 9'b101110110;
      13'h1099: filaimg <= 9'b101110110;
      13'h109A: filaimg <= 9'b101110110;
      13'h109B: filaimg <= 9'b101110110;
      13'h109C: filaimg <= 9'b101110110;
      13'h109D: filaimg <= 9'b101110110;
      13'h109E: filaimg <= 9'b101110110;
      13'h109F: filaimg <= 9'b101110110;
      13'h10A0: filaimg <= 9'b101110110;
      13'h10A1: filaimg <= 9'b101110110;
      13'h10A2: filaimg <= 9'b101110110;
      13'h10A3: filaimg <= 9'b101110110;
      13'h10A4: filaimg <= 9'b101110110;
      13'h10A5: filaimg <= 9'b101110110;
      13'h10A6: filaimg <= 9'b101110110;
      13'h10A7: filaimg <= 9'b101110110;
      13'h10A8: filaimg <= 9'b101110110;
      13'h10A9: filaimg <= 9'b101110110;
      13'h10AA: filaimg <= 9'b101110110;
      13'h10AB: filaimg <= 9'b101110110;
      13'h10AC: filaimg <= 9'b101110110;
      13'h10AD: filaimg <= 9'b101110110;
      13'h10AE: filaimg <= 9'b101110110;
      13'h10AF: filaimg <= 9'b101110110;
      13'h10B0: filaimg <= 9'b101110110;
      13'h10B1: filaimg <= 9'b101110110;
      13'h10B2: filaimg <= 9'b101110110;
      13'h10B3: filaimg <= 9'b101110110;
      13'h10B4: filaimg <= 9'b101110110;
      13'h10B5: filaimg <= 9'b101110110;
      13'h10B6: filaimg <= 9'b101110110;
      13'h10B7: filaimg <= 9'b101110110;
      13'h10B8: filaimg <= 9'b101110110;
      13'h10B9: filaimg <= 9'b101110110;
      13'h10BA: filaimg <= 9'b101110110;
      13'h10BB: filaimg <= 9'b101110110;
      13'h10BC: filaimg <= 9'b101110110;
      13'h10BD: filaimg <= 9'b101110110;
      13'h10BE: filaimg <= 9'b101110110;
      13'h10BF: filaimg <= 9'b101110110;
      13'h10C0: filaimg <= 9'b101110110;
      13'h10C1: filaimg <= 9'b101110110;
      13'h10C2: filaimg <= 9'b101110110;
      13'h10C3: filaimg <= 9'b101110110;
      13'h10C4: filaimg <= 9'b101110110;
      13'h10C5: filaimg <= 9'b101110110;
      13'h10C6: filaimg <= 9'b101110110;
      13'h10C7: filaimg <= 9'b101110110;
      13'h10C8: filaimg <= 9'b101110110;
      13'h10C9: filaimg <= 9'b101110110;
      13'h10CA: filaimg <= 9'b101110110;
      13'h10CB: filaimg <= 9'b101110110;
      13'h10CC: filaimg <= 9'b101110110;
      13'h10CD: filaimg <= 9'b101110110;
      13'h10CE: filaimg <= 9'b101110110;
      13'h10CF: filaimg <= 9'b101110110;
      13'h10D0: filaimg <= 9'b101110110;
      13'h10D1: filaimg <= 9'b101110110;
      13'h10D2: filaimg <= 9'b101110110;
      13'h10D3: filaimg <= 9'b101110110;
      13'h10D4: filaimg <= 9'b101110110;
      13'h10D5: filaimg <= 9'b101110110;
      13'h10D6: filaimg <= 9'b101110110;
      13'h10D7: filaimg <= 9'b101110110;
      13'h10D8: filaimg <= 9'b101110110;
      13'h10D9: filaimg <= 9'b101110110;
      13'h10DA: filaimg <= 9'b101110110;
      13'h10DB: filaimg <= 9'b101110110;
      13'h10DC: filaimg <= 9'b101110110;
      13'h10DD: filaimg <= 9'b101110110;
      13'h10DE: filaimg <= 9'b101110110;
      13'h10DF: filaimg <= 9'b101110110;
      13'h10E0: filaimg <= 9'b101110110;
      13'h10E1: filaimg <= 9'b101110110;
      13'h10E2: filaimg <= 9'b101110110;
      13'h10E3: filaimg <= 9'b101110110;
      13'h10E4: filaimg <= 9'b101110110;
      13'h10E5: filaimg <= 9'b101110110;
      13'h10E6: filaimg <= 9'b101110110;
      13'h10E7: filaimg <= 9'b101110110;
      13'h10E8: filaimg <= 9'b101110110;
      13'h10E9: filaimg <= 9'b101110110;
      13'h10EA: filaimg <= 9'b101110110;
      13'h10EB: filaimg <= 9'b101110110;
      13'h10EC: filaimg <= 9'b101110110;
      13'h10ED: filaimg <= 9'b101110110;
      13'h10EE: filaimg <= 9'b101110110;
      13'h10EF: filaimg <= 9'b101110110;
      13'h10F0: filaimg <= 9'b101110110;
      13'h10F1: filaimg <= 9'b101110110;
      13'h10F2: filaimg <= 9'b101110110;
      13'h10F3: filaimg <= 9'b101110110;
      13'h10F4: filaimg <= 9'b101110110;
      13'h10F5: filaimg <= 9'b101110110;
      13'h10F6: filaimg <= 9'b101110110;
      13'h10F7: filaimg <= 9'b101110110;
      13'h10F8: filaimg <= 9'b101110110;
      13'h10F9: filaimg <= 9'b101110110;
      13'h10FA: filaimg <= 9'b101110110;
      13'h10FB: filaimg <= 9'b101110110;
      13'h10FC: filaimg <= 9'b101110110;
      13'h10FD: filaimg <= 9'b101110110;
      13'h10FE: filaimg <= 9'b101110110;
      13'h10FF: filaimg <= 9'b101110110;
      13'h1100: filaimg <= 9'b101110110;
      13'h1101: filaimg <= 9'b101110110;
      13'h1102: filaimg <= 9'b101110110;
      13'h1103: filaimg <= 9'b101110110;
      13'h1104: filaimg <= 9'b101110110;
      13'h1105: filaimg <= 9'b101110110;
      13'h1106: filaimg <= 9'b101110110;
      13'h1107: filaimg <= 9'b101110110;
      13'h1108: filaimg <= 9'b101110110;
      13'h1109: filaimg <= 9'b101110110;
      13'h110A: filaimg <= 9'b101110110;
      13'h110B: filaimg <= 9'b101110110;
      13'h110C: filaimg <= 9'b101110110;
      13'h110D: filaimg <= 9'b101110110;
      13'h110E: filaimg <= 9'b101110110;
      13'h110F: filaimg <= 9'b101110110;
      13'h1110: filaimg <= 9'b101110110;
      13'h1111: filaimg <= 9'b101110110;
      13'h1112: filaimg <= 9'b101110110;
      13'h1113: filaimg <= 9'b101110110;
      13'h1114: filaimg <= 9'b101110110;
      13'h1115: filaimg <= 9'b101110110;
      13'h1116: filaimg <= 9'b101110110;
      13'h1117: filaimg <= 9'b101110110;
      13'h1118: filaimg <= 9'b101110110;
      13'h1119: filaimg <= 9'b101110110;
      13'h111A: filaimg <= 9'b101110110;
      13'h111B: filaimg <= 9'b101110110;
      13'h111C: filaimg <= 9'b101110110;
      13'h111D: filaimg <= 9'b101110110;
      13'h111E: filaimg <= 9'b101110110;
      13'h111F: filaimg <= 9'b101110110;
      13'h1120: filaimg <= 9'b101110110;
      13'h1121: filaimg <= 9'b101110110;
      13'h1122: filaimg <= 9'b101110110;
      13'h1123: filaimg <= 9'b101110110;
      13'h1124: filaimg <= 9'b101110110;
      13'h1125: filaimg <= 9'b101110110;
      13'h1126: filaimg <= 9'b101110110;
      13'h1127: filaimg <= 9'b101110110;
      13'h1128: filaimg <= 9'b101110110;
      13'h1129: filaimg <= 9'b101110110;
      13'h112A: filaimg <= 9'b101110110;
      13'h112B: filaimg <= 9'b101110110;
      13'h112C: filaimg <= 9'b101110110;
      13'h112D: filaimg <= 9'b101110110;
      13'h112E: filaimg <= 9'b101110110;
      13'h112F: filaimg <= 9'b101110110;
      13'h1130: filaimg <= 9'b101110110;
      13'h1131: filaimg <= 9'b101110110;
      13'h1132: filaimg <= 9'b101110110;
      13'h1133: filaimg <= 9'b101110110;
      13'h1134: filaimg <= 9'b101110110;
      13'h1135: filaimg <= 9'b101110110;
      13'h1136: filaimg <= 9'b101110110;
      13'h1137: filaimg <= 9'b101110110;
      13'h1138: filaimg <= 9'b101110110;
      13'h1139: filaimg <= 9'b101110110;
      13'h113A: filaimg <= 9'b101110110;
      13'h113B: filaimg <= 9'b101110110;
      13'h113C: filaimg <= 9'b101110110;
      13'h113D: filaimg <= 9'b101110110;
      13'h113E: filaimg <= 9'b101110110;
      13'h113F: filaimg <= 9'b101110110;
      13'h1140: filaimg <= 9'b101110110;
      13'h1141: filaimg <= 9'b101110110;
      13'h1142: filaimg <= 9'b101110110;
      13'h1143: filaimg <= 9'b101110110;
      13'h1144: filaimg <= 9'b101110110;
      13'h1145: filaimg <= 9'b101110110;
      13'h1146: filaimg <= 9'b101110110;
      13'h1147: filaimg <= 9'b101110110;
      13'h1148: filaimg <= 9'b101110110;
      13'h1149: filaimg <= 9'b101110110;
      13'h114A: filaimg <= 9'b101110110;
      13'h114B: filaimg <= 9'b101110110;
      13'h114C: filaimg <= 9'b101110110;
      13'h114D: filaimg <= 9'b101110110;
      13'h114E: filaimg <= 9'b101110110;
      13'h114F: filaimg <= 9'b101110110;
      13'h1150: filaimg <= 9'b101110110;
      13'h1151: filaimg <= 9'b101110110;
      13'h1152: filaimg <= 9'b101110110;
      13'h1153: filaimg <= 9'b101110110;
      13'h1154: filaimg <= 9'b101110110;
      13'h1155: filaimg <= 9'b101110110;
      13'h1156: filaimg <= 9'b101110110;
      13'h1157: filaimg <= 9'b101110110;
      13'h1158: filaimg <= 9'b101110110;
      13'h1159: filaimg <= 9'b101110110;
      13'h115A: filaimg <= 9'b101110110;
      13'h115B: filaimg <= 9'b101110110;
      13'h115C: filaimg <= 9'b101110110;
      13'h115D: filaimg <= 9'b101110110;
      13'h115E: filaimg <= 9'b101110110;
      13'h115F: filaimg <= 9'b101110110;
      13'h1160: filaimg <= 9'b101110110;
      13'h1161: filaimg <= 9'b101110110;
      13'h1162: filaimg <= 9'b101110110;
      13'h1163: filaimg <= 9'b101110110;
      13'h1164: filaimg <= 9'b101110110;
      13'h1165: filaimg <= 9'b101110110;
      13'h1166: filaimg <= 9'b101110110;
      13'h1167: filaimg <= 9'b101110110;
      13'h1168: filaimg <= 9'b101110110;
      13'h1169: filaimg <= 9'b101110110;
      13'h116A: filaimg <= 9'b101110110;
      13'h116B: filaimg <= 9'b101110110;
      13'h116C: filaimg <= 9'b101110110;
      13'h116D: filaimg <= 9'b101110110;
      13'h116E: filaimg <= 9'b101110110;
      13'h116F: filaimg <= 9'b101110110;
      13'h1170: filaimg <= 9'b101110110;
      13'h1171: filaimg <= 9'b101110110;
      13'h1172: filaimg <= 9'b101110110;
      13'h1173: filaimg <= 9'b101110110;
      13'h1174: filaimg <= 9'b101110110;
      13'h1175: filaimg <= 9'b101110110;
      13'h1176: filaimg <= 9'b101110110;
      13'h1177: filaimg <= 9'b101110110;
      13'h1178: filaimg <= 9'b101110110;
      13'h1179: filaimg <= 9'b101110110;
      13'h117A: filaimg <= 9'b101110110;
      13'h117B: filaimg <= 9'b101110110;
      13'h117C: filaimg <= 9'b101110110;
      13'h117D: filaimg <= 9'b101110110;
      13'h117E: filaimg <= 9'b101110110;
      13'h117F: filaimg <= 9'b101110110;
      13'h1180: filaimg <= 9'b101110110;
      13'h1181: filaimg <= 9'b101110110;
      13'h1182: filaimg <= 9'b101110110;
      13'h1183: filaimg <= 9'b101110110;
      13'h1184: filaimg <= 9'b101110110;
      13'h1185: filaimg <= 9'b101110110;
      13'h1186: filaimg <= 9'b101110110;
      13'h1187: filaimg <= 9'b101110110;
      13'h1188: filaimg <= 9'b101110110;
      13'h1189: filaimg <= 9'b101110110;
      13'h118A: filaimg <= 9'b101110110;
      13'h118B: filaimg <= 9'b101110110;
      13'h118C: filaimg <= 9'b101110110;
      13'h118D: filaimg <= 9'b101110110;
      13'h118E: filaimg <= 9'b101110110;
      13'h118F: filaimg <= 9'b101110110;
      13'h1190: filaimg <= 9'b101110110;
      13'h1191: filaimg <= 9'b101110110;
      13'h1192: filaimg <= 9'b101110110;
      13'h1193: filaimg <= 9'b101110110;
      13'h1194: filaimg <= 9'b101110110;
      13'h1195: filaimg <= 9'b101110110;
      13'h1196: filaimg <= 9'b101110110;
      13'h1197: filaimg <= 9'b101110110;
      13'h1198: filaimg <= 9'b101110110;
      13'h1199: filaimg <= 9'b101110110;
      13'h119A: filaimg <= 9'b101110110;
      13'h119B: filaimg <= 9'b101110110;
      13'h119C: filaimg <= 9'b101110110;
      13'h119D: filaimg <= 9'b101110110;
      13'h119E: filaimg <= 9'b101110110;
      13'h119F: filaimg <= 9'b101110110;
      13'h11A0: filaimg <= 9'b101110110;
      13'h11A1: filaimg <= 9'b101110110;
      13'h11A2: filaimg <= 9'b101110110;
      13'h11A3: filaimg <= 9'b101110110;
      13'h11A4: filaimg <= 9'b101110110;
      13'h11A5: filaimg <= 9'b101110110;
      13'h11A6: filaimg <= 9'b101110110;
      13'h11A7: filaimg <= 9'b101110110;
      13'h11A8: filaimg <= 9'b101110110;
      13'h11A9: filaimg <= 9'b101110110;
      13'h11AA: filaimg <= 9'b101110110;
      13'h11AB: filaimg <= 9'b101110110;
      13'h11AC: filaimg <= 9'b101110110;
      13'h11AD: filaimg <= 9'b101110110;
      13'h11AE: filaimg <= 9'b101110110;
      13'h11AF: filaimg <= 9'b101110110;
      13'h11B0: filaimg <= 9'b101110110;
      13'h11B1: filaimg <= 9'b101110110;
      13'h11B2: filaimg <= 9'b101110110;
      13'h11B3: filaimg <= 9'b101110110;
      13'h11B4: filaimg <= 9'b101110110;
      13'h11B5: filaimg <= 9'b101110110;
      13'h11B6: filaimg <= 9'b101110110;
      13'h11B7: filaimg <= 9'b101110110;
      13'h11B8: filaimg <= 9'b101110110;
      13'h11B9: filaimg <= 9'b101110110;
      13'h11BA: filaimg <= 9'b101110110;
      13'h11BB: filaimg <= 9'b101110110;
      13'h11BC: filaimg <= 9'b101110110;
      13'h11BD: filaimg <= 9'b101110110;
      13'h11BE: filaimg <= 9'b101110110;
      13'h11BF: filaimg <= 9'b101110110;
      13'h11C0: filaimg <= 9'b101110110;
      13'h11C1: filaimg <= 9'b101110110;
      13'h11C2: filaimg <= 9'b101110110;
      13'h11C3: filaimg <= 9'b101110110;
      13'h11C4: filaimg <= 9'b101110110;
      13'h11C5: filaimg <= 9'b101110110;
      13'h11C6: filaimg <= 9'b101110110;
      13'h11C7: filaimg <= 9'b101110110;
      13'h11C8: filaimg <= 9'b101110110;
      13'h11C9: filaimg <= 9'b101110110;
      13'h11CA: filaimg <= 9'b101110110;
      13'h11CB: filaimg <= 9'b101110110;
      13'h11CC: filaimg <= 9'b101110110;
      13'h11CD: filaimg <= 9'b101110110;
      13'h11CE: filaimg <= 9'b101110110;
      13'h11CF: filaimg <= 9'b101110110;
      13'h11D0: filaimg <= 9'b101110110;
      13'h11D1: filaimg <= 9'b101110110;
      13'h11D2: filaimg <= 9'b101110110;
      13'h11D3: filaimg <= 9'b101110110;
      13'h11D4: filaimg <= 9'b101110110;
      13'h11D5: filaimg <= 9'b101110110;
      13'h11D6: filaimg <= 9'b101110110;
      13'h11D7: filaimg <= 9'b101110110;
      13'h11D8: filaimg <= 9'b101110110;
      13'h11D9: filaimg <= 9'b101110110;
      13'h11DA: filaimg <= 9'b101110110;
      13'h11DB: filaimg <= 9'b101110110;
      13'h11DC: filaimg <= 9'b101110110;
      13'h11DD: filaimg <= 9'b101110110;
      13'h11DE: filaimg <= 9'b101110110;
      13'h11DF: filaimg <= 9'b101110110;
      13'h11E0: filaimg <= 9'b101110110;
      13'h11E1: filaimg <= 9'b101110110;
      13'h11E2: filaimg <= 9'b101110110;
      13'h11E3: filaimg <= 9'b101110110;
      13'h11E4: filaimg <= 9'b101110110;
      13'h11E5: filaimg <= 9'b101110110;
      13'h11E6: filaimg <= 9'b101110110;
      13'h11E7: filaimg <= 9'b101110110;
      13'h11E8: filaimg <= 9'b101110110;
      13'h11E9: filaimg <= 9'b101110110;
      13'h11EA: filaimg <= 9'b101110110;
      13'h11EB: filaimg <= 9'b101110110;
      13'h11EC: filaimg <= 9'b101110110;
      13'h11ED: filaimg <= 9'b101110110;
      13'h11EE: filaimg <= 9'b101110110;
      13'h11EF: filaimg <= 9'b101110110;
      13'h11F0: filaimg <= 9'b101110110;
      13'h11F1: filaimg <= 9'b101110110;
      13'h11F2: filaimg <= 9'b101110110;
      13'h11F3: filaimg <= 9'b101110110;
      13'h11F4: filaimg <= 9'b101110110;
      13'h11F5: filaimg <= 9'b101110110;
      13'h11F6: filaimg <= 9'b101110110;
      13'h11F7: filaimg <= 9'b101110110;
      13'h11F8: filaimg <= 9'b101110110;
      13'h11F9: filaimg <= 9'b101110110;
      13'h11FA: filaimg <= 9'b101110110;
      13'h11FB: filaimg <= 9'b101110110;
      13'h11FC: filaimg <= 9'b101110110;
      13'h11FD: filaimg <= 9'b101110110;
      13'h11FE: filaimg <= 9'b101110110;
      13'h11FF: filaimg <= 9'b101110110;
      13'h1200: filaimg <= 9'b101110110;
      13'h1201: filaimg <= 9'b101110110;
      13'h1202: filaimg <= 9'b101110110;
      13'h1203: filaimg <= 9'b101110110;
      13'h1204: filaimg <= 9'b101110110;
      13'h1205: filaimg <= 9'b101110110;
      13'h1206: filaimg <= 9'b101110110;
      13'h1207: filaimg <= 9'b101110110;
      13'h1208: filaimg <= 9'b101110110;
      13'h1209: filaimg <= 9'b101110110;
      13'h120A: filaimg <= 9'b101110110;
      13'h120B: filaimg <= 9'b101110110;
      13'h120C: filaimg <= 9'b101110110;
      13'h120D: filaimg <= 9'b101110110;
      13'h120E: filaimg <= 9'b101110110;
      13'h120F: filaimg <= 9'b101110110;
      13'h1210: filaimg <= 9'b101110110;
      13'h1211: filaimg <= 9'b101110110;
      13'h1212: filaimg <= 9'b101110110;
      13'h1213: filaimg <= 9'b101110110;
      13'h1214: filaimg <= 9'b101110110;
      13'h1215: filaimg <= 9'b101110110;
      13'h1216: filaimg <= 9'b101110110;
      13'h1217: filaimg <= 9'b101110110;
      13'h1218: filaimg <= 9'b101110110;
      13'h1219: filaimg <= 9'b101110110;
      13'h121A: filaimg <= 9'b101110110;
      13'h121B: filaimg <= 9'b101110110;
      13'h121C: filaimg <= 9'b101110110;
      13'h121D: filaimg <= 9'b101110110;
      13'h121E: filaimg <= 9'b101110110;
      13'h121F: filaimg <= 9'b101110110;
      13'h1220: filaimg <= 9'b101110110;
      13'h1221: filaimg <= 9'b101110110;
      13'h1222: filaimg <= 9'b101110110;
      13'h1223: filaimg <= 9'b101110110;
      13'h1224: filaimg <= 9'b101110110;
      13'h1225: filaimg <= 9'b101110110;
      13'h1226: filaimg <= 9'b101110110;
      13'h1227: filaimg <= 9'b101110110;
      13'h1228: filaimg <= 9'b101110110;
      13'h1229: filaimg <= 9'b101110110;
      13'h122A: filaimg <= 9'b101110110;
      13'h122B: filaimg <= 9'b101110110;
      13'h122C: filaimg <= 9'b101110110;
      13'h122D: filaimg <= 9'b101110110;
      13'h122E: filaimg <= 9'b101110110;
      13'h122F: filaimg <= 9'b101110110;
      13'h1230: filaimg <= 9'b101110110;
      13'h1231: filaimg <= 9'b101110110;
      13'h1232: filaimg <= 9'b101110110;
      13'h1233: filaimg <= 9'b101110110;
      13'h1234: filaimg <= 9'b101110110;
      13'h1235: filaimg <= 9'b101110110;
      13'h1236: filaimg <= 9'b101110110;
      13'h1237: filaimg <= 9'b101110110;
      13'h1238: filaimg <= 9'b101110110;
      13'h1239: filaimg <= 9'b101110110;
      13'h123A: filaimg <= 9'b101110110;
      13'h123B: filaimg <= 9'b101110110;
      13'h123C: filaimg <= 9'b101110110;
      13'h123D: filaimg <= 9'b101110110;
      13'h123E: filaimg <= 9'b101110110;
      13'h123F: filaimg <= 9'b101110110;
      13'h1240: filaimg <= 9'b101110110;
      13'h1241: filaimg <= 9'b101110110;
      13'h1242: filaimg <= 9'b101110110;
      13'h1243: filaimg <= 9'b101110110;
      13'h1244: filaimg <= 9'b101110110;
      13'h1245: filaimg <= 9'b101110110;
      13'h1246: filaimg <= 9'b101110110;
      13'h1247: filaimg <= 9'b101110110;
      13'h1248: filaimg <= 9'b101110110;
      13'h1249: filaimg <= 9'b101110110;
      13'h124A: filaimg <= 9'b101110110;
      13'h124B: filaimg <= 9'b101110110;
      13'h124C: filaimg <= 9'b101110110;
      13'h124D: filaimg <= 9'b101110110;
      13'h124E: filaimg <= 9'b101110110;
      13'h124F: filaimg <= 9'b101110110;
      13'h1250: filaimg <= 9'b101110110;
      13'h1251: filaimg <= 9'b101110110;
      13'h1252: filaimg <= 9'b101110110;
      13'h1253: filaimg <= 9'b101110110;
      13'h1254: filaimg <= 9'b101110110;
      13'h1255: filaimg <= 9'b101110110;
      13'h1256: filaimg <= 9'b101110110;
      13'h1257: filaimg <= 9'b101110110;
      13'h1258: filaimg <= 9'b101110110;
      13'h1259: filaimg <= 9'b101110110;
      13'h125A: filaimg <= 9'b101110110;
      13'h125B: filaimg <= 9'b101110110;
      13'h125C: filaimg <= 9'b101110110;
      13'h125D: filaimg <= 9'b101110110;
      13'h125E: filaimg <= 9'b101110110;
      13'h125F: filaimg <= 9'b101110110;
      13'h1260: filaimg <= 9'b101110110;
      13'h1261: filaimg <= 9'b101110110;
      13'h1262: filaimg <= 9'b101110110;
      13'h1263: filaimg <= 9'b101110110;
      13'h1264: filaimg <= 9'b101110110;
      13'h1265: filaimg <= 9'b101110110;
      13'h1266: filaimg <= 9'b101110110;
      13'h1267: filaimg <= 9'b101110110;
      13'h1268: filaimg <= 9'b101110110;
      13'h1269: filaimg <= 9'b101110110;
      13'h126A: filaimg <= 9'b101110110;
      13'h126B: filaimg <= 9'b101110110;
      13'h126C: filaimg <= 9'b101110110;
      13'h126D: filaimg <= 9'b101110110;
      13'h126E: filaimg <= 9'b101110110;
      13'h126F: filaimg <= 9'b101110110;
      13'h1270: filaimg <= 9'b101110110;
      13'h1271: filaimg <= 9'b101110110;
      13'h1272: filaimg <= 9'b101110110;
      13'h1273: filaimg <= 9'b101110110;
      13'h1274: filaimg <= 9'b101110110;
      13'h1275: filaimg <= 9'b101110110;
      13'h1276: filaimg <= 9'b101110110;
      13'h1277: filaimg <= 9'b101110110;
      13'h1278: filaimg <= 9'b101110110;
      13'h1279: filaimg <= 9'b101110110;
      13'h127A: filaimg <= 9'b101110110;
      13'h127B: filaimg <= 9'b101110110;
      13'h127C: filaimg <= 9'b101110110;
      13'h127D: filaimg <= 9'b101110110;
      13'h127E: filaimg <= 9'b101110110;
      13'h127F: filaimg <= 9'b101110110;
      13'h1280: filaimg <= 9'b101110110;
      13'h1281: filaimg <= 9'b101110110;
      13'h1282: filaimg <= 9'b101110110;
      13'h1283: filaimg <= 9'b101110110;
      13'h1284: filaimg <= 9'b101110110;
      13'h1285: filaimg <= 9'b101110110;
      13'h1286: filaimg <= 9'b101110110;
      13'h1287: filaimg <= 9'b101110110;
      13'h1288: filaimg <= 9'b101110110;
      13'h1289: filaimg <= 9'b101110110;
      13'h128A: filaimg <= 9'b101110110;
      13'h128B: filaimg <= 9'b101110110;
      13'h128C: filaimg <= 9'b101110110;
      13'h128D: filaimg <= 9'b101110110;
      13'h128E: filaimg <= 9'b101110110;
      13'h128F: filaimg <= 9'b101110110;
      13'h1290: filaimg <= 9'b101110110;
      13'h1291: filaimg <= 9'b101110110;
      13'h1292: filaimg <= 9'b101110110;
      13'h1293: filaimg <= 9'b101110110;
      13'h1294: filaimg <= 9'b101110110;
      13'h1295: filaimg <= 9'b101110110;
      13'h1296: filaimg <= 9'b101110110;
      13'h1297: filaimg <= 9'b101110110;
      13'h1298: filaimg <= 9'b101110110;
      13'h1299: filaimg <= 9'b101110110;
      13'h129A: filaimg <= 9'b101110110;
      13'h129B: filaimg <= 9'b101110110;
      13'h129C: filaimg <= 9'b101110110;
      13'h129D: filaimg <= 9'b101110110;
      13'h129E: filaimg <= 9'b101110110;
      13'h129F: filaimg <= 9'b101110110;
      13'h12A0: filaimg <= 9'b101110110;
      13'h12A1: filaimg <= 9'b101110110;
      13'h12A2: filaimg <= 9'b101110110;
      13'h12A3: filaimg <= 9'b101110110;
      13'h12A4: filaimg <= 9'b101110110;
      13'h12A5: filaimg <= 9'b101110110;
      13'h12A6: filaimg <= 9'b101110110;
      13'h12A7: filaimg <= 9'b101110110;
      13'h12A8: filaimg <= 9'b101110110;
      13'h12A9: filaimg <= 9'b101110110;
      13'h12AA: filaimg <= 9'b101110110;
      13'h12AB: filaimg <= 9'b101110110;
      13'h12AC: filaimg <= 9'b101110110;
      13'h12AD: filaimg <= 9'b101110110;
      13'h12AE: filaimg <= 9'b101110110;
      13'h12AF: filaimg <= 9'b101110110;
      13'h12B0: filaimg <= 9'b101110110;
      13'h12B1: filaimg <= 9'b101110110;
      13'h12B2: filaimg <= 9'b101110110;
      13'h12B3: filaimg <= 9'b101110110;
      13'h12B4: filaimg <= 9'b101110110;
      13'h12B5: filaimg <= 9'b101110110;
      13'h12B6: filaimg <= 9'b101110110;
      13'h12B7: filaimg <= 9'b101110110;
      13'h12B8: filaimg <= 9'b101110110;
      13'h12B9: filaimg <= 9'b101110110;
      13'h12BA: filaimg <= 9'b101110110;
      13'h12BB: filaimg <= 9'b101110110;
      13'h12BC: filaimg <= 9'b101110110;
      13'h12BD: filaimg <= 9'b101110110;
      13'h12BE: filaimg <= 9'b101110110;
      13'h12BF: filaimg <= 9'b101110110;
      default: filaimg <= 9'b101110110;
    endcase
  end

endmodule
