// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jul 16 2019 20:09:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__84558;
    wire N__84544;
    wire N__84543;
    wire N__84542;
    wire N__84535;
    wire N__84534;
    wire N__84533;
    wire N__84526;
    wire N__84525;
    wire N__84524;
    wire N__84517;
    wire N__84516;
    wire N__84515;
    wire N__84508;
    wire N__84507;
    wire N__84506;
    wire N__84499;
    wire N__84498;
    wire N__84497;
    wire N__84490;
    wire N__84489;
    wire N__84488;
    wire N__84481;
    wire N__84480;
    wire N__84479;
    wire N__84472;
    wire N__84471;
    wire N__84470;
    wire N__84463;
    wire N__84462;
    wire N__84461;
    wire N__84444;
    wire N__84441;
    wire N__84438;
    wire N__84435;
    wire N__84434;
    wire N__84433;
    wire N__84426;
    wire N__84423;
    wire N__84420;
    wire N__84417;
    wire N__84414;
    wire N__84411;
    wire N__84408;
    wire N__84405;
    wire N__84402;
    wire N__84399;
    wire N__84396;
    wire N__84395;
    wire N__84394;
    wire N__84391;
    wire N__84386;
    wire N__84383;
    wire N__84380;
    wire N__84377;
    wire N__84374;
    wire N__84371;
    wire N__84368;
    wire N__84363;
    wire N__84360;
    wire N__84357;
    wire N__84354;
    wire N__84351;
    wire N__84350;
    wire N__84349;
    wire N__84346;
    wire N__84341;
    wire N__84338;
    wire N__84335;
    wire N__84332;
    wire N__84329;
    wire N__84326;
    wire N__84323;
    wire N__84318;
    wire N__84315;
    wire N__84312;
    wire N__84309;
    wire N__84306;
    wire N__84303;
    wire N__84302;
    wire N__84301;
    wire N__84300;
    wire N__84297;
    wire N__84296;
    wire N__84295;
    wire N__84294;
    wire N__84293;
    wire N__84292;
    wire N__84291;
    wire N__84290;
    wire N__84289;
    wire N__84288;
    wire N__84287;
    wire N__84284;
    wire N__84281;
    wire N__84272;
    wire N__84263;
    wire N__84260;
    wire N__84253;
    wire N__84250;
    wire N__84245;
    wire N__84240;
    wire N__84237;
    wire N__84234;
    wire N__84229;
    wire N__84226;
    wire N__84221;
    wire N__84218;
    wire N__84215;
    wire N__84212;
    wire N__84209;
    wire N__84204;
    wire N__84201;
    wire N__84198;
    wire N__84195;
    wire N__84194;
    wire N__84193;
    wire N__84186;
    wire N__84183;
    wire N__84180;
    wire N__84177;
    wire N__84174;
    wire N__84171;
    wire N__84168;
    wire N__84165;
    wire N__84162;
    wire N__84161;
    wire N__84160;
    wire N__84153;
    wire N__84150;
    wire N__84147;
    wire N__84144;
    wire N__84141;
    wire N__84138;
    wire N__84135;
    wire N__84134;
    wire N__84133;
    wire N__84126;
    wire N__84123;
    wire N__84120;
    wire N__84117;
    wire N__84114;
    wire N__84113;
    wire N__84112;
    wire N__84111;
    wire N__84110;
    wire N__84109;
    wire N__84108;
    wire N__84107;
    wire N__84106;
    wire N__84105;
    wire N__84104;
    wire N__84103;
    wire N__84102;
    wire N__84101;
    wire N__84100;
    wire N__84099;
    wire N__84098;
    wire N__84097;
    wire N__84096;
    wire N__84095;
    wire N__84094;
    wire N__84093;
    wire N__84092;
    wire N__84091;
    wire N__84090;
    wire N__84089;
    wire N__84088;
    wire N__84087;
    wire N__84086;
    wire N__84085;
    wire N__84084;
    wire N__84083;
    wire N__84082;
    wire N__84081;
    wire N__84080;
    wire N__84079;
    wire N__84078;
    wire N__84077;
    wire N__84076;
    wire N__84075;
    wire N__84074;
    wire N__84073;
    wire N__84072;
    wire N__84071;
    wire N__84070;
    wire N__84069;
    wire N__84068;
    wire N__84067;
    wire N__84066;
    wire N__84065;
    wire N__84064;
    wire N__84063;
    wire N__84062;
    wire N__84061;
    wire N__84060;
    wire N__84059;
    wire N__84058;
    wire N__84057;
    wire N__84056;
    wire N__84055;
    wire N__84054;
    wire N__84053;
    wire N__84052;
    wire N__84051;
    wire N__84050;
    wire N__84049;
    wire N__84048;
    wire N__84047;
    wire N__84046;
    wire N__84045;
    wire N__84044;
    wire N__84043;
    wire N__84042;
    wire N__84041;
    wire N__84040;
    wire N__84039;
    wire N__84038;
    wire N__84037;
    wire N__84036;
    wire N__84035;
    wire N__84034;
    wire N__84033;
    wire N__84032;
    wire N__84031;
    wire N__84030;
    wire N__84029;
    wire N__84028;
    wire N__84027;
    wire N__84026;
    wire N__84025;
    wire N__84024;
    wire N__84023;
    wire N__84022;
    wire N__84021;
    wire N__84020;
    wire N__84019;
    wire N__84018;
    wire N__84017;
    wire N__84016;
    wire N__84015;
    wire N__84014;
    wire N__84013;
    wire N__84012;
    wire N__84011;
    wire N__84010;
    wire N__84009;
    wire N__84008;
    wire N__84007;
    wire N__84006;
    wire N__84005;
    wire N__84004;
    wire N__84003;
    wire N__84002;
    wire N__84001;
    wire N__84000;
    wire N__83999;
    wire N__83998;
    wire N__83997;
    wire N__83996;
    wire N__83995;
    wire N__83994;
    wire N__83993;
    wire N__83992;
    wire N__83991;
    wire N__83990;
    wire N__83989;
    wire N__83988;
    wire N__83987;
    wire N__83986;
    wire N__83985;
    wire N__83984;
    wire N__83983;
    wire N__83982;
    wire N__83981;
    wire N__83980;
    wire N__83979;
    wire N__83978;
    wire N__83977;
    wire N__83976;
    wire N__83975;
    wire N__83974;
    wire N__83973;
    wire N__83972;
    wire N__83971;
    wire N__83970;
    wire N__83969;
    wire N__83968;
    wire N__83967;
    wire N__83966;
    wire N__83965;
    wire N__83964;
    wire N__83963;
    wire N__83962;
    wire N__83961;
    wire N__83960;
    wire N__83959;
    wire N__83958;
    wire N__83957;
    wire N__83956;
    wire N__83955;
    wire N__83954;
    wire N__83953;
    wire N__83952;
    wire N__83951;
    wire N__83950;
    wire N__83949;
    wire N__83948;
    wire N__83947;
    wire N__83946;
    wire N__83945;
    wire N__83944;
    wire N__83943;
    wire N__83942;
    wire N__83941;
    wire N__83940;
    wire N__83939;
    wire N__83938;
    wire N__83937;
    wire N__83936;
    wire N__83935;
    wire N__83934;
    wire N__83933;
    wire N__83932;
    wire N__83931;
    wire N__83930;
    wire N__83929;
    wire N__83928;
    wire N__83927;
    wire N__83926;
    wire N__83925;
    wire N__83924;
    wire N__83923;
    wire N__83922;
    wire N__83921;
    wire N__83920;
    wire N__83919;
    wire N__83918;
    wire N__83917;
    wire N__83916;
    wire N__83915;
    wire N__83914;
    wire N__83913;
    wire N__83912;
    wire N__83911;
    wire N__83910;
    wire N__83909;
    wire N__83908;
    wire N__83907;
    wire N__83906;
    wire N__83905;
    wire N__83904;
    wire N__83903;
    wire N__83902;
    wire N__83901;
    wire N__83900;
    wire N__83899;
    wire N__83898;
    wire N__83897;
    wire N__83896;
    wire N__83895;
    wire N__83894;
    wire N__83893;
    wire N__83892;
    wire N__83891;
    wire N__83890;
    wire N__83889;
    wire N__83888;
    wire N__83887;
    wire N__83886;
    wire N__83885;
    wire N__83884;
    wire N__83883;
    wire N__83882;
    wire N__83881;
    wire N__83880;
    wire N__83879;
    wire N__83878;
    wire N__83877;
    wire N__83876;
    wire N__83875;
    wire N__83874;
    wire N__83873;
    wire N__83872;
    wire N__83871;
    wire N__83870;
    wire N__83869;
    wire N__83868;
    wire N__83867;
    wire N__83866;
    wire N__83865;
    wire N__83864;
    wire N__83863;
    wire N__83862;
    wire N__83861;
    wire N__83860;
    wire N__83859;
    wire N__83858;
    wire N__83857;
    wire N__83856;
    wire N__83855;
    wire N__83854;
    wire N__83853;
    wire N__83852;
    wire N__83851;
    wire N__83850;
    wire N__83849;
    wire N__83848;
    wire N__83847;
    wire N__83846;
    wire N__83845;
    wire N__83844;
    wire N__83843;
    wire N__83842;
    wire N__83841;
    wire N__83840;
    wire N__83839;
    wire N__83838;
    wire N__83837;
    wire N__83836;
    wire N__83835;
    wire N__83834;
    wire N__83833;
    wire N__83832;
    wire N__83831;
    wire N__83830;
    wire N__83829;
    wire N__83828;
    wire N__83827;
    wire N__83826;
    wire N__83825;
    wire N__83824;
    wire N__83823;
    wire N__83822;
    wire N__83821;
    wire N__83820;
    wire N__83819;
    wire N__83818;
    wire N__83817;
    wire N__83816;
    wire N__83815;
    wire N__83214;
    wire N__83211;
    wire N__83208;
    wire N__83205;
    wire N__83204;
    wire N__83203;
    wire N__83202;
    wire N__83201;
    wire N__83198;
    wire N__83195;
    wire N__83192;
    wire N__83189;
    wire N__83188;
    wire N__83185;
    wire N__83184;
    wire N__83183;
    wire N__83182;
    wire N__83175;
    wire N__83172;
    wire N__83169;
    wire N__83166;
    wire N__83163;
    wire N__83160;
    wire N__83157;
    wire N__83156;
    wire N__83149;
    wire N__83146;
    wire N__83141;
    wire N__83138;
    wire N__83135;
    wire N__83134;
    wire N__83133;
    wire N__83132;
    wire N__83131;
    wire N__83128;
    wire N__83119;
    wire N__83116;
    wire N__83113;
    wire N__83110;
    wire N__83107;
    wire N__83106;
    wire N__83103;
    wire N__83100;
    wire N__83097;
    wire N__83094;
    wire N__83091;
    wire N__83090;
    wire N__83087;
    wire N__83084;
    wire N__83077;
    wire N__83072;
    wire N__83069;
    wire N__83066;
    wire N__83063;
    wire N__83056;
    wire N__83051;
    wire N__83048;
    wire N__83043;
    wire N__83042;
    wire N__83041;
    wire N__83040;
    wire N__83039;
    wire N__83038;
    wire N__83037;
    wire N__83036;
    wire N__83035;
    wire N__83034;
    wire N__83033;
    wire N__83032;
    wire N__83031;
    wire N__83030;
    wire N__83029;
    wire N__83028;
    wire N__83027;
    wire N__83026;
    wire N__83025;
    wire N__83024;
    wire N__83023;
    wire N__83022;
    wire N__83021;
    wire N__83020;
    wire N__83019;
    wire N__83018;
    wire N__83017;
    wire N__83016;
    wire N__83015;
    wire N__83014;
    wire N__83013;
    wire N__83012;
    wire N__83011;
    wire N__83010;
    wire N__83009;
    wire N__83008;
    wire N__83007;
    wire N__83006;
    wire N__83005;
    wire N__83004;
    wire N__83003;
    wire N__83002;
    wire N__83001;
    wire N__82990;
    wire N__82985;
    wire N__82968;
    wire N__82965;
    wire N__82962;
    wire N__82959;
    wire N__82956;
    wire N__82951;
    wire N__82936;
    wire N__82933;
    wire N__82928;
    wire N__82925;
    wire N__82916;
    wire N__82913;
    wire N__82910;
    wire N__82907;
    wire N__82904;
    wire N__82901;
    wire N__82898;
    wire N__82895;
    wire N__82894;
    wire N__82893;
    wire N__82892;
    wire N__82891;
    wire N__82890;
    wire N__82889;
    wire N__82888;
    wire N__82887;
    wire N__82886;
    wire N__82885;
    wire N__82884;
    wire N__82883;
    wire N__82882;
    wire N__82881;
    wire N__82880;
    wire N__82879;
    wire N__82878;
    wire N__82877;
    wire N__82876;
    wire N__82875;
    wire N__82874;
    wire N__82873;
    wire N__82872;
    wire N__82871;
    wire N__82870;
    wire N__82869;
    wire N__82868;
    wire N__82867;
    wire N__82866;
    wire N__82865;
    wire N__82864;
    wire N__82863;
    wire N__82862;
    wire N__82861;
    wire N__82860;
    wire N__82859;
    wire N__82858;
    wire N__82857;
    wire N__82856;
    wire N__82855;
    wire N__82854;
    wire N__82853;
    wire N__82852;
    wire N__82851;
    wire N__82850;
    wire N__82849;
    wire N__82846;
    wire N__82843;
    wire N__82840;
    wire N__82837;
    wire N__82834;
    wire N__82831;
    wire N__82828;
    wire N__82825;
    wire N__82822;
    wire N__82819;
    wire N__82816;
    wire N__82813;
    wire N__82810;
    wire N__82807;
    wire N__82804;
    wire N__82801;
    wire N__82798;
    wire N__82795;
    wire N__82792;
    wire N__82789;
    wire N__82656;
    wire N__82653;
    wire N__82650;
    wire N__82647;
    wire N__82644;
    wire N__82641;
    wire N__82640;
    wire N__82637;
    wire N__82634;
    wire N__82633;
    wire N__82632;
    wire N__82627;
    wire N__82624;
    wire N__82621;
    wire N__82620;
    wire N__82619;
    wire N__82618;
    wire N__82617;
    wire N__82614;
    wire N__82609;
    wire N__82604;
    wire N__82599;
    wire N__82590;
    wire N__82587;
    wire N__82584;
    wire N__82583;
    wire N__82582;
    wire N__82579;
    wire N__82576;
    wire N__82573;
    wire N__82572;
    wire N__82569;
    wire N__82566;
    wire N__82561;
    wire N__82558;
    wire N__82553;
    wire N__82548;
    wire N__82545;
    wire N__82542;
    wire N__82541;
    wire N__82536;
    wire N__82535;
    wire N__82532;
    wire N__82529;
    wire N__82524;
    wire N__82521;
    wire N__82518;
    wire N__82515;
    wire N__82514;
    wire N__82513;
    wire N__82506;
    wire N__82503;
    wire N__82500;
    wire N__82497;
    wire N__82494;
    wire N__82491;
    wire N__82488;
    wire N__82487;
    wire N__82482;
    wire N__82479;
    wire N__82476;
    wire N__82475;
    wire N__82472;
    wire N__82469;
    wire N__82464;
    wire N__82461;
    wire N__82460;
    wire N__82459;
    wire N__82458;
    wire N__82457;
    wire N__82456;
    wire N__82455;
    wire N__82454;
    wire N__82453;
    wire N__82452;
    wire N__82451;
    wire N__82448;
    wire N__82445;
    wire N__82442;
    wire N__82439;
    wire N__82436;
    wire N__82433;
    wire N__82432;
    wire N__82431;
    wire N__82428;
    wire N__82425;
    wire N__82422;
    wire N__82419;
    wire N__82416;
    wire N__82415;
    wire N__82414;
    wire N__82409;
    wire N__82406;
    wire N__82403;
    wire N__82400;
    wire N__82397;
    wire N__82394;
    wire N__82391;
    wire N__82386;
    wire N__82383;
    wire N__82380;
    wire N__82377;
    wire N__82374;
    wire N__82371;
    wire N__82368;
    wire N__82363;
    wire N__82354;
    wire N__82343;
    wire N__82340;
    wire N__82337;
    wire N__82332;
    wire N__82327;
    wire N__82320;
    wire N__82317;
    wire N__82314;
    wire N__82311;
    wire N__82308;
    wire N__82307;
    wire N__82302;
    wire N__82299;
    wire N__82298;
    wire N__82297;
    wire N__82294;
    wire N__82289;
    wire N__82286;
    wire N__82283;
    wire N__82280;
    wire N__82277;
    wire N__82272;
    wire N__82269;
    wire N__82266;
    wire N__82263;
    wire N__82260;
    wire N__82259;
    wire N__82258;
    wire N__82251;
    wire N__82248;
    wire N__82245;
    wire N__82242;
    wire N__82239;
    wire N__82236;
    wire N__82233;
    wire N__82230;
    wire N__82229;
    wire N__82228;
    wire N__82223;
    wire N__82220;
    wire N__82217;
    wire N__82214;
    wire N__82211;
    wire N__82208;
    wire N__82205;
    wire N__82202;
    wire N__82199;
    wire N__82196;
    wire N__82191;
    wire N__82190;
    wire N__82187;
    wire N__82184;
    wire N__82179;
    wire N__82176;
    wire N__82173;
    wire N__82172;
    wire N__82169;
    wire N__82166;
    wire N__82161;
    wire N__82158;
    wire N__82157;
    wire N__82154;
    wire N__82151;
    wire N__82146;
    wire N__82143;
    wire N__82140;
    wire N__82137;
    wire N__82134;
    wire N__82131;
    wire N__82128;
    wire N__82127;
    wire N__82126;
    wire N__82123;
    wire N__82118;
    wire N__82113;
    wire N__82112;
    wire N__82107;
    wire N__82104;
    wire N__82101;
    wire N__82100;
    wire N__82099;
    wire N__82096;
    wire N__82091;
    wire N__82086;
    wire N__82085;
    wire N__82084;
    wire N__82079;
    wire N__82076;
    wire N__82071;
    wire N__82070;
    wire N__82069;
    wire N__82066;
    wire N__82063;
    wire N__82060;
    wire N__82059;
    wire N__82056;
    wire N__82051;
    wire N__82048;
    wire N__82043;
    wire N__82038;
    wire N__82035;
    wire N__82032;
    wire N__82029;
    wire N__82026;
    wire N__82025;
    wire N__82024;
    wire N__82019;
    wire N__82016;
    wire N__82011;
    wire N__82008;
    wire N__82005;
    wire N__82004;
    wire N__82001;
    wire N__81998;
    wire N__81995;
    wire N__81992;
    wire N__81987;
    wire N__81984;
    wire N__81981;
    wire N__81980;
    wire N__81977;
    wire N__81974;
    wire N__81971;
    wire N__81966;
    wire N__81963;
    wire N__81962;
    wire N__81959;
    wire N__81956;
    wire N__81951;
    wire N__81948;
    wire N__81945;
    wire N__81942;
    wire N__81939;
    wire N__81936;
    wire N__81935;
    wire N__81930;
    wire N__81929;
    wire N__81928;
    wire N__81927;
    wire N__81924;
    wire N__81917;
    wire N__81914;
    wire N__81911;
    wire N__81906;
    wire N__81903;
    wire N__81900;
    wire N__81899;
    wire N__81898;
    wire N__81895;
    wire N__81890;
    wire N__81889;
    wire N__81888;
    wire N__81887;
    wire N__81882;
    wire N__81875;
    wire N__81872;
    wire N__81869;
    wire N__81864;
    wire N__81861;
    wire N__81858;
    wire N__81855;
    wire N__81852;
    wire N__81851;
    wire N__81848;
    wire N__81845;
    wire N__81842;
    wire N__81839;
    wire N__81838;
    wire N__81837;
    wire N__81836;
    wire N__81833;
    wire N__81830;
    wire N__81823;
    wire N__81816;
    wire N__81813;
    wire N__81810;
    wire N__81809;
    wire N__81808;
    wire N__81805;
    wire N__81802;
    wire N__81799;
    wire N__81794;
    wire N__81791;
    wire N__81788;
    wire N__81783;
    wire N__81780;
    wire N__81777;
    wire N__81774;
    wire N__81773;
    wire N__81770;
    wire N__81767;
    wire N__81764;
    wire N__81759;
    wire N__81756;
    wire N__81753;
    wire N__81750;
    wire N__81747;
    wire N__81744;
    wire N__81741;
    wire N__81738;
    wire N__81735;
    wire N__81734;
    wire N__81731;
    wire N__81728;
    wire N__81723;
    wire N__81720;
    wire N__81717;
    wire N__81714;
    wire N__81711;
    wire N__81708;
    wire N__81705;
    wire N__81704;
    wire N__81703;
    wire N__81700;
    wire N__81697;
    wire N__81694;
    wire N__81691;
    wire N__81688;
    wire N__81683;
    wire N__81680;
    wire N__81675;
    wire N__81672;
    wire N__81669;
    wire N__81666;
    wire N__81665;
    wire N__81664;
    wire N__81657;
    wire N__81654;
    wire N__81651;
    wire N__81648;
    wire N__81645;
    wire N__81644;
    wire N__81643;
    wire N__81636;
    wire N__81633;
    wire N__81630;
    wire N__81627;
    wire N__81624;
    wire N__81621;
    wire N__81620;
    wire N__81619;
    wire N__81612;
    wire N__81609;
    wire N__81606;
    wire N__81603;
    wire N__81600;
    wire N__81597;
    wire N__81594;
    wire N__81593;
    wire N__81592;
    wire N__81591;
    wire N__81588;
    wire N__81587;
    wire N__81586;
    wire N__81585;
    wire N__81578;
    wire N__81575;
    wire N__81574;
    wire N__81573;
    wire N__81572;
    wire N__81571;
    wire N__81570;
    wire N__81563;
    wire N__81558;
    wire N__81553;
    wire N__81550;
    wire N__81547;
    wire N__81544;
    wire N__81543;
    wire N__81542;
    wire N__81539;
    wire N__81534;
    wire N__81523;
    wire N__81520;
    wire N__81517;
    wire N__81514;
    wire N__81511;
    wire N__81508;
    wire N__81505;
    wire N__81498;
    wire N__81495;
    wire N__81492;
    wire N__81489;
    wire N__81488;
    wire N__81483;
    wire N__81480;
    wire N__81477;
    wire N__81474;
    wire N__81471;
    wire N__81468;
    wire N__81465;
    wire N__81464;
    wire N__81459;
    wire N__81456;
    wire N__81453;
    wire N__81450;
    wire N__81447;
    wire N__81444;
    wire N__81441;
    wire N__81438;
    wire N__81435;
    wire N__81434;
    wire N__81429;
    wire N__81426;
    wire N__81423;
    wire N__81420;
    wire N__81417;
    wire N__81414;
    wire N__81411;
    wire N__81408;
    wire N__81407;
    wire N__81404;
    wire N__81401;
    wire N__81396;
    wire N__81393;
    wire N__81390;
    wire N__81387;
    wire N__81384;
    wire N__81383;
    wire N__81378;
    wire N__81375;
    wire N__81372;
    wire N__81369;
    wire N__81366;
    wire N__81363;
    wire N__81362;
    wire N__81359;
    wire N__81354;
    wire N__81351;
    wire N__81348;
    wire N__81345;
    wire N__81342;
    wire N__81339;
    wire N__81336;
    wire N__81335;
    wire N__81330;
    wire N__81327;
    wire N__81324;
    wire N__81321;
    wire N__81318;
    wire N__81315;
    wire N__81312;
    wire N__81309;
    wire N__81308;
    wire N__81305;
    wire N__81304;
    wire N__81303;
    wire N__81300;
    wire N__81297;
    wire N__81296;
    wire N__81295;
    wire N__81292;
    wire N__81289;
    wire N__81288;
    wire N__81285;
    wire N__81282;
    wire N__81279;
    wire N__81276;
    wire N__81269;
    wire N__81258;
    wire N__81257;
    wire N__81256;
    wire N__81253;
    wire N__81250;
    wire N__81249;
    wire N__81248;
    wire N__81247;
    wire N__81244;
    wire N__81243;
    wire N__81240;
    wire N__81237;
    wire N__81234;
    wire N__81231;
    wire N__81230;
    wire N__81227;
    wire N__81224;
    wire N__81221;
    wire N__81216;
    wire N__81211;
    wire N__81208;
    wire N__81205;
    wire N__81200;
    wire N__81199;
    wire N__81192;
    wire N__81191;
    wire N__81190;
    wire N__81189;
    wire N__81186;
    wire N__81183;
    wire N__81180;
    wire N__81177;
    wire N__81174;
    wire N__81171;
    wire N__81168;
    wire N__81153;
    wire N__81150;
    wire N__81149;
    wire N__81148;
    wire N__81147;
    wire N__81146;
    wire N__81145;
    wire N__81144;
    wire N__81143;
    wire N__81142;
    wire N__81141;
    wire N__81140;
    wire N__81139;
    wire N__81138;
    wire N__81135;
    wire N__81108;
    wire N__81105;
    wire N__81102;
    wire N__81101;
    wire N__81100;
    wire N__81097;
    wire N__81094;
    wire N__81093;
    wire N__81090;
    wire N__81087;
    wire N__81086;
    wire N__81085;
    wire N__81082;
    wire N__81081;
    wire N__81080;
    wire N__81077;
    wire N__81076;
    wire N__81075;
    wire N__81072;
    wire N__81069;
    wire N__81066;
    wire N__81063;
    wire N__81060;
    wire N__81059;
    wire N__81056;
    wire N__81053;
    wire N__81050;
    wire N__81047;
    wire N__81044;
    wire N__81041;
    wire N__81038;
    wire N__81035;
    wire N__81032;
    wire N__81029;
    wire N__81026;
    wire N__81023;
    wire N__81020;
    wire N__81017;
    wire N__81014;
    wire N__81011;
    wire N__81010;
    wire N__81007;
    wire N__81000;
    wire N__80997;
    wire N__80992;
    wire N__80989;
    wire N__80986;
    wire N__80983;
    wire N__80982;
    wire N__80979;
    wire N__80976;
    wire N__80971;
    wire N__80964;
    wire N__80959;
    wire N__80956;
    wire N__80943;
    wire N__80940;
    wire N__80939;
    wire N__80936;
    wire N__80933;
    wire N__80930;
    wire N__80927;
    wire N__80922;
    wire N__80919;
    wire N__80918;
    wire N__80915;
    wire N__80914;
    wire N__80913;
    wire N__80912;
    wire N__80909;
    wire N__80906;
    wire N__80903;
    wire N__80900;
    wire N__80897;
    wire N__80894;
    wire N__80891;
    wire N__80886;
    wire N__80883;
    wire N__80878;
    wire N__80875;
    wire N__80872;
    wire N__80869;
    wire N__80866;
    wire N__80863;
    wire N__80858;
    wire N__80855;
    wire N__80852;
    wire N__80849;
    wire N__80844;
    wire N__80841;
    wire N__80838;
    wire N__80835;
    wire N__80834;
    wire N__80833;
    wire N__80832;
    wire N__80831;
    wire N__80830;
    wire N__80827;
    wire N__80822;
    wire N__80815;
    wire N__80814;
    wire N__80813;
    wire N__80812;
    wire N__80811;
    wire N__80810;
    wire N__80809;
    wire N__80808;
    wire N__80807;
    wire N__80806;
    wire N__80799;
    wire N__80788;
    wire N__80779;
    wire N__80774;
    wire N__80771;
    wire N__80768;
    wire N__80765;
    wire N__80762;
    wire N__80759;
    wire N__80756;
    wire N__80753;
    wire N__80748;
    wire N__80745;
    wire N__80742;
    wire N__80739;
    wire N__80738;
    wire N__80737;
    wire N__80734;
    wire N__80729;
    wire N__80726;
    wire N__80723;
    wire N__80720;
    wire N__80717;
    wire N__80714;
    wire N__80711;
    wire N__80706;
    wire N__80703;
    wire N__80700;
    wire N__80697;
    wire N__80696;
    wire N__80693;
    wire N__80690;
    wire N__80687;
    wire N__80682;
    wire N__80679;
    wire N__80676;
    wire N__80673;
    wire N__80670;
    wire N__80669;
    wire N__80664;
    wire N__80661;
    wire N__80658;
    wire N__80655;
    wire N__80652;
    wire N__80651;
    wire N__80646;
    wire N__80643;
    wire N__80640;
    wire N__80637;
    wire N__80636;
    wire N__80633;
    wire N__80630;
    wire N__80627;
    wire N__80624;
    wire N__80619;
    wire N__80616;
    wire N__80615;
    wire N__80612;
    wire N__80609;
    wire N__80604;
    wire N__80601;
    wire N__80598;
    wire N__80595;
    wire N__80592;
    wire N__80589;
    wire N__80586;
    wire N__80585;
    wire N__80582;
    wire N__80579;
    wire N__80574;
    wire N__80571;
    wire N__80568;
    wire N__80567;
    wire N__80562;
    wire N__80559;
    wire N__80556;
    wire N__80553;
    wire N__80550;
    wire N__80547;
    wire N__80546;
    wire N__80545;
    wire N__80542;
    wire N__80539;
    wire N__80536;
    wire N__80529;
    wire N__80526;
    wire N__80523;
    wire N__80520;
    wire N__80517;
    wire N__80516;
    wire N__80515;
    wire N__80514;
    wire N__80511;
    wire N__80510;
    wire N__80509;
    wire N__80506;
    wire N__80505;
    wire N__80504;
    wire N__80501;
    wire N__80500;
    wire N__80497;
    wire N__80494;
    wire N__80493;
    wire N__80488;
    wire N__80485;
    wire N__80482;
    wire N__80481;
    wire N__80478;
    wire N__80475;
    wire N__80472;
    wire N__80471;
    wire N__80468;
    wire N__80467;
    wire N__80464;
    wire N__80463;
    wire N__80460;
    wire N__80457;
    wire N__80454;
    wire N__80451;
    wire N__80448;
    wire N__80445;
    wire N__80440;
    wire N__80437;
    wire N__80434;
    wire N__80433;
    wire N__80432;
    wire N__80429;
    wire N__80426;
    wire N__80423;
    wire N__80420;
    wire N__80417;
    wire N__80414;
    wire N__80413;
    wire N__80412;
    wire N__80409;
    wire N__80404;
    wire N__80401;
    wire N__80396;
    wire N__80395;
    wire N__80390;
    wire N__80381;
    wire N__80376;
    wire N__80373;
    wire N__80370;
    wire N__80367;
    wire N__80362;
    wire N__80359;
    wire N__80356;
    wire N__80347;
    wire N__80334;
    wire N__80331;
    wire N__80330;
    wire N__80327;
    wire N__80324;
    wire N__80321;
    wire N__80318;
    wire N__80313;
    wire N__80310;
    wire N__80309;
    wire N__80308;
    wire N__80307;
    wire N__80298;
    wire N__80297;
    wire N__80296;
    wire N__80295;
    wire N__80292;
    wire N__80291;
    wire N__80288;
    wire N__80285;
    wire N__80282;
    wire N__80279;
    wire N__80276;
    wire N__80275;
    wire N__80272;
    wire N__80269;
    wire N__80266;
    wire N__80263;
    wire N__80262;
    wire N__80259;
    wire N__80258;
    wire N__80255;
    wire N__80250;
    wire N__80249;
    wire N__80248;
    wire N__80245;
    wire N__80242;
    wire N__80239;
    wire N__80238;
    wire N__80235;
    wire N__80232;
    wire N__80229;
    wire N__80226;
    wire N__80223;
    wire N__80220;
    wire N__80217;
    wire N__80212;
    wire N__80209;
    wire N__80206;
    wire N__80205;
    wire N__80204;
    wire N__80203;
    wire N__80200;
    wire N__80199;
    wire N__80196;
    wire N__80191;
    wire N__80188;
    wire N__80187;
    wire N__80178;
    wire N__80173;
    wire N__80170;
    wire N__80167;
    wire N__80164;
    wire N__80161;
    wire N__80156;
    wire N__80153;
    wire N__80146;
    wire N__80133;
    wire N__80130;
    wire N__80129;
    wire N__80126;
    wire N__80123;
    wire N__80120;
    wire N__80117;
    wire N__80112;
    wire N__80109;
    wire N__80108;
    wire N__80107;
    wire N__80106;
    wire N__80105;
    wire N__80104;
    wire N__80101;
    wire N__80100;
    wire N__80099;
    wire N__80096;
    wire N__80093;
    wire N__80090;
    wire N__80089;
    wire N__80088;
    wire N__80085;
    wire N__80082;
    wire N__80081;
    wire N__80078;
    wire N__80075;
    wire N__80074;
    wire N__80071;
    wire N__80068;
    wire N__80063;
    wire N__80060;
    wire N__80057;
    wire N__80052;
    wire N__80049;
    wire N__80046;
    wire N__80045;
    wire N__80044;
    wire N__80041;
    wire N__80038;
    wire N__80037;
    wire N__80034;
    wire N__80031;
    wire N__80028;
    wire N__80025;
    wire N__80022;
    wire N__80019;
    wire N__80014;
    wire N__80009;
    wire N__80004;
    wire N__80003;
    wire N__80000;
    wire N__79995;
    wire N__79990;
    wire N__79983;
    wire N__79978;
    wire N__79975;
    wire N__79962;
    wire N__79961;
    wire N__79958;
    wire N__79955;
    wire N__79952;
    wire N__79949;
    wire N__79946;
    wire N__79943;
    wire N__79938;
    wire N__79935;
    wire N__79932;
    wire N__79931;
    wire N__79930;
    wire N__79927;
    wire N__79924;
    wire N__79921;
    wire N__79918;
    wire N__79915;
    wire N__79910;
    wire N__79909;
    wire N__79908;
    wire N__79905;
    wire N__79902;
    wire N__79899;
    wire N__79896;
    wire N__79893;
    wire N__79892;
    wire N__79891;
    wire N__79890;
    wire N__79889;
    wire N__79888;
    wire N__79885;
    wire N__79882;
    wire N__79877;
    wire N__79874;
    wire N__79871;
    wire N__79870;
    wire N__79867;
    wire N__79866;
    wire N__79865;
    wire N__79864;
    wire N__79861;
    wire N__79858;
    wire N__79857;
    wire N__79852;
    wire N__79847;
    wire N__79844;
    wire N__79841;
    wire N__79838;
    wire N__79837;
    wire N__79832;
    wire N__79829;
    wire N__79826;
    wire N__79823;
    wire N__79820;
    wire N__79817;
    wire N__79814;
    wire N__79809;
    wire N__79806;
    wire N__79803;
    wire N__79800;
    wire N__79797;
    wire N__79794;
    wire N__79791;
    wire N__79784;
    wire N__79779;
    wire N__79776;
    wire N__79771;
    wire N__79758;
    wire N__79755;
    wire N__79754;
    wire N__79751;
    wire N__79748;
    wire N__79745;
    wire N__79742;
    wire N__79737;
    wire N__79734;
    wire N__79731;
    wire N__79730;
    wire N__79727;
    wire N__79726;
    wire N__79725;
    wire N__79724;
    wire N__79721;
    wire N__79720;
    wire N__79717;
    wire N__79716;
    wire N__79715;
    wire N__79714;
    wire N__79713;
    wire N__79710;
    wire N__79707;
    wire N__79704;
    wire N__79701;
    wire N__79698;
    wire N__79697;
    wire N__79694;
    wire N__79691;
    wire N__79688;
    wire N__79685;
    wire N__79684;
    wire N__79681;
    wire N__79678;
    wire N__79675;
    wire N__79672;
    wire N__79669;
    wire N__79666;
    wire N__79663;
    wire N__79658;
    wire N__79655;
    wire N__79652;
    wire N__79649;
    wire N__79644;
    wire N__79641;
    wire N__79636;
    wire N__79631;
    wire N__79630;
    wire N__79623;
    wire N__79618;
    wire N__79611;
    wire N__79608;
    wire N__79599;
    wire N__79596;
    wire N__79595;
    wire N__79592;
    wire N__79589;
    wire N__79586;
    wire N__79583;
    wire N__79578;
    wire N__79575;
    wire N__79572;
    wire N__79569;
    wire N__79566;
    wire N__79563;
    wire N__79562;
    wire N__79561;
    wire N__79554;
    wire N__79551;
    wire N__79548;
    wire N__79545;
    wire N__79542;
    wire N__79539;
    wire N__79536;
    wire N__79533;
    wire N__79530;
    wire N__79527;
    wire N__79526;
    wire N__79523;
    wire N__79522;
    wire N__79519;
    wire N__79516;
    wire N__79513;
    wire N__79510;
    wire N__79503;
    wire N__79502;
    wire N__79499;
    wire N__79496;
    wire N__79491;
    wire N__79490;
    wire N__79485;
    wire N__79482;
    wire N__79479;
    wire N__79478;
    wire N__79473;
    wire N__79470;
    wire N__79467;
    wire N__79466;
    wire N__79463;
    wire N__79460;
    wire N__79457;
    wire N__79454;
    wire N__79449;
    wire N__79446;
    wire N__79445;
    wire N__79442;
    wire N__79439;
    wire N__79436;
    wire N__79433;
    wire N__79430;
    wire N__79427;
    wire N__79422;
    wire N__79419;
    wire N__79416;
    wire N__79415;
    wire N__79412;
    wire N__79411;
    wire N__79410;
    wire N__79407;
    wire N__79406;
    wire N__79403;
    wire N__79398;
    wire N__79395;
    wire N__79392;
    wire N__79383;
    wire N__79380;
    wire N__79377;
    wire N__79374;
    wire N__79371;
    wire N__79370;
    wire N__79369;
    wire N__79364;
    wire N__79361;
    wire N__79358;
    wire N__79353;
    wire N__79350;
    wire N__79347;
    wire N__79344;
    wire N__79341;
    wire N__79338;
    wire N__79337;
    wire N__79334;
    wire N__79331;
    wire N__79328;
    wire N__79323;
    wire N__79320;
    wire N__79317;
    wire N__79316;
    wire N__79313;
    wire N__79310;
    wire N__79305;
    wire N__79302;
    wire N__79299;
    wire N__79296;
    wire N__79293;
    wire N__79290;
    wire N__79289;
    wire N__79288;
    wire N__79285;
    wire N__79284;
    wire N__79281;
    wire N__79278;
    wire N__79277;
    wire N__79276;
    wire N__79275;
    wire N__79272;
    wire N__79269;
    wire N__79268;
    wire N__79265;
    wire N__79262;
    wire N__79259;
    wire N__79258;
    wire N__79255;
    wire N__79252;
    wire N__79249;
    wire N__79246;
    wire N__79243;
    wire N__79242;
    wire N__79239;
    wire N__79234;
    wire N__79231;
    wire N__79228;
    wire N__79227;
    wire N__79224;
    wire N__79221;
    wire N__79216;
    wire N__79213;
    wire N__79208;
    wire N__79205;
    wire N__79202;
    wire N__79199;
    wire N__79198;
    wire N__79197;
    wire N__79192;
    wire N__79187;
    wire N__79184;
    wire N__79181;
    wire N__79176;
    wire N__79173;
    wire N__79170;
    wire N__79167;
    wire N__79160;
    wire N__79155;
    wire N__79146;
    wire N__79143;
    wire N__79142;
    wire N__79139;
    wire N__79136;
    wire N__79133;
    wire N__79130;
    wire N__79125;
    wire N__79122;
    wire N__79121;
    wire N__79116;
    wire N__79113;
    wire N__79110;
    wire N__79107;
    wire N__79106;
    wire N__79103;
    wire N__79100;
    wire N__79095;
    wire N__79094;
    wire N__79091;
    wire N__79088;
    wire N__79083;
    wire N__79082;
    wire N__79077;
    wire N__79074;
    wire N__79071;
    wire N__79068;
    wire N__79065;
    wire N__79064;
    wire N__79061;
    wire N__79058;
    wire N__79053;
    wire N__79050;
    wire N__79047;
    wire N__79044;
    wire N__79043;
    wire N__79040;
    wire N__79037;
    wire N__79032;
    wire N__79029;
    wire N__79026;
    wire N__79023;
    wire N__79022;
    wire N__79017;
    wire N__79014;
    wire N__79013;
    wire N__79008;
    wire N__79005;
    wire N__79002;
    wire N__78999;
    wire N__78998;
    wire N__78993;
    wire N__78990;
    wire N__78987;
    wire N__78984;
    wire N__78981;
    wire N__78978;
    wire N__78975;
    wire N__78974;
    wire N__78973;
    wire N__78970;
    wire N__78965;
    wire N__78964;
    wire N__78959;
    wire N__78956;
    wire N__78951;
    wire N__78950;
    wire N__78949;
    wire N__78946;
    wire N__78941;
    wire N__78938;
    wire N__78935;
    wire N__78930;
    wire N__78927;
    wire N__78924;
    wire N__78921;
    wire N__78918;
    wire N__78917;
    wire N__78914;
    wire N__78911;
    wire N__78908;
    wire N__78905;
    wire N__78900;
    wire N__78897;
    wire N__78894;
    wire N__78891;
    wire N__78888;
    wire N__78885;
    wire N__78882;
    wire N__78881;
    wire N__78880;
    wire N__78879;
    wire N__78876;
    wire N__78869;
    wire N__78864;
    wire N__78863;
    wire N__78860;
    wire N__78857;
    wire N__78856;
    wire N__78849;
    wire N__78846;
    wire N__78843;
    wire N__78840;
    wire N__78837;
    wire N__78834;
    wire N__78831;
    wire N__78830;
    wire N__78829;
    wire N__78828;
    wire N__78825;
    wire N__78822;
    wire N__78821;
    wire N__78818;
    wire N__78817;
    wire N__78814;
    wire N__78809;
    wire N__78802;
    wire N__78795;
    wire N__78792;
    wire N__78789;
    wire N__78786;
    wire N__78783;
    wire N__78780;
    wire N__78777;
    wire N__78774;
    wire N__78771;
    wire N__78770;
    wire N__78769;
    wire N__78768;
    wire N__78767;
    wire N__78766;
    wire N__78765;
    wire N__78762;
    wire N__78753;
    wire N__78750;
    wire N__78749;
    wire N__78746;
    wire N__78743;
    wire N__78738;
    wire N__78735;
    wire N__78728;
    wire N__78725;
    wire N__78722;
    wire N__78719;
    wire N__78716;
    wire N__78711;
    wire N__78708;
    wire N__78705;
    wire N__78702;
    wire N__78699;
    wire N__78698;
    wire N__78697;
    wire N__78696;
    wire N__78691;
    wire N__78686;
    wire N__78683;
    wire N__78680;
    wire N__78675;
    wire N__78672;
    wire N__78669;
    wire N__78666;
    wire N__78663;
    wire N__78660;
    wire N__78657;
    wire N__78656;
    wire N__78651;
    wire N__78648;
    wire N__78647;
    wire N__78644;
    wire N__78641;
    wire N__78636;
    wire N__78633;
    wire N__78630;
    wire N__78627;
    wire N__78624;
    wire N__78621;
    wire N__78620;
    wire N__78615;
    wire N__78614;
    wire N__78613;
    wire N__78610;
    wire N__78605;
    wire N__78600;
    wire N__78597;
    wire N__78594;
    wire N__78591;
    wire N__78588;
    wire N__78587;
    wire N__78586;
    wire N__78585;
    wire N__78584;
    wire N__78573;
    wire N__78570;
    wire N__78567;
    wire N__78564;
    wire N__78561;
    wire N__78558;
    wire N__78555;
    wire N__78552;
    wire N__78551;
    wire N__78550;
    wire N__78547;
    wire N__78544;
    wire N__78541;
    wire N__78538;
    wire N__78533;
    wire N__78528;
    wire N__78525;
    wire N__78522;
    wire N__78519;
    wire N__78516;
    wire N__78515;
    wire N__78510;
    wire N__78509;
    wire N__78508;
    wire N__78507;
    wire N__78506;
    wire N__78503;
    wire N__78494;
    wire N__78489;
    wire N__78486;
    wire N__78485;
    wire N__78482;
    wire N__78479;
    wire N__78474;
    wire N__78471;
    wire N__78468;
    wire N__78465;
    wire N__78462;
    wire N__78459;
    wire N__78458;
    wire N__78455;
    wire N__78452;
    wire N__78447;
    wire N__78444;
    wire N__78441;
    wire N__78438;
    wire N__78435;
    wire N__78432;
    wire N__78429;
    wire N__78426;
    wire N__78423;
    wire N__78420;
    wire N__78417;
    wire N__78416;
    wire N__78415;
    wire N__78414;
    wire N__78405;
    wire N__78402;
    wire N__78401;
    wire N__78396;
    wire N__78393;
    wire N__78390;
    wire N__78389;
    wire N__78384;
    wire N__78381;
    wire N__78380;
    wire N__78377;
    wire N__78374;
    wire N__78369;
    wire N__78368;
    wire N__78365;
    wire N__78362;
    wire N__78361;
    wire N__78360;
    wire N__78359;
    wire N__78358;
    wire N__78357;
    wire N__78356;
    wire N__78355;
    wire N__78354;
    wire N__78353;
    wire N__78352;
    wire N__78349;
    wire N__78346;
    wire N__78321;
    wire N__78318;
    wire N__78315;
    wire N__78314;
    wire N__78313;
    wire N__78312;
    wire N__78311;
    wire N__78308;
    wire N__78305;
    wire N__78298;
    wire N__78291;
    wire N__78290;
    wire N__78289;
    wire N__78288;
    wire N__78285;
    wire N__78278;
    wire N__78273;
    wire N__78270;
    wire N__78267;
    wire N__78266;
    wire N__78263;
    wire N__78260;
    wire N__78259;
    wire N__78256;
    wire N__78253;
    wire N__78250;
    wire N__78243;
    wire N__78240;
    wire N__78237;
    wire N__78234;
    wire N__78231;
    wire N__78230;
    wire N__78229;
    wire N__78228;
    wire N__78227;
    wire N__78224;
    wire N__78221;
    wire N__78216;
    wire N__78213;
    wire N__78204;
    wire N__78203;
    wire N__78202;
    wire N__78201;
    wire N__78200;
    wire N__78199;
    wire N__78198;
    wire N__78197;
    wire N__78196;
    wire N__78187;
    wire N__78186;
    wire N__78185;
    wire N__78184;
    wire N__78183;
    wire N__78182;
    wire N__78179;
    wire N__78178;
    wire N__78169;
    wire N__78166;
    wire N__78163;
    wire N__78154;
    wire N__78151;
    wire N__78148;
    wire N__78145;
    wire N__78138;
    wire N__78135;
    wire N__78130;
    wire N__78127;
    wire N__78124;
    wire N__78121;
    wire N__78118;
    wire N__78113;
    wire N__78110;
    wire N__78105;
    wire N__78102;
    wire N__78099;
    wire N__78096;
    wire N__78093;
    wire N__78090;
    wire N__78087;
    wire N__78084;
    wire N__78081;
    wire N__78078;
    wire N__78075;
    wire N__78072;
    wire N__78069;
    wire N__78066;
    wire N__78063;
    wire N__78060;
    wire N__78057;
    wire N__78054;
    wire N__78051;
    wire N__78048;
    wire N__78045;
    wire N__78042;
    wire N__78039;
    wire N__78036;
    wire N__78033;
    wire N__78030;
    wire N__78027;
    wire N__78024;
    wire N__78021;
    wire N__78018;
    wire N__78015;
    wire N__78012;
    wire N__78009;
    wire N__78006;
    wire N__78003;
    wire N__78000;
    wire N__77997;
    wire N__77994;
    wire N__77991;
    wire N__77988;
    wire N__77985;
    wire N__77982;
    wire N__77979;
    wire N__77976;
    wire N__77973;
    wire N__77970;
    wire N__77967;
    wire N__77964;
    wire N__77961;
    wire N__77958;
    wire N__77955;
    wire N__77952;
    wire N__77949;
    wire N__77948;
    wire N__77945;
    wire N__77942;
    wire N__77941;
    wire N__77938;
    wire N__77935;
    wire N__77932;
    wire N__77929;
    wire N__77926;
    wire N__77923;
    wire N__77918;
    wire N__77913;
    wire N__77910;
    wire N__77907;
    wire N__77906;
    wire N__77905;
    wire N__77904;
    wire N__77903;
    wire N__77902;
    wire N__77901;
    wire N__77898;
    wire N__77893;
    wire N__77884;
    wire N__77877;
    wire N__77874;
    wire N__77871;
    wire N__77868;
    wire N__77865;
    wire N__77862;
    wire N__77859;
    wire N__77856;
    wire N__77853;
    wire N__77850;
    wire N__77847;
    wire N__77844;
    wire N__77841;
    wire N__77838;
    wire N__77835;
    wire N__77832;
    wire N__77829;
    wire N__77826;
    wire N__77823;
    wire N__77820;
    wire N__77817;
    wire N__77814;
    wire N__77811;
    wire N__77808;
    wire N__77805;
    wire N__77802;
    wire N__77799;
    wire N__77796;
    wire N__77793;
    wire N__77790;
    wire N__77787;
    wire N__77784;
    wire N__77781;
    wire N__77778;
    wire N__77775;
    wire N__77772;
    wire N__77769;
    wire N__77766;
    wire N__77763;
    wire N__77760;
    wire N__77757;
    wire N__77754;
    wire N__77751;
    wire N__77748;
    wire N__77745;
    wire N__77742;
    wire N__77739;
    wire N__77736;
    wire N__77733;
    wire N__77730;
    wire N__77727;
    wire N__77724;
    wire N__77721;
    wire N__77718;
    wire N__77715;
    wire N__77712;
    wire N__77709;
    wire N__77706;
    wire N__77703;
    wire N__77700;
    wire N__77697;
    wire N__77694;
    wire N__77691;
    wire N__77688;
    wire N__77685;
    wire N__77682;
    wire N__77679;
    wire N__77676;
    wire N__77673;
    wire N__77670;
    wire N__77667;
    wire N__77666;
    wire N__77665;
    wire N__77664;
    wire N__77663;
    wire N__77662;
    wire N__77661;
    wire N__77660;
    wire N__77659;
    wire N__77658;
    wire N__77657;
    wire N__77656;
    wire N__77655;
    wire N__77654;
    wire N__77653;
    wire N__77650;
    wire N__77649;
    wire N__77648;
    wire N__77647;
    wire N__77646;
    wire N__77643;
    wire N__77642;
    wire N__77641;
    wire N__77640;
    wire N__77639;
    wire N__77638;
    wire N__77637;
    wire N__77636;
    wire N__77635;
    wire N__77634;
    wire N__77633;
    wire N__77632;
    wire N__77631;
    wire N__77630;
    wire N__77629;
    wire N__77628;
    wire N__77627;
    wire N__77626;
    wire N__77625;
    wire N__77624;
    wire N__77623;
    wire N__77622;
    wire N__77621;
    wire N__77620;
    wire N__77619;
    wire N__77618;
    wire N__77617;
    wire N__77616;
    wire N__77615;
    wire N__77614;
    wire N__77613;
    wire N__77612;
    wire N__77611;
    wire N__77610;
    wire N__77609;
    wire N__77608;
    wire N__77607;
    wire N__77606;
    wire N__77605;
    wire N__77604;
    wire N__77603;
    wire N__77602;
    wire N__77601;
    wire N__77600;
    wire N__77597;
    wire N__77594;
    wire N__77593;
    wire N__77592;
    wire N__77591;
    wire N__77590;
    wire N__77589;
    wire N__77588;
    wire N__77587;
    wire N__77586;
    wire N__77583;
    wire N__77580;
    wire N__77571;
    wire N__77568;
    wire N__77563;
    wire N__77560;
    wire N__77553;
    wire N__77546;
    wire N__77541;
    wire N__77534;
    wire N__77525;
    wire N__77522;
    wire N__77519;
    wire N__77516;
    wire N__77513;
    wire N__77510;
    wire N__77507;
    wire N__77500;
    wire N__77497;
    wire N__77492;
    wire N__77487;
    wire N__77484;
    wire N__77481;
    wire N__77478;
    wire N__77475;
    wire N__77472;
    wire N__77469;
    wire N__77462;
    wire N__77455;
    wire N__77452;
    wire N__77449;
    wire N__77446;
    wire N__77443;
    wire N__77440;
    wire N__77437;
    wire N__77434;
    wire N__77431;
    wire N__77422;
    wire N__77415;
    wire N__77412;
    wire N__77409;
    wire N__77406;
    wire N__77403;
    wire N__77402;
    wire N__77401;
    wire N__77400;
    wire N__77399;
    wire N__77398;
    wire N__77397;
    wire N__77396;
    wire N__77395;
    wire N__77394;
    wire N__77393;
    wire N__77392;
    wire N__77391;
    wire N__77390;
    wire N__77389;
    wire N__77388;
    wire N__77387;
    wire N__77386;
    wire N__77385;
    wire N__77384;
    wire N__77383;
    wire N__77382;
    wire N__77381;
    wire N__77380;
    wire N__77379;
    wire N__77378;
    wire N__77377;
    wire N__77376;
    wire N__77375;
    wire N__77374;
    wire N__77373;
    wire N__77372;
    wire N__77371;
    wire N__77370;
    wire N__77369;
    wire N__77368;
    wire N__77367;
    wire N__77366;
    wire N__77365;
    wire N__77364;
    wire N__77363;
    wire N__77362;
    wire N__77361;
    wire N__77360;
    wire N__77359;
    wire N__77358;
    wire N__77357;
    wire N__77356;
    wire N__77355;
    wire N__77354;
    wire N__77353;
    wire N__77352;
    wire N__77351;
    wire N__77350;
    wire N__77349;
    wire N__77348;
    wire N__77347;
    wire N__77346;
    wire N__77345;
    wire N__77344;
    wire N__77343;
    wire N__77342;
    wire N__77341;
    wire N__77340;
    wire N__77339;
    wire N__77338;
    wire N__77337;
    wire N__77336;
    wire N__77335;
    wire N__77334;
    wire N__77333;
    wire N__77332;
    wire N__77331;
    wire N__77330;
    wire N__77329;
    wire N__77328;
    wire N__77327;
    wire N__77326;
    wire N__77325;
    wire N__77324;
    wire N__77323;
    wire N__77322;
    wire N__77321;
    wire N__77320;
    wire N__77319;
    wire N__77318;
    wire N__77317;
    wire N__77316;
    wire N__77315;
    wire N__77314;
    wire N__77313;
    wire N__77312;
    wire N__77311;
    wire N__77310;
    wire N__77309;
    wire N__77308;
    wire N__77307;
    wire N__77306;
    wire N__77305;
    wire N__77304;
    wire N__77303;
    wire N__77302;
    wire N__77301;
    wire N__77300;
    wire N__77299;
    wire N__77298;
    wire N__77297;
    wire N__77296;
    wire N__77295;
    wire N__77294;
    wire N__77293;
    wire N__77292;
    wire N__77291;
    wire N__77290;
    wire N__77289;
    wire N__77288;
    wire N__77287;
    wire N__77286;
    wire N__77285;
    wire N__77284;
    wire N__77283;
    wire N__77282;
    wire N__77281;
    wire N__77280;
    wire N__77279;
    wire N__77278;
    wire N__77277;
    wire N__77276;
    wire N__77275;
    wire N__77274;
    wire N__77273;
    wire N__77272;
    wire N__77271;
    wire N__77270;
    wire N__77269;
    wire N__77268;
    wire N__77267;
    wire N__77266;
    wire N__77265;
    wire N__77264;
    wire N__77263;
    wire N__77262;
    wire N__77261;
    wire N__77260;
    wire N__77259;
    wire N__77258;
    wire N__77257;
    wire N__77256;
    wire N__77255;
    wire N__77254;
    wire N__77253;
    wire N__77252;
    wire N__77251;
    wire N__77250;
    wire N__77249;
    wire N__77248;
    wire N__77247;
    wire N__77246;
    wire N__77243;
    wire N__77240;
    wire N__77237;
    wire N__77234;
    wire N__77231;
    wire N__77228;
    wire N__77225;
    wire N__77222;
    wire N__77219;
    wire N__77216;
    wire N__77213;
    wire N__77210;
    wire N__77207;
    wire N__77204;
    wire N__77201;
    wire N__77198;
    wire N__77195;
    wire N__77192;
    wire N__77189;
    wire N__77186;
    wire N__77183;
    wire N__77180;
    wire N__77177;
    wire N__77174;
    wire N__77171;
    wire N__77168;
    wire N__77165;
    wire N__77162;
    wire N__77159;
    wire N__77156;
    wire N__77153;
    wire N__77150;
    wire N__77147;
    wire N__77144;
    wire N__77141;
    wire N__77138;
    wire N__77135;
    wire N__77132;
    wire N__77129;
    wire N__77126;
    wire N__77123;
    wire N__77120;
    wire N__77117;
    wire N__76716;
    wire N__76713;
    wire N__76710;
    wire N__76707;
    wire N__76704;
    wire N__76701;
    wire N__76698;
    wire N__76695;
    wire N__76694;
    wire N__76693;
    wire N__76690;
    wire N__76687;
    wire N__76684;
    wire N__76681;
    wire N__76674;
    wire N__76671;
    wire N__76670;
    wire N__76667;
    wire N__76664;
    wire N__76661;
    wire N__76658;
    wire N__76657;
    wire N__76654;
    wire N__76651;
    wire N__76648;
    wire N__76641;
    wire N__76640;
    wire N__76639;
    wire N__76638;
    wire N__76635;
    wire N__76634;
    wire N__76633;
    wire N__76632;
    wire N__76631;
    wire N__76630;
    wire N__76629;
    wire N__76628;
    wire N__76627;
    wire N__76626;
    wire N__76625;
    wire N__76624;
    wire N__76623;
    wire N__76622;
    wire N__76621;
    wire N__76620;
    wire N__76619;
    wire N__76618;
    wire N__76617;
    wire N__76616;
    wire N__76615;
    wire N__76614;
    wire N__76613;
    wire N__76612;
    wire N__76611;
    wire N__76610;
    wire N__76609;
    wire N__76608;
    wire N__76601;
    wire N__76596;
    wire N__76585;
    wire N__76576;
    wire N__76569;
    wire N__76568;
    wire N__76567;
    wire N__76566;
    wire N__76565;
    wire N__76564;
    wire N__76563;
    wire N__76560;
    wire N__76555;
    wire N__76548;
    wire N__76535;
    wire N__76534;
    wire N__76531;
    wire N__76530;
    wire N__76529;
    wire N__76528;
    wire N__76527;
    wire N__76524;
    wire N__76521;
    wire N__76518;
    wire N__76511;
    wire N__76502;
    wire N__76497;
    wire N__76494;
    wire N__76493;
    wire N__76492;
    wire N__76491;
    wire N__76490;
    wire N__76489;
    wire N__76488;
    wire N__76481;
    wire N__76480;
    wire N__76479;
    wire N__76478;
    wire N__76477;
    wire N__76476;
    wire N__76475;
    wire N__76466;
    wire N__76463;
    wire N__76462;
    wire N__76461;
    wire N__76458;
    wire N__76457;
    wire N__76454;
    wire N__76445;
    wire N__76440;
    wire N__76433;
    wire N__76426;
    wire N__76423;
    wire N__76410;
    wire N__76409;
    wire N__76408;
    wire N__76407;
    wire N__76406;
    wire N__76403;
    wire N__76402;
    wire N__76401;
    wire N__76400;
    wire N__76399;
    wire N__76398;
    wire N__76395;
    wire N__76392;
    wire N__76389;
    wire N__76386;
    wire N__76383;
    wire N__76376;
    wire N__76367;
    wire N__76358;
    wire N__76355;
    wire N__76344;
    wire N__76323;
    wire N__76320;
    wire N__76319;
    wire N__76316;
    wire N__76313;
    wire N__76310;
    wire N__76307;
    wire N__76306;
    wire N__76301;
    wire N__76298;
    wire N__76293;
    wire N__76292;
    wire N__76291;
    wire N__76288;
    wire N__76287;
    wire N__76286;
    wire N__76285;
    wire N__76284;
    wire N__76283;
    wire N__76280;
    wire N__76279;
    wire N__76278;
    wire N__76277;
    wire N__76276;
    wire N__76273;
    wire N__76272;
    wire N__76271;
    wire N__76270;
    wire N__76269;
    wire N__76264;
    wire N__76263;
    wire N__76262;
    wire N__76259;
    wire N__76256;
    wire N__76255;
    wire N__76254;
    wire N__76251;
    wire N__76250;
    wire N__76247;
    wire N__76246;
    wire N__76245;
    wire N__76242;
    wire N__76237;
    wire N__76234;
    wire N__76227;
    wire N__76226;
    wire N__76225;
    wire N__76224;
    wire N__76221;
    wire N__76220;
    wire N__76219;
    wire N__76214;
    wire N__76211;
    wire N__76200;
    wire N__76195;
    wire N__76188;
    wire N__76185;
    wire N__76176;
    wire N__76175;
    wire N__76174;
    wire N__76171;
    wire N__76170;
    wire N__76167;
    wire N__76166;
    wire N__76163;
    wire N__76160;
    wire N__76159;
    wire N__76158;
    wire N__76157;
    wire N__76156;
    wire N__76155;
    wire N__76152;
    wire N__76151;
    wire N__76148;
    wire N__76147;
    wire N__76144;
    wire N__76133;
    wire N__76130;
    wire N__76125;
    wire N__76118;
    wire N__76115;
    wire N__76110;
    wire N__76107;
    wire N__76098;
    wire N__76097;
    wire N__76094;
    wire N__76091;
    wire N__76088;
    wire N__76085;
    wire N__76082;
    wire N__76079;
    wire N__76064;
    wire N__76061;
    wire N__76044;
    wire N__76041;
    wire N__76038;
    wire N__76035;
    wire N__76032;
    wire N__76029;
    wire N__76026;
    wire N__76023;
    wire N__76020;
    wire N__76017;
    wire N__76014;
    wire N__76011;
    wire N__76008;
    wire N__76005;
    wire N__76002;
    wire N__75999;
    wire N__75996;
    wire N__75993;
    wire N__75990;
    wire N__75987;
    wire N__75984;
    wire N__75981;
    wire N__75978;
    wire N__75975;
    wire N__75972;
    wire N__75969;
    wire N__75966;
    wire N__75963;
    wire N__75960;
    wire N__75957;
    wire N__75954;
    wire N__75951;
    wire N__75948;
    wire N__75945;
    wire N__75942;
    wire N__75939;
    wire N__75936;
    wire N__75933;
    wire N__75930;
    wire N__75927;
    wire N__75926;
    wire N__75923;
    wire N__75920;
    wire N__75915;
    wire N__75912;
    wire N__75911;
    wire N__75906;
    wire N__75903;
    wire N__75900;
    wire N__75897;
    wire N__75894;
    wire N__75893;
    wire N__75890;
    wire N__75887;
    wire N__75884;
    wire N__75881;
    wire N__75876;
    wire N__75873;
    wire N__75870;
    wire N__75867;
    wire N__75864;
    wire N__75861;
    wire N__75860;
    wire N__75859;
    wire N__75852;
    wire N__75849;
    wire N__75846;
    wire N__75843;
    wire N__75840;
    wire N__75837;
    wire N__75834;
    wire N__75831;
    wire N__75828;
    wire N__75827;
    wire N__75826;
    wire N__75819;
    wire N__75816;
    wire N__75813;
    wire N__75810;
    wire N__75807;
    wire N__75804;
    wire N__75801;
    wire N__75798;
    wire N__75795;
    wire N__75792;
    wire N__75791;
    wire N__75790;
    wire N__75785;
    wire N__75784;
    wire N__75783;
    wire N__75780;
    wire N__75777;
    wire N__75772;
    wire N__75769;
    wire N__75764;
    wire N__75761;
    wire N__75758;
    wire N__75755;
    wire N__75752;
    wire N__75747;
    wire N__75744;
    wire N__75741;
    wire N__75738;
    wire N__75735;
    wire N__75732;
    wire N__75731;
    wire N__75730;
    wire N__75727;
    wire N__75722;
    wire N__75719;
    wire N__75716;
    wire N__75711;
    wire N__75708;
    wire N__75705;
    wire N__75702;
    wire N__75699;
    wire N__75696;
    wire N__75693;
    wire N__75690;
    wire N__75687;
    wire N__75686;
    wire N__75685;
    wire N__75678;
    wire N__75675;
    wire N__75672;
    wire N__75669;
    wire N__75666;
    wire N__75663;
    wire N__75660;
    wire N__75659;
    wire N__75656;
    wire N__75653;
    wire N__75648;
    wire N__75645;
    wire N__75642;
    wire N__75641;
    wire N__75636;
    wire N__75635;
    wire N__75634;
    wire N__75631;
    wire N__75626;
    wire N__75621;
    wire N__75620;
    wire N__75619;
    wire N__75618;
    wire N__75615;
    wire N__75608;
    wire N__75603;
    wire N__75600;
    wire N__75597;
    wire N__75594;
    wire N__75591;
    wire N__75590;
    wire N__75585;
    wire N__75582;
    wire N__75579;
    wire N__75578;
    wire N__75575;
    wire N__75572;
    wire N__75569;
    wire N__75566;
    wire N__75561;
    wire N__75558;
    wire N__75555;
    wire N__75552;
    wire N__75549;
    wire N__75546;
    wire N__75545;
    wire N__75544;
    wire N__75539;
    wire N__75536;
    wire N__75533;
    wire N__75530;
    wire N__75527;
    wire N__75522;
    wire N__75519;
    wire N__75516;
    wire N__75513;
    wire N__75512;
    wire N__75509;
    wire N__75506;
    wire N__75503;
    wire N__75498;
    wire N__75495;
    wire N__75492;
    wire N__75491;
    wire N__75486;
    wire N__75483;
    wire N__75480;
    wire N__75477;
    wire N__75474;
    wire N__75473;
    wire N__75470;
    wire N__75469;
    wire N__75468;
    wire N__75461;
    wire N__75458;
    wire N__75455;
    wire N__75450;
    wire N__75449;
    wire N__75448;
    wire N__75447;
    wire N__75438;
    wire N__75435;
    wire N__75432;
    wire N__75429;
    wire N__75426;
    wire N__75423;
    wire N__75420;
    wire N__75417;
    wire N__75414;
    wire N__75411;
    wire N__75410;
    wire N__75409;
    wire N__75406;
    wire N__75403;
    wire N__75400;
    wire N__75397;
    wire N__75394;
    wire N__75389;
    wire N__75384;
    wire N__75381;
    wire N__75378;
    wire N__75375;
    wire N__75372;
    wire N__75369;
    wire N__75368;
    wire N__75365;
    wire N__75364;
    wire N__75361;
    wire N__75358;
    wire N__75355;
    wire N__75352;
    wire N__75349;
    wire N__75346;
    wire N__75343;
    wire N__75340;
    wire N__75335;
    wire N__75330;
    wire N__75327;
    wire N__75324;
    wire N__75321;
    wire N__75318;
    wire N__75315;
    wire N__75312;
    wire N__75309;
    wire N__75308;
    wire N__75305;
    wire N__75302;
    wire N__75299;
    wire N__75296;
    wire N__75291;
    wire N__75288;
    wire N__75287;
    wire N__75284;
    wire N__75281;
    wire N__75278;
    wire N__75273;
    wire N__75270;
    wire N__75267;
    wire N__75264;
    wire N__75261;
    wire N__75258;
    wire N__75255;
    wire N__75252;
    wire N__75249;
    wire N__75248;
    wire N__75247;
    wire N__75242;
    wire N__75239;
    wire N__75236;
    wire N__75233;
    wire N__75230;
    wire N__75227;
    wire N__75224;
    wire N__75219;
    wire N__75216;
    wire N__75213;
    wire N__75210;
    wire N__75207;
    wire N__75206;
    wire N__75203;
    wire N__75202;
    wire N__75195;
    wire N__75192;
    wire N__75189;
    wire N__75186;
    wire N__75183;
    wire N__75180;
    wire N__75177;
    wire N__75176;
    wire N__75173;
    wire N__75170;
    wire N__75167;
    wire N__75162;
    wire N__75159;
    wire N__75158;
    wire N__75157;
    wire N__75154;
    wire N__75151;
    wire N__75148;
    wire N__75145;
    wire N__75142;
    wire N__75139;
    wire N__75134;
    wire N__75129;
    wire N__75126;
    wire N__75123;
    wire N__75120;
    wire N__75117;
    wire N__75114;
    wire N__75111;
    wire N__75108;
    wire N__75105;
    wire N__75102;
    wire N__75099;
    wire N__75096;
    wire N__75093;
    wire N__75090;
    wire N__75087;
    wire N__75084;
    wire N__75081;
    wire N__75080;
    wire N__75077;
    wire N__75076;
    wire N__75073;
    wire N__75070;
    wire N__75067;
    wire N__75062;
    wire N__75059;
    wire N__75056;
    wire N__75051;
    wire N__75048;
    wire N__75047;
    wire N__75044;
    wire N__75041;
    wire N__75036;
    wire N__75033;
    wire N__75030;
    wire N__75027;
    wire N__75024;
    wire N__75021;
    wire N__75018;
    wire N__75017;
    wire N__75012;
    wire N__75009;
    wire N__75006;
    wire N__75005;
    wire N__75004;
    wire N__74997;
    wire N__74996;
    wire N__74993;
    wire N__74990;
    wire N__74987;
    wire N__74984;
    wire N__74981;
    wire N__74976;
    wire N__74973;
    wire N__74972;
    wire N__74969;
    wire N__74966;
    wire N__74963;
    wire N__74960;
    wire N__74955;
    wire N__74952;
    wire N__74949;
    wire N__74946;
    wire N__74943;
    wire N__74940;
    wire N__74937;
    wire N__74934;
    wire N__74933;
    wire N__74930;
    wire N__74927;
    wire N__74924;
    wire N__74921;
    wire N__74918;
    wire N__74915;
    wire N__74912;
    wire N__74909;
    wire N__74904;
    wire N__74903;
    wire N__74900;
    wire N__74899;
    wire N__74898;
    wire N__74895;
    wire N__74894;
    wire N__74891;
    wire N__74886;
    wire N__74883;
    wire N__74880;
    wire N__74879;
    wire N__74874;
    wire N__74873;
    wire N__74870;
    wire N__74865;
    wire N__74862;
    wire N__74859;
    wire N__74858;
    wire N__74857;
    wire N__74856;
    wire N__74855;
    wire N__74854;
    wire N__74853;
    wire N__74852;
    wire N__74849;
    wire N__74846;
    wire N__74841;
    wire N__74836;
    wire N__74831;
    wire N__74828;
    wire N__74823;
    wire N__74808;
    wire N__74807;
    wire N__74804;
    wire N__74803;
    wire N__74796;
    wire N__74793;
    wire N__74790;
    wire N__74789;
    wire N__74788;
    wire N__74787;
    wire N__74786;
    wire N__74785;
    wire N__74782;
    wire N__74779;
    wire N__74776;
    wire N__74771;
    wire N__74770;
    wire N__74767;
    wire N__74766;
    wire N__74763;
    wire N__74760;
    wire N__74759;
    wire N__74754;
    wire N__74749;
    wire N__74748;
    wire N__74745;
    wire N__74744;
    wire N__74743;
    wire N__74742;
    wire N__74739;
    wire N__74736;
    wire N__74733;
    wire N__74732;
    wire N__74727;
    wire N__74724;
    wire N__74721;
    wire N__74718;
    wire N__74715;
    wire N__74714;
    wire N__74711;
    wire N__74706;
    wire N__74703;
    wire N__74702;
    wire N__74701;
    wire N__74700;
    wire N__74697;
    wire N__74694;
    wire N__74689;
    wire N__74684;
    wire N__74679;
    wire N__74674;
    wire N__74667;
    wire N__74652;
    wire N__74649;
    wire N__74646;
    wire N__74645;
    wire N__74642;
    wire N__74639;
    wire N__74634;
    wire N__74631;
    wire N__74628;
    wire N__74625;
    wire N__74622;
    wire N__74619;
    wire N__74616;
    wire N__74613;
    wire N__74610;
    wire N__74607;
    wire N__74604;
    wire N__74603;
    wire N__74602;
    wire N__74599;
    wire N__74594;
    wire N__74591;
    wire N__74588;
    wire N__74585;
    wire N__74582;
    wire N__74579;
    wire N__74576;
    wire N__74571;
    wire N__74570;
    wire N__74569;
    wire N__74568;
    wire N__74565;
    wire N__74564;
    wire N__74563;
    wire N__74562;
    wire N__74561;
    wire N__74560;
    wire N__74557;
    wire N__74554;
    wire N__74551;
    wire N__74550;
    wire N__74547;
    wire N__74544;
    wire N__74541;
    wire N__74540;
    wire N__74537;
    wire N__74532;
    wire N__74529;
    wire N__74524;
    wire N__74521;
    wire N__74518;
    wire N__74513;
    wire N__74508;
    wire N__74507;
    wire N__74506;
    wire N__74505;
    wire N__74504;
    wire N__74503;
    wire N__74496;
    wire N__74493;
    wire N__74486;
    wire N__74483;
    wire N__74480;
    wire N__74477;
    wire N__74474;
    wire N__74473;
    wire N__74470;
    wire N__74469;
    wire N__74464;
    wire N__74461;
    wire N__74458;
    wire N__74453;
    wire N__74450;
    wire N__74445;
    wire N__74442;
    wire N__74427;
    wire N__74426;
    wire N__74423;
    wire N__74422;
    wire N__74421;
    wire N__74420;
    wire N__74419;
    wire N__74418;
    wire N__74417;
    wire N__74416;
    wire N__74415;
    wire N__74414;
    wire N__74413;
    wire N__74412;
    wire N__74411;
    wire N__74410;
    wire N__74403;
    wire N__74400;
    wire N__74395;
    wire N__74386;
    wire N__74385;
    wire N__74384;
    wire N__74379;
    wire N__74378;
    wire N__74371;
    wire N__74368;
    wire N__74365;
    wire N__74362;
    wire N__74359;
    wire N__74354;
    wire N__74351;
    wire N__74348;
    wire N__74343;
    wire N__74334;
    wire N__74331;
    wire N__74326;
    wire N__74323;
    wire N__74316;
    wire N__74313;
    wire N__74310;
    wire N__74307;
    wire N__74304;
    wire N__74303;
    wire N__74300;
    wire N__74299;
    wire N__74296;
    wire N__74293;
    wire N__74290;
    wire N__74287;
    wire N__74282;
    wire N__74277;
    wire N__74274;
    wire N__74271;
    wire N__74268;
    wire N__74265;
    wire N__74262;
    wire N__74261;
    wire N__74256;
    wire N__74253;
    wire N__74250;
    wire N__74247;
    wire N__74244;
    wire N__74241;
    wire N__74238;
    wire N__74235;
    wire N__74232;
    wire N__74229;
    wire N__74226;
    wire N__74225;
    wire N__74222;
    wire N__74219;
    wire N__74216;
    wire N__74213;
    wire N__74212;
    wire N__74207;
    wire N__74204;
    wire N__74199;
    wire N__74196;
    wire N__74193;
    wire N__74192;
    wire N__74191;
    wire N__74188;
    wire N__74183;
    wire N__74178;
    wire N__74177;
    wire N__74176;
    wire N__74175;
    wire N__74174;
    wire N__74169;
    wire N__74168;
    wire N__74165;
    wire N__74164;
    wire N__74161;
    wire N__74158;
    wire N__74155;
    wire N__74154;
    wire N__74151;
    wire N__74150;
    wire N__74145;
    wire N__74140;
    wire N__74137;
    wire N__74134;
    wire N__74129;
    wire N__74126;
    wire N__74117;
    wire N__74114;
    wire N__74109;
    wire N__74108;
    wire N__74105;
    wire N__74102;
    wire N__74099;
    wire N__74096;
    wire N__74095;
    wire N__74092;
    wire N__74089;
    wire N__74086;
    wire N__74079;
    wire N__74076;
    wire N__74073;
    wire N__74070;
    wire N__74069;
    wire N__74066;
    wire N__74063;
    wire N__74060;
    wire N__74057;
    wire N__74054;
    wire N__74051;
    wire N__74046;
    wire N__74045;
    wire N__74044;
    wire N__74037;
    wire N__74034;
    wire N__74031;
    wire N__74030;
    wire N__74027;
    wire N__74026;
    wire N__74023;
    wire N__74020;
    wire N__74017;
    wire N__74010;
    wire N__74007;
    wire N__74004;
    wire N__74001;
    wire N__73998;
    wire N__73995;
    wire N__73992;
    wire N__73989;
    wire N__73986;
    wire N__73983;
    wire N__73980;
    wire N__73977;
    wire N__73976;
    wire N__73975;
    wire N__73972;
    wire N__73969;
    wire N__73966;
    wire N__73959;
    wire N__73958;
    wire N__73955;
    wire N__73952;
    wire N__73949;
    wire N__73946;
    wire N__73943;
    wire N__73938;
    wire N__73935;
    wire N__73934;
    wire N__73933;
    wire N__73930;
    wire N__73927;
    wire N__73924;
    wire N__73923;
    wire N__73920;
    wire N__73917;
    wire N__73914;
    wire N__73911;
    wire N__73908;
    wire N__73905;
    wire N__73900;
    wire N__73897;
    wire N__73890;
    wire N__73887;
    wire N__73884;
    wire N__73881;
    wire N__73878;
    wire N__73877;
    wire N__73874;
    wire N__73871;
    wire N__73870;
    wire N__73867;
    wire N__73864;
    wire N__73861;
    wire N__73858;
    wire N__73855;
    wire N__73852;
    wire N__73847;
    wire N__73842;
    wire N__73839;
    wire N__73836;
    wire N__73833;
    wire N__73830;
    wire N__73827;
    wire N__73824;
    wire N__73823;
    wire N__73822;
    wire N__73819;
    wire N__73816;
    wire N__73813;
    wire N__73810;
    wire N__73805;
    wire N__73800;
    wire N__73797;
    wire N__73794;
    wire N__73791;
    wire N__73788;
    wire N__73787;
    wire N__73784;
    wire N__73781;
    wire N__73778;
    wire N__73775;
    wire N__73772;
    wire N__73771;
    wire N__73770;
    wire N__73769;
    wire N__73764;
    wire N__73761;
    wire N__73756;
    wire N__73751;
    wire N__73750;
    wire N__73747;
    wire N__73744;
    wire N__73741;
    wire N__73740;
    wire N__73739;
    wire N__73732;
    wire N__73729;
    wire N__73728;
    wire N__73727;
    wire N__73726;
    wire N__73725;
    wire N__73722;
    wire N__73721;
    wire N__73718;
    wire N__73717;
    wire N__73714;
    wire N__73711;
    wire N__73708;
    wire N__73705;
    wire N__73702;
    wire N__73699;
    wire N__73696;
    wire N__73693;
    wire N__73692;
    wire N__73689;
    wire N__73686;
    wire N__73683;
    wire N__73680;
    wire N__73677;
    wire N__73674;
    wire N__73671;
    wire N__73666;
    wire N__73663;
    wire N__73662;
    wire N__73659;
    wire N__73654;
    wire N__73649;
    wire N__73646;
    wire N__73643;
    wire N__73640;
    wire N__73637;
    wire N__73634;
    wire N__73631;
    wire N__73628;
    wire N__73623;
    wire N__73620;
    wire N__73615;
    wire N__73602;
    wire N__73601;
    wire N__73600;
    wire N__73599;
    wire N__73596;
    wire N__73595;
    wire N__73594;
    wire N__73593;
    wire N__73592;
    wire N__73591;
    wire N__73590;
    wire N__73587;
    wire N__73584;
    wire N__73581;
    wire N__73580;
    wire N__73575;
    wire N__73574;
    wire N__73573;
    wire N__73572;
    wire N__73569;
    wire N__73568;
    wire N__73567;
    wire N__73564;
    wire N__73561;
    wire N__73556;
    wire N__73553;
    wire N__73548;
    wire N__73545;
    wire N__73544;
    wire N__73541;
    wire N__73536;
    wire N__73535;
    wire N__73532;
    wire N__73529;
    wire N__73524;
    wire N__73521;
    wire N__73518;
    wire N__73515;
    wire N__73508;
    wire N__73507;
    wire N__73506;
    wire N__73505;
    wire N__73504;
    wire N__73503;
    wire N__73500;
    wire N__73495;
    wire N__73492;
    wire N__73489;
    wire N__73488;
    wire N__73487;
    wire N__73484;
    wire N__73481;
    wire N__73472;
    wire N__73465;
    wire N__73462;
    wire N__73459;
    wire N__73454;
    wire N__73449;
    wire N__73446;
    wire N__73443;
    wire N__73438;
    wire N__73435;
    wire N__73424;
    wire N__73413;
    wire N__73412;
    wire N__73411;
    wire N__73408;
    wire N__73405;
    wire N__73404;
    wire N__73403;
    wire N__73402;
    wire N__73399;
    wire N__73396;
    wire N__73393;
    wire N__73390;
    wire N__73387;
    wire N__73384;
    wire N__73383;
    wire N__73380;
    wire N__73377;
    wire N__73372;
    wire N__73369;
    wire N__73366;
    wire N__73363;
    wire N__73360;
    wire N__73357;
    wire N__73354;
    wire N__73349;
    wire N__73346;
    wire N__73341;
    wire N__73336;
    wire N__73333;
    wire N__73330;
    wire N__73327;
    wire N__73324;
    wire N__73317;
    wire N__73314;
    wire N__73311;
    wire N__73308;
    wire N__73307;
    wire N__73306;
    wire N__73305;
    wire N__73304;
    wire N__73303;
    wire N__73300;
    wire N__73299;
    wire N__73296;
    wire N__73295;
    wire N__73292;
    wire N__73289;
    wire N__73288;
    wire N__73287;
    wire N__73286;
    wire N__73283;
    wire N__73280;
    wire N__73277;
    wire N__73274;
    wire N__73271;
    wire N__73266;
    wire N__73263;
    wire N__73258;
    wire N__73255;
    wire N__73254;
    wire N__73251;
    wire N__73248;
    wire N__73245;
    wire N__73242;
    wire N__73237;
    wire N__73234;
    wire N__73229;
    wire N__73228;
    wire N__73227;
    wire N__73224;
    wire N__73221;
    wire N__73214;
    wire N__73207;
    wire N__73206;
    wire N__73205;
    wire N__73202;
    wire N__73199;
    wire N__73194;
    wire N__73191;
    wire N__73188;
    wire N__73183;
    wire N__73170;
    wire N__73167;
    wire N__73166;
    wire N__73165;
    wire N__73162;
    wire N__73161;
    wire N__73160;
    wire N__73159;
    wire N__73158;
    wire N__73155;
    wire N__73154;
    wire N__73151;
    wire N__73148;
    wire N__73145;
    wire N__73140;
    wire N__73137;
    wire N__73136;
    wire N__73133;
    wire N__73130;
    wire N__73127;
    wire N__73124;
    wire N__73121;
    wire N__73118;
    wire N__73115;
    wire N__73112;
    wire N__73109;
    wire N__73104;
    wire N__73101;
    wire N__73096;
    wire N__73091;
    wire N__73080;
    wire N__73077;
    wire N__73074;
    wire N__73071;
    wire N__73070;
    wire N__73069;
    wire N__73068;
    wire N__73065;
    wire N__73062;
    wire N__73059;
    wire N__73056;
    wire N__73055;
    wire N__73054;
    wire N__73053;
    wire N__73052;
    wire N__73051;
    wire N__73046;
    wire N__73043;
    wire N__73040;
    wire N__73037;
    wire N__73034;
    wire N__73031;
    wire N__73026;
    wire N__73023;
    wire N__73012;
    wire N__73009;
    wire N__73004;
    wire N__72999;
    wire N__72998;
    wire N__72995;
    wire N__72994;
    wire N__72993;
    wire N__72992;
    wire N__72991;
    wire N__72990;
    wire N__72989;
    wire N__72988;
    wire N__72985;
    wire N__72984;
    wire N__72983;
    wire N__72982;
    wire N__72981;
    wire N__72978;
    wire N__72973;
    wire N__72972;
    wire N__72971;
    wire N__72968;
    wire N__72965;
    wire N__72960;
    wire N__72959;
    wire N__72958;
    wire N__72951;
    wire N__72948;
    wire N__72943;
    wire N__72940;
    wire N__72937;
    wire N__72934;
    wire N__72931;
    wire N__72928;
    wire N__72923;
    wire N__72922;
    wire N__72919;
    wire N__72918;
    wire N__72915;
    wire N__72912;
    wire N__72909;
    wire N__72908;
    wire N__72907;
    wire N__72904;
    wire N__72901;
    wire N__72898;
    wire N__72895;
    wire N__72888;
    wire N__72887;
    wire N__72886;
    wire N__72885;
    wire N__72884;
    wire N__72883;
    wire N__72880;
    wire N__72877;
    wire N__72872;
    wire N__72867;
    wire N__72864;
    wire N__72861;
    wire N__72854;
    wire N__72849;
    wire N__72840;
    wire N__72835;
    wire N__72830;
    wire N__72825;
    wire N__72810;
    wire N__72807;
    wire N__72804;
    wire N__72801;
    wire N__72798;
    wire N__72797;
    wire N__72794;
    wire N__72791;
    wire N__72790;
    wire N__72789;
    wire N__72788;
    wire N__72787;
    wire N__72786;
    wire N__72785;
    wire N__72782;
    wire N__72779;
    wire N__72776;
    wire N__72773;
    wire N__72770;
    wire N__72769;
    wire N__72766;
    wire N__72763;
    wire N__72760;
    wire N__72757;
    wire N__72754;
    wire N__72747;
    wire N__72744;
    wire N__72737;
    wire N__72734;
    wire N__72731;
    wire N__72726;
    wire N__72723;
    wire N__72714;
    wire N__72711;
    wire N__72708;
    wire N__72707;
    wire N__72704;
    wire N__72703;
    wire N__72700;
    wire N__72699;
    wire N__72698;
    wire N__72697;
    wire N__72696;
    wire N__72695;
    wire N__72692;
    wire N__72689;
    wire N__72686;
    wire N__72683;
    wire N__72680;
    wire N__72679;
    wire N__72678;
    wire N__72677;
    wire N__72676;
    wire N__72675;
    wire N__72668;
    wire N__72665;
    wire N__72664;
    wire N__72663;
    wire N__72660;
    wire N__72657;
    wire N__72652;
    wire N__72649;
    wire N__72644;
    wire N__72639;
    wire N__72634;
    wire N__72631;
    wire N__72628;
    wire N__72621;
    wire N__72616;
    wire N__72613;
    wire N__72608;
    wire N__72605;
    wire N__72598;
    wire N__72595;
    wire N__72588;
    wire N__72585;
    wire N__72584;
    wire N__72583;
    wire N__72582;
    wire N__72581;
    wire N__72580;
    wire N__72577;
    wire N__72574;
    wire N__72573;
    wire N__72570;
    wire N__72569;
    wire N__72566;
    wire N__72563;
    wire N__72560;
    wire N__72557;
    wire N__72554;
    wire N__72551;
    wire N__72548;
    wire N__72545;
    wire N__72538;
    wire N__72535;
    wire N__72526;
    wire N__72523;
    wire N__72516;
    wire N__72513;
    wire N__72512;
    wire N__72509;
    wire N__72506;
    wire N__72505;
    wire N__72504;
    wire N__72503;
    wire N__72502;
    wire N__72501;
    wire N__72498;
    wire N__72495;
    wire N__72492;
    wire N__72489;
    wire N__72488;
    wire N__72485;
    wire N__72482;
    wire N__72479;
    wire N__72476;
    wire N__72473;
    wire N__72468;
    wire N__72465;
    wire N__72458;
    wire N__72455;
    wire N__72452;
    wire N__72447;
    wire N__72444;
    wire N__72435;
    wire N__72432;
    wire N__72431;
    wire N__72430;
    wire N__72427;
    wire N__72426;
    wire N__72425;
    wire N__72422;
    wire N__72421;
    wire N__72418;
    wire N__72415;
    wire N__72412;
    wire N__72411;
    wire N__72410;
    wire N__72407;
    wire N__72404;
    wire N__72399;
    wire N__72396;
    wire N__72393;
    wire N__72390;
    wire N__72387;
    wire N__72384;
    wire N__72381;
    wire N__72378;
    wire N__72375;
    wire N__72370;
    wire N__72367;
    wire N__72356;
    wire N__72351;
    wire N__72348;
    wire N__72347;
    wire N__72346;
    wire N__72345;
    wire N__72344;
    wire N__72341;
    wire N__72338;
    wire N__72337;
    wire N__72336;
    wire N__72335;
    wire N__72332;
    wire N__72329;
    wire N__72326;
    wire N__72321;
    wire N__72318;
    wire N__72315;
    wire N__72312;
    wire N__72307;
    wire N__72304;
    wire N__72301;
    wire N__72294;
    wire N__72289;
    wire N__72284;
    wire N__72279;
    wire N__72276;
    wire N__72275;
    wire N__72274;
    wire N__72273;
    wire N__72272;
    wire N__72271;
    wire N__72270;
    wire N__72269;
    wire N__72266;
    wire N__72261;
    wire N__72260;
    wire N__72257;
    wire N__72254;
    wire N__72253;
    wire N__72250;
    wire N__72247;
    wire N__72246;
    wire N__72245;
    wire N__72244;
    wire N__72241;
    wire N__72238;
    wire N__72235;
    wire N__72230;
    wire N__72227;
    wire N__72222;
    wire N__72221;
    wire N__72220;
    wire N__72219;
    wire N__72218;
    wire N__72215;
    wire N__72212;
    wire N__72211;
    wire N__72210;
    wire N__72209;
    wire N__72204;
    wire N__72201;
    wire N__72198;
    wire N__72193;
    wire N__72188;
    wire N__72187;
    wire N__72184;
    wire N__72181;
    wire N__72180;
    wire N__72179;
    wire N__72178;
    wire N__72175;
    wire N__72172;
    wire N__72169;
    wire N__72166;
    wire N__72163;
    wire N__72160;
    wire N__72157;
    wire N__72152;
    wire N__72145;
    wire N__72140;
    wire N__72137;
    wire N__72134;
    wire N__72127;
    wire N__72102;
    wire N__72099;
    wire N__72096;
    wire N__72093;
    wire N__72092;
    wire N__72089;
    wire N__72086;
    wire N__72081;
    wire N__72078;
    wire N__72075;
    wire N__72072;
    wire N__72071;
    wire N__72070;
    wire N__72067;
    wire N__72060;
    wire N__72057;
    wire N__72056;
    wire N__72055;
    wire N__72054;
    wire N__72051;
    wire N__72044;
    wire N__72043;
    wire N__72042;
    wire N__72037;
    wire N__72032;
    wire N__72029;
    wire N__72026;
    wire N__72025;
    wire N__72022;
    wire N__72019;
    wire N__72016;
    wire N__72013;
    wire N__72008;
    wire N__72003;
    wire N__72000;
    wire N__71999;
    wire N__71996;
    wire N__71993;
    wire N__71990;
    wire N__71985;
    wire N__71984;
    wire N__71983;
    wire N__71980;
    wire N__71979;
    wire N__71978;
    wire N__71977;
    wire N__71976;
    wire N__71973;
    wire N__71972;
    wire N__71971;
    wire N__71970;
    wire N__71961;
    wire N__71960;
    wire N__71959;
    wire N__71958;
    wire N__71957;
    wire N__71956;
    wire N__71947;
    wire N__71946;
    wire N__71943;
    wire N__71940;
    wire N__71939;
    wire N__71936;
    wire N__71927;
    wire N__71924;
    wire N__71921;
    wire N__71912;
    wire N__71911;
    wire N__71908;
    wire N__71905;
    wire N__71902;
    wire N__71897;
    wire N__71894;
    wire N__71893;
    wire N__71888;
    wire N__71885;
    wire N__71882;
    wire N__71877;
    wire N__71876;
    wire N__71875;
    wire N__71872;
    wire N__71867;
    wire N__71864;
    wire N__71859;
    wire N__71856;
    wire N__71851;
    wire N__71844;
    wire N__71843;
    wire N__71842;
    wire N__71839;
    wire N__71838;
    wire N__71837;
    wire N__71834;
    wire N__71833;
    wire N__71830;
    wire N__71827;
    wire N__71824;
    wire N__71821;
    wire N__71818;
    wire N__71813;
    wire N__71810;
    wire N__71805;
    wire N__71802;
    wire N__71799;
    wire N__71798;
    wire N__71791;
    wire N__71788;
    wire N__71785;
    wire N__71782;
    wire N__71777;
    wire N__71774;
    wire N__71771;
    wire N__71766;
    wire N__71765;
    wire N__71762;
    wire N__71761;
    wire N__71760;
    wire N__71757;
    wire N__71756;
    wire N__71755;
    wire N__71754;
    wire N__71753;
    wire N__71752;
    wire N__71751;
    wire N__71742;
    wire N__71733;
    wire N__71730;
    wire N__71729;
    wire N__71728;
    wire N__71725;
    wire N__71724;
    wire N__71721;
    wire N__71718;
    wire N__71709;
    wire N__71706;
    wire N__71699;
    wire N__71694;
    wire N__71693;
    wire N__71688;
    wire N__71685;
    wire N__71682;
    wire N__71679;
    wire N__71676;
    wire N__71675;
    wire N__71672;
    wire N__71671;
    wire N__71670;
    wire N__71669;
    wire N__71668;
    wire N__71665;
    wire N__71662;
    wire N__71661;
    wire N__71660;
    wire N__71659;
    wire N__71654;
    wire N__71651;
    wire N__71648;
    wire N__71645;
    wire N__71642;
    wire N__71637;
    wire N__71634;
    wire N__71631;
    wire N__71628;
    wire N__71625;
    wire N__71622;
    wire N__71619;
    wire N__71610;
    wire N__71605;
    wire N__71602;
    wire N__71599;
    wire N__71592;
    wire N__71589;
    wire N__71586;
    wire N__71585;
    wire N__71584;
    wire N__71583;
    wire N__71582;
    wire N__71579;
    wire N__71578;
    wire N__71577;
    wire N__71574;
    wire N__71571;
    wire N__71566;
    wire N__71563;
    wire N__71560;
    wire N__71559;
    wire N__71558;
    wire N__71557;
    wire N__71554;
    wire N__71553;
    wire N__71552;
    wire N__71549;
    wire N__71546;
    wire N__71543;
    wire N__71542;
    wire N__71541;
    wire N__71538;
    wire N__71535;
    wire N__71532;
    wire N__71527;
    wire N__71526;
    wire N__71525;
    wire N__71518;
    wire N__71511;
    wire N__71508;
    wire N__71505;
    wire N__71496;
    wire N__71491;
    wire N__71488;
    wire N__71485;
    wire N__71476;
    wire N__71469;
    wire N__71468;
    wire N__71467;
    wire N__71464;
    wire N__71463;
    wire N__71462;
    wire N__71461;
    wire N__71458;
    wire N__71455;
    wire N__71454;
    wire N__71453;
    wire N__71452;
    wire N__71451;
    wire N__71450;
    wire N__71449;
    wire N__71448;
    wire N__71447;
    wire N__71444;
    wire N__71437;
    wire N__71434;
    wire N__71431;
    wire N__71428;
    wire N__71423;
    wire N__71420;
    wire N__71417;
    wire N__71412;
    wire N__71409;
    wire N__71404;
    wire N__71399;
    wire N__71398;
    wire N__71397;
    wire N__71394;
    wire N__71389;
    wire N__71384;
    wire N__71381;
    wire N__71376;
    wire N__71371;
    wire N__71368;
    wire N__71365;
    wire N__71360;
    wire N__71357;
    wire N__71354;
    wire N__71349;
    wire N__71346;
    wire N__71337;
    wire N__71334;
    wire N__71331;
    wire N__71330;
    wire N__71327;
    wire N__71326;
    wire N__71323;
    wire N__71320;
    wire N__71317;
    wire N__71314;
    wire N__71311;
    wire N__71310;
    wire N__71309;
    wire N__71308;
    wire N__71305;
    wire N__71304;
    wire N__71303;
    wire N__71302;
    wire N__71299;
    wire N__71296;
    wire N__71291;
    wire N__71288;
    wire N__71285;
    wire N__71282;
    wire N__71277;
    wire N__71274;
    wire N__71271;
    wire N__71268;
    wire N__71253;
    wire N__71250;
    wire N__71247;
    wire N__71244;
    wire N__71241;
    wire N__71240;
    wire N__71237;
    wire N__71236;
    wire N__71233;
    wire N__71230;
    wire N__71227;
    wire N__71224;
    wire N__71223;
    wire N__71220;
    wire N__71217;
    wire N__71216;
    wire N__71213;
    wire N__71212;
    wire N__71209;
    wire N__71206;
    wire N__71203;
    wire N__71200;
    wire N__71199;
    wire N__71198;
    wire N__71195;
    wire N__71192;
    wire N__71189;
    wire N__71184;
    wire N__71177;
    wire N__71166;
    wire N__71165;
    wire N__71162;
    wire N__71161;
    wire N__71160;
    wire N__71157;
    wire N__71156;
    wire N__71155;
    wire N__71154;
    wire N__71151;
    wire N__71150;
    wire N__71149;
    wire N__71148;
    wire N__71147;
    wire N__71146;
    wire N__71143;
    wire N__71140;
    wire N__71137;
    wire N__71134;
    wire N__71131;
    wire N__71128;
    wire N__71127;
    wire N__71124;
    wire N__71121;
    wire N__71118;
    wire N__71117;
    wire N__71116;
    wire N__71113;
    wire N__71110;
    wire N__71109;
    wire N__71104;
    wire N__71101;
    wire N__71098;
    wire N__71093;
    wire N__71090;
    wire N__71089;
    wire N__71086;
    wire N__71083;
    wire N__71080;
    wire N__71077;
    wire N__71076;
    wire N__71071;
    wire N__71068;
    wire N__71065;
    wire N__71064;
    wire N__71061;
    wire N__71060;
    wire N__71059;
    wire N__71056;
    wire N__71047;
    wire N__71044;
    wire N__71035;
    wire N__71032;
    wire N__71029;
    wire N__71024;
    wire N__71019;
    wire N__71014;
    wire N__71009;
    wire N__70992;
    wire N__70989;
    wire N__70988;
    wire N__70985;
    wire N__70984;
    wire N__70981;
    wire N__70978;
    wire N__70977;
    wire N__70974;
    wire N__70971;
    wire N__70968;
    wire N__70967;
    wire N__70966;
    wire N__70963;
    wire N__70962;
    wire N__70961;
    wire N__70958;
    wire N__70955;
    wire N__70952;
    wire N__70949;
    wire N__70946;
    wire N__70943;
    wire N__70938;
    wire N__70935;
    wire N__70920;
    wire N__70919;
    wire N__70916;
    wire N__70915;
    wire N__70914;
    wire N__70911;
    wire N__70908;
    wire N__70907;
    wire N__70904;
    wire N__70901;
    wire N__70898;
    wire N__70895;
    wire N__70894;
    wire N__70893;
    wire N__70892;
    wire N__70889;
    wire N__70886;
    wire N__70883;
    wire N__70880;
    wire N__70877;
    wire N__70874;
    wire N__70869;
    wire N__70866;
    wire N__70863;
    wire N__70858;
    wire N__70855;
    wire N__70842;
    wire N__70839;
    wire N__70836;
    wire N__70833;
    wire N__70832;
    wire N__70829;
    wire N__70826;
    wire N__70825;
    wire N__70824;
    wire N__70823;
    wire N__70818;
    wire N__70815;
    wire N__70810;
    wire N__70809;
    wire N__70808;
    wire N__70807;
    wire N__70804;
    wire N__70801;
    wire N__70798;
    wire N__70795;
    wire N__70792;
    wire N__70789;
    wire N__70782;
    wire N__70773;
    wire N__70770;
    wire N__70769;
    wire N__70766;
    wire N__70763;
    wire N__70758;
    wire N__70755;
    wire N__70752;
    wire N__70749;
    wire N__70748;
    wire N__70747;
    wire N__70746;
    wire N__70743;
    wire N__70742;
    wire N__70741;
    wire N__70738;
    wire N__70737;
    wire N__70734;
    wire N__70733;
    wire N__70732;
    wire N__70731;
    wire N__70728;
    wire N__70725;
    wire N__70722;
    wire N__70719;
    wire N__70716;
    wire N__70713;
    wire N__70710;
    wire N__70707;
    wire N__70706;
    wire N__70705;
    wire N__70704;
    wire N__70703;
    wire N__70702;
    wire N__70699;
    wire N__70698;
    wire N__70697;
    wire N__70696;
    wire N__70693;
    wire N__70690;
    wire N__70687;
    wire N__70684;
    wire N__70673;
    wire N__70670;
    wire N__70667;
    wire N__70664;
    wire N__70661;
    wire N__70660;
    wire N__70657;
    wire N__70656;
    wire N__70651;
    wire N__70648;
    wire N__70647;
    wire N__70646;
    wire N__70645;
    wire N__70644;
    wire N__70643;
    wire N__70640;
    wire N__70639;
    wire N__70638;
    wire N__70629;
    wire N__70626;
    wire N__70617;
    wire N__70616;
    wire N__70615;
    wire N__70614;
    wire N__70611;
    wire N__70608;
    wire N__70605;
    wire N__70600;
    wire N__70595;
    wire N__70586;
    wire N__70583;
    wire N__70580;
    wire N__70577;
    wire N__70572;
    wire N__70569;
    wire N__70566;
    wire N__70563;
    wire N__70556;
    wire N__70551;
    wire N__70530;
    wire N__70529;
    wire N__70528;
    wire N__70527;
    wire N__70526;
    wire N__70525;
    wire N__70522;
    wire N__70521;
    wire N__70518;
    wire N__70517;
    wire N__70516;
    wire N__70515;
    wire N__70514;
    wire N__70513;
    wire N__70512;
    wire N__70511;
    wire N__70510;
    wire N__70509;
    wire N__70506;
    wire N__70503;
    wire N__70502;
    wire N__70501;
    wire N__70500;
    wire N__70499;
    wire N__70498;
    wire N__70497;
    wire N__70496;
    wire N__70495;
    wire N__70494;
    wire N__70493;
    wire N__70492;
    wire N__70491;
    wire N__70486;
    wire N__70481;
    wire N__70478;
    wire N__70475;
    wire N__70472;
    wire N__70471;
    wire N__70470;
    wire N__70469;
    wire N__70468;
    wire N__70467;
    wire N__70466;
    wire N__70463;
    wire N__70460;
    wire N__70459;
    wire N__70458;
    wire N__70457;
    wire N__70454;
    wire N__70453;
    wire N__70446;
    wire N__70443;
    wire N__70438;
    wire N__70435;
    wire N__70434;
    wire N__70433;
    wire N__70432;
    wire N__70431;
    wire N__70428;
    wire N__70427;
    wire N__70422;
    wire N__70417;
    wire N__70416;
    wire N__70415;
    wire N__70412;
    wire N__70411;
    wire N__70410;
    wire N__70409;
    wire N__70408;
    wire N__70407;
    wire N__70404;
    wire N__70403;
    wire N__70400;
    wire N__70393;
    wire N__70384;
    wire N__70381;
    wire N__70380;
    wire N__70379;
    wire N__70376;
    wire N__70371;
    wire N__70366;
    wire N__70361;
    wire N__70360;
    wire N__70359;
    wire N__70358;
    wire N__70355;
    wire N__70352;
    wire N__70347;
    wire N__70344;
    wire N__70341;
    wire N__70332;
    wire N__70327;
    wire N__70318;
    wire N__70313;
    wire N__70312;
    wire N__70309;
    wire N__70308;
    wire N__70305;
    wire N__70300;
    wire N__70297;
    wire N__70296;
    wire N__70295;
    wire N__70292;
    wire N__70283;
    wire N__70280;
    wire N__70273;
    wire N__70268;
    wire N__70265;
    wire N__70260;
    wire N__70257;
    wire N__70254;
    wire N__70253;
    wire N__70252;
    wire N__70251;
    wire N__70250;
    wire N__70247;
    wire N__70246;
    wire N__70245;
    wire N__70244;
    wire N__70241;
    wire N__70236;
    wire N__70233;
    wire N__70228;
    wire N__70219;
    wire N__70216;
    wire N__70209;
    wire N__70206;
    wire N__70199;
    wire N__70188;
    wire N__70179;
    wire N__70174;
    wire N__70169;
    wire N__70166;
    wire N__70161;
    wire N__70158;
    wire N__70147;
    wire N__70142;
    wire N__70137;
    wire N__70130;
    wire N__70125;
    wire N__70110;
    wire N__70107;
    wire N__70104;
    wire N__70101;
    wire N__70100;
    wire N__70099;
    wire N__70096;
    wire N__70093;
    wire N__70092;
    wire N__70091;
    wire N__70090;
    wire N__70089;
    wire N__70088;
    wire N__70087;
    wire N__70084;
    wire N__70083;
    wire N__70082;
    wire N__70081;
    wire N__70080;
    wire N__70079;
    wire N__70074;
    wire N__70069;
    wire N__70060;
    wire N__70057;
    wire N__70054;
    wire N__70051;
    wire N__70046;
    wire N__70043;
    wire N__70042;
    wire N__70041;
    wire N__70040;
    wire N__70039;
    wire N__70038;
    wire N__70035;
    wire N__70030;
    wire N__70019;
    wire N__70014;
    wire N__70013;
    wire N__70012;
    wire N__70009;
    wire N__70004;
    wire N__69999;
    wire N__69994;
    wire N__69989;
    wire N__69978;
    wire N__69977;
    wire N__69974;
    wire N__69971;
    wire N__69970;
    wire N__69969;
    wire N__69966;
    wire N__69961;
    wire N__69958;
    wire N__69957;
    wire N__69956;
    wire N__69955;
    wire N__69954;
    wire N__69953;
    wire N__69952;
    wire N__69951;
    wire N__69950;
    wire N__69949;
    wire N__69946;
    wire N__69943;
    wire N__69940;
    wire N__69937;
    wire N__69934;
    wire N__69933;
    wire N__69930;
    wire N__69929;
    wire N__69928;
    wire N__69925;
    wire N__69922;
    wire N__69919;
    wire N__69916;
    wire N__69915;
    wire N__69914;
    wire N__69909;
    wire N__69898;
    wire N__69893;
    wire N__69890;
    wire N__69887;
    wire N__69886;
    wire N__69883;
    wire N__69880;
    wire N__69877;
    wire N__69874;
    wire N__69873;
    wire N__69872;
    wire N__69869;
    wire N__69868;
    wire N__69867;
    wire N__69866;
    wire N__69865;
    wire N__69862;
    wire N__69861;
    wire N__69854;
    wire N__69853;
    wire N__69852;
    wire N__69851;
    wire N__69848;
    wire N__69847;
    wire N__69844;
    wire N__69841;
    wire N__69832;
    wire N__69829;
    wire N__69826;
    wire N__69823;
    wire N__69820;
    wire N__69817;
    wire N__69816;
    wire N__69813;
    wire N__69810;
    wire N__69805;
    wire N__69802;
    wire N__69799;
    wire N__69796;
    wire N__69793;
    wire N__69790;
    wire N__69787;
    wire N__69786;
    wire N__69781;
    wire N__69778;
    wire N__69775;
    wire N__69770;
    wire N__69767;
    wire N__69766;
    wire N__69765;
    wire N__69762;
    wire N__69759;
    wire N__69748;
    wire N__69745;
    wire N__69740;
    wire N__69737;
    wire N__69734;
    wire N__69723;
    wire N__69718;
    wire N__69711;
    wire N__69696;
    wire N__69695;
    wire N__69692;
    wire N__69689;
    wire N__69688;
    wire N__69683;
    wire N__69682;
    wire N__69681;
    wire N__69680;
    wire N__69679;
    wire N__69676;
    wire N__69673;
    wire N__69668;
    wire N__69667;
    wire N__69666;
    wire N__69663;
    wire N__69662;
    wire N__69661;
    wire N__69660;
    wire N__69659;
    wire N__69658;
    wire N__69657;
    wire N__69656;
    wire N__69655;
    wire N__69654;
    wire N__69653;
    wire N__69652;
    wire N__69651;
    wire N__69648;
    wire N__69645;
    wire N__69640;
    wire N__69637;
    wire N__69636;
    wire N__69635;
    wire N__69634;
    wire N__69633;
    wire N__69632;
    wire N__69627;
    wire N__69626;
    wire N__69625;
    wire N__69620;
    wire N__69617;
    wire N__69614;
    wire N__69611;
    wire N__69608;
    wire N__69603;
    wire N__69602;
    wire N__69601;
    wire N__69600;
    wire N__69599;
    wire N__69596;
    wire N__69591;
    wire N__69588;
    wire N__69587;
    wire N__69586;
    wire N__69577;
    wire N__69576;
    wire N__69573;
    wire N__69570;
    wire N__69567;
    wire N__69566;
    wire N__69565;
    wire N__69560;
    wire N__69557;
    wire N__69554;
    wire N__69551;
    wire N__69550;
    wire N__69545;
    wire N__69538;
    wire N__69537;
    wire N__69536;
    wire N__69535;
    wire N__69534;
    wire N__69531;
    wire N__69528;
    wire N__69523;
    wire N__69520;
    wire N__69513;
    wire N__69508;
    wire N__69505;
    wire N__69502;
    wire N__69501;
    wire N__69500;
    wire N__69497;
    wire N__69494;
    wire N__69491;
    wire N__69486;
    wire N__69481;
    wire N__69480;
    wire N__69477;
    wire N__69474;
    wire N__69471;
    wire N__69466;
    wire N__69459;
    wire N__69456;
    wire N__69453;
    wire N__69450;
    wire N__69447;
    wire N__69444;
    wire N__69435;
    wire N__69430;
    wire N__69425;
    wire N__69418;
    wire N__69415;
    wire N__69410;
    wire N__69403;
    wire N__69400;
    wire N__69395;
    wire N__69388;
    wire N__69379;
    wire N__69374;
    wire N__69367;
    wire N__69364;
    wire N__69357;
    wire N__69354;
    wire N__69351;
    wire N__69348;
    wire N__69345;
    wire N__69342;
    wire N__69339;
    wire N__69336;
    wire N__69333;
    wire N__69330;
    wire N__69327;
    wire N__69324;
    wire N__69323;
    wire N__69322;
    wire N__69321;
    wire N__69318;
    wire N__69317;
    wire N__69316;
    wire N__69313;
    wire N__69310;
    wire N__69307;
    wire N__69306;
    wire N__69305;
    wire N__69304;
    wire N__69303;
    wire N__69300;
    wire N__69299;
    wire N__69296;
    wire N__69293;
    wire N__69290;
    wire N__69287;
    wire N__69284;
    wire N__69281;
    wire N__69278;
    wire N__69275;
    wire N__69272;
    wire N__69269;
    wire N__69266;
    wire N__69261;
    wire N__69260;
    wire N__69257;
    wire N__69254;
    wire N__69249;
    wire N__69246;
    wire N__69243;
    wire N__69236;
    wire N__69233;
    wire N__69230;
    wire N__69225;
    wire N__69222;
    wire N__69219;
    wire N__69216;
    wire N__69213;
    wire N__69210;
    wire N__69207;
    wire N__69202;
    wire N__69199;
    wire N__69194;
    wire N__69191;
    wire N__69188;
    wire N__69185;
    wire N__69182;
    wire N__69177;
    wire N__69172;
    wire N__69165;
    wire N__69164;
    wire N__69163;
    wire N__69162;
    wire N__69159;
    wire N__69158;
    wire N__69157;
    wire N__69156;
    wire N__69153;
    wire N__69150;
    wire N__69147;
    wire N__69146;
    wire N__69143;
    wire N__69142;
    wire N__69137;
    wire N__69134;
    wire N__69133;
    wire N__69130;
    wire N__69125;
    wire N__69122;
    wire N__69119;
    wire N__69116;
    wire N__69111;
    wire N__69108;
    wire N__69105;
    wire N__69102;
    wire N__69099;
    wire N__69094;
    wire N__69091;
    wire N__69078;
    wire N__69075;
    wire N__69072;
    wire N__69069;
    wire N__69066;
    wire N__69063;
    wire N__69060;
    wire N__69057;
    wire N__69054;
    wire N__69051;
    wire N__69048;
    wire N__69045;
    wire N__69042;
    wire N__69041;
    wire N__69040;
    wire N__69039;
    wire N__69038;
    wire N__69037;
    wire N__69036;
    wire N__69033;
    wire N__69032;
    wire N__69029;
    wire N__69020;
    wire N__69017;
    wire N__69016;
    wire N__69013;
    wire N__69010;
    wire N__69007;
    wire N__69004;
    wire N__68999;
    wire N__68996;
    wire N__68991;
    wire N__68988;
    wire N__68979;
    wire N__68976;
    wire N__68973;
    wire N__68970;
    wire N__68967;
    wire N__68964;
    wire N__68961;
    wire N__68958;
    wire N__68955;
    wire N__68952;
    wire N__68949;
    wire N__68946;
    wire N__68943;
    wire N__68942;
    wire N__68941;
    wire N__68940;
    wire N__68937;
    wire N__68930;
    wire N__68925;
    wire N__68922;
    wire N__68919;
    wire N__68916;
    wire N__68913;
    wire N__68910;
    wire N__68909;
    wire N__68908;
    wire N__68905;
    wire N__68900;
    wire N__68895;
    wire N__68892;
    wire N__68889;
    wire N__68886;
    wire N__68883;
    wire N__68880;
    wire N__68877;
    wire N__68876;
    wire N__68873;
    wire N__68870;
    wire N__68865;
    wire N__68864;
    wire N__68861;
    wire N__68860;
    wire N__68855;
    wire N__68852;
    wire N__68849;
    wire N__68844;
    wire N__68841;
    wire N__68838;
    wire N__68835;
    wire N__68832;
    wire N__68829;
    wire N__68826;
    wire N__68823;
    wire N__68820;
    wire N__68817;
    wire N__68814;
    wire N__68811;
    wire N__68808;
    wire N__68805;
    wire N__68802;
    wire N__68799;
    wire N__68796;
    wire N__68793;
    wire N__68790;
    wire N__68787;
    wire N__68784;
    wire N__68781;
    wire N__68778;
    wire N__68775;
    wire N__68772;
    wire N__68769;
    wire N__68766;
    wire N__68763;
    wire N__68760;
    wire N__68757;
    wire N__68754;
    wire N__68751;
    wire N__68748;
    wire N__68745;
    wire N__68742;
    wire N__68739;
    wire N__68736;
    wire N__68733;
    wire N__68730;
    wire N__68727;
    wire N__68724;
    wire N__68721;
    wire N__68718;
    wire N__68715;
    wire N__68712;
    wire N__68709;
    wire N__68706;
    wire N__68703;
    wire N__68700;
    wire N__68697;
    wire N__68694;
    wire N__68693;
    wire N__68692;
    wire N__68689;
    wire N__68686;
    wire N__68683;
    wire N__68678;
    wire N__68673;
    wire N__68670;
    wire N__68667;
    wire N__68666;
    wire N__68663;
    wire N__68660;
    wire N__68655;
    wire N__68654;
    wire N__68651;
    wire N__68648;
    wire N__68643;
    wire N__68640;
    wire N__68639;
    wire N__68638;
    wire N__68637;
    wire N__68636;
    wire N__68633;
    wire N__68632;
    wire N__68627;
    wire N__68622;
    wire N__68619;
    wire N__68616;
    wire N__68613;
    wire N__68610;
    wire N__68605;
    wire N__68600;
    wire N__68597;
    wire N__68592;
    wire N__68591;
    wire N__68586;
    wire N__68583;
    wire N__68582;
    wire N__68577;
    wire N__68574;
    wire N__68573;
    wire N__68570;
    wire N__68565;
    wire N__68564;
    wire N__68563;
    wire N__68562;
    wire N__68561;
    wire N__68558;
    wire N__68555;
    wire N__68552;
    wire N__68547;
    wire N__68544;
    wire N__68543;
    wire N__68542;
    wire N__68539;
    wire N__68536;
    wire N__68533;
    wire N__68530;
    wire N__68525;
    wire N__68522;
    wire N__68519;
    wire N__68516;
    wire N__68511;
    wire N__68508;
    wire N__68505;
    wire N__68502;
    wire N__68499;
    wire N__68490;
    wire N__68489;
    wire N__68484;
    wire N__68481;
    wire N__68478;
    wire N__68475;
    wire N__68472;
    wire N__68471;
    wire N__68468;
    wire N__68465;
    wire N__68460;
    wire N__68457;
    wire N__68454;
    wire N__68451;
    wire N__68450;
    wire N__68447;
    wire N__68444;
    wire N__68441;
    wire N__68438;
    wire N__68433;
    wire N__68430;
    wire N__68427;
    wire N__68424;
    wire N__68421;
    wire N__68418;
    wire N__68415;
    wire N__68414;
    wire N__68411;
    wire N__68408;
    wire N__68405;
    wire N__68402;
    wire N__68399;
    wire N__68394;
    wire N__68391;
    wire N__68390;
    wire N__68387;
    wire N__68384;
    wire N__68381;
    wire N__68376;
    wire N__68373;
    wire N__68370;
    wire N__68367;
    wire N__68364;
    wire N__68361;
    wire N__68358;
    wire N__68355;
    wire N__68352;
    wire N__68349;
    wire N__68346;
    wire N__68343;
    wire N__68342;
    wire N__68339;
    wire N__68336;
    wire N__68333;
    wire N__68330;
    wire N__68327;
    wire N__68322;
    wire N__68319;
    wire N__68316;
    wire N__68315;
    wire N__68314;
    wire N__68309;
    wire N__68306;
    wire N__68303;
    wire N__68300;
    wire N__68297;
    wire N__68292;
    wire N__68289;
    wire N__68288;
    wire N__68285;
    wire N__68282;
    wire N__68277;
    wire N__68276;
    wire N__68273;
    wire N__68270;
    wire N__68269;
    wire N__68264;
    wire N__68261;
    wire N__68256;
    wire N__68253;
    wire N__68250;
    wire N__68247;
    wire N__68246;
    wire N__68243;
    wire N__68240;
    wire N__68235;
    wire N__68232;
    wire N__68231;
    wire N__68228;
    wire N__68225;
    wire N__68220;
    wire N__68219;
    wire N__68216;
    wire N__68213;
    wire N__68212;
    wire N__68209;
    wire N__68206;
    wire N__68203;
    wire N__68200;
    wire N__68193;
    wire N__68190;
    wire N__68189;
    wire N__68186;
    wire N__68183;
    wire N__68178;
    wire N__68175;
    wire N__68172;
    wire N__68169;
    wire N__68166;
    wire N__68165;
    wire N__68162;
    wire N__68159;
    wire N__68154;
    wire N__68153;
    wire N__68152;
    wire N__68151;
    wire N__68144;
    wire N__68141;
    wire N__68138;
    wire N__68133;
    wire N__68130;
    wire N__68129;
    wire N__68124;
    wire N__68121;
    wire N__68118;
    wire N__68115;
    wire N__68114;
    wire N__68113;
    wire N__68110;
    wire N__68107;
    wire N__68104;
    wire N__68101;
    wire N__68098;
    wire N__68095;
    wire N__68092;
    wire N__68087;
    wire N__68082;
    wire N__68079;
    wire N__68076;
    wire N__68073;
    wire N__68070;
    wire N__68067;
    wire N__68064;
    wire N__68063;
    wire N__68060;
    wire N__68057;
    wire N__68052;
    wire N__68049;
    wire N__68048;
    wire N__68045;
    wire N__68042;
    wire N__68037;
    wire N__68034;
    wire N__68031;
    wire N__68028;
    wire N__68025;
    wire N__68022;
    wire N__68019;
    wire N__68018;
    wire N__68015;
    wire N__68012;
    wire N__68007;
    wire N__68004;
    wire N__68001;
    wire N__67998;
    wire N__67997;
    wire N__67996;
    wire N__67993;
    wire N__67990;
    wire N__67987;
    wire N__67984;
    wire N__67979;
    wire N__67976;
    wire N__67973;
    wire N__67968;
    wire N__67967;
    wire N__67966;
    wire N__67959;
    wire N__67956;
    wire N__67953;
    wire N__67952;
    wire N__67949;
    wire N__67946;
    wire N__67941;
    wire N__67938;
    wire N__67935;
    wire N__67932;
    wire N__67931;
    wire N__67930;
    wire N__67927;
    wire N__67922;
    wire N__67919;
    wire N__67916;
    wire N__67911;
    wire N__67908;
    wire N__67905;
    wire N__67902;
    wire N__67899;
    wire N__67896;
    wire N__67893;
    wire N__67892;
    wire N__67887;
    wire N__67884;
    wire N__67881;
    wire N__67878;
    wire N__67877;
    wire N__67872;
    wire N__67869;
    wire N__67866;
    wire N__67863;
    wire N__67862;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67852;
    wire N__67849;
    wire N__67846;
    wire N__67843;
    wire N__67836;
    wire N__67833;
    wire N__67830;
    wire N__67827;
    wire N__67826;
    wire N__67823;
    wire N__67820;
    wire N__67815;
    wire N__67812;
    wire N__67809;
    wire N__67808;
    wire N__67805;
    wire N__67802;
    wire N__67797;
    wire N__67794;
    wire N__67791;
    wire N__67788;
    wire N__67785;
    wire N__67782;
    wire N__67779;
    wire N__67778;
    wire N__67773;
    wire N__67770;
    wire N__67767;
    wire N__67764;
    wire N__67761;
    wire N__67760;
    wire N__67759;
    wire N__67758;
    wire N__67757;
    wire N__67756;
    wire N__67753;
    wire N__67752;
    wire N__67749;
    wire N__67746;
    wire N__67743;
    wire N__67742;
    wire N__67741;
    wire N__67732;
    wire N__67731;
    wire N__67730;
    wire N__67729;
    wire N__67718;
    wire N__67715;
    wire N__67708;
    wire N__67703;
    wire N__67698;
    wire N__67695;
    wire N__67694;
    wire N__67693;
    wire N__67690;
    wire N__67685;
    wire N__67682;
    wire N__67679;
    wire N__67674;
    wire N__67673;
    wire N__67670;
    wire N__67667;
    wire N__67662;
    wire N__67659;
    wire N__67656;
    wire N__67655;
    wire N__67652;
    wire N__67651;
    wire N__67650;
    wire N__67649;
    wire N__67648;
    wire N__67647;
    wire N__67646;
    wire N__67645;
    wire N__67644;
    wire N__67643;
    wire N__67636;
    wire N__67633;
    wire N__67632;
    wire N__67631;
    wire N__67628;
    wire N__67627;
    wire N__67626;
    wire N__67625;
    wire N__67624;
    wire N__67623;
    wire N__67620;
    wire N__67609;
    wire N__67606;
    wire N__67599;
    wire N__67586;
    wire N__67583;
    wire N__67580;
    wire N__67573;
    wire N__67570;
    wire N__67565;
    wire N__67560;
    wire N__67559;
    wire N__67556;
    wire N__67553;
    wire N__67550;
    wire N__67547;
    wire N__67546;
    wire N__67545;
    wire N__67542;
    wire N__67539;
    wire N__67534;
    wire N__67527;
    wire N__67526;
    wire N__67525;
    wire N__67520;
    wire N__67519;
    wire N__67518;
    wire N__67517;
    wire N__67514;
    wire N__67511;
    wire N__67506;
    wire N__67503;
    wire N__67500;
    wire N__67497;
    wire N__67492;
    wire N__67485;
    wire N__67482;
    wire N__67479;
    wire N__67478;
    wire N__67475;
    wire N__67472;
    wire N__67467;
    wire N__67464;
    wire N__67461;
    wire N__67458;
    wire N__67457;
    wire N__67454;
    wire N__67451;
    wire N__67446;
    wire N__67445;
    wire N__67444;
    wire N__67441;
    wire N__67438;
    wire N__67435;
    wire N__67428;
    wire N__67427;
    wire N__67426;
    wire N__67425;
    wire N__67422;
    wire N__67419;
    wire N__67416;
    wire N__67413;
    wire N__67410;
    wire N__67405;
    wire N__67398;
    wire N__67395;
    wire N__67392;
    wire N__67389;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67379;
    wire N__67378;
    wire N__67377;
    wire N__67374;
    wire N__67371;
    wire N__67370;
    wire N__67369;
    wire N__67368;
    wire N__67367;
    wire N__67364;
    wire N__67361;
    wire N__67356;
    wire N__67353;
    wire N__67348;
    wire N__67345;
    wire N__67344;
    wire N__67343;
    wire N__67342;
    wire N__67339;
    wire N__67334;
    wire N__67329;
    wire N__67326;
    wire N__67319;
    wire N__67316;
    wire N__67313;
    wire N__67312;
    wire N__67309;
    wire N__67304;
    wire N__67299;
    wire N__67296;
    wire N__67293;
    wire N__67288;
    wire N__67281;
    wire N__67280;
    wire N__67279;
    wire N__67274;
    wire N__67273;
    wire N__67272;
    wire N__67269;
    wire N__67268;
    wire N__67265;
    wire N__67262;
    wire N__67261;
    wire N__67260;
    wire N__67257;
    wire N__67254;
    wire N__67251;
    wire N__67248;
    wire N__67245;
    wire N__67242;
    wire N__67237;
    wire N__67232;
    wire N__67227;
    wire N__67218;
    wire N__67217;
    wire N__67214;
    wire N__67211;
    wire N__67208;
    wire N__67205;
    wire N__67202;
    wire N__67199;
    wire N__67196;
    wire N__67191;
    wire N__67188;
    wire N__67187;
    wire N__67182;
    wire N__67179;
    wire N__67176;
    wire N__67173;
    wire N__67170;
    wire N__67169;
    wire N__67166;
    wire N__67165;
    wire N__67162;
    wire N__67159;
    wire N__67154;
    wire N__67151;
    wire N__67148;
    wire N__67143;
    wire N__67140;
    wire N__67139;
    wire N__67138;
    wire N__67137;
    wire N__67136;
    wire N__67133;
    wire N__67130;
    wire N__67129;
    wire N__67128;
    wire N__67125;
    wire N__67122;
    wire N__67121;
    wire N__67118;
    wire N__67117;
    wire N__67116;
    wire N__67113;
    wire N__67110;
    wire N__67095;
    wire N__67094;
    wire N__67091;
    wire N__67088;
    wire N__67083;
    wire N__67078;
    wire N__67077;
    wire N__67076;
    wire N__67069;
    wire N__67066;
    wire N__67063;
    wire N__67060;
    wire N__67059;
    wire N__67058;
    wire N__67055;
    wire N__67050;
    wire N__67045;
    wire N__67038;
    wire N__67037;
    wire N__67036;
    wire N__67035;
    wire N__67026;
    wire N__67023;
    wire N__67020;
    wire N__67017;
    wire N__67014;
    wire N__67011;
    wire N__67010;
    wire N__67007;
    wire N__67004;
    wire N__67001;
    wire N__66996;
    wire N__66993;
    wire N__66990;
    wire N__66987;
    wire N__66984;
    wire N__66983;
    wire N__66980;
    wire N__66977;
    wire N__66974;
    wire N__66971;
    wire N__66968;
    wire N__66965;
    wire N__66960;
    wire N__66957;
    wire N__66954;
    wire N__66951;
    wire N__66950;
    wire N__66947;
    wire N__66944;
    wire N__66941;
    wire N__66936;
    wire N__66933;
    wire N__66930;
    wire N__66927;
    wire N__66926;
    wire N__66925;
    wire N__66922;
    wire N__66917;
    wire N__66912;
    wire N__66909;
    wire N__66906;
    wire N__66905;
    wire N__66902;
    wire N__66899;
    wire N__66894;
    wire N__66891;
    wire N__66888;
    wire N__66887;
    wire N__66886;
    wire N__66883;
    wire N__66878;
    wire N__66873;
    wire N__66870;
    wire N__66869;
    wire N__66866;
    wire N__66863;
    wire N__66860;
    wire N__66857;
    wire N__66852;
    wire N__66849;
    wire N__66848;
    wire N__66847;
    wire N__66846;
    wire N__66839;
    wire N__66838;
    wire N__66835;
    wire N__66832;
    wire N__66831;
    wire N__66828;
    wire N__66825;
    wire N__66822;
    wire N__66819;
    wire N__66810;
    wire N__66809;
    wire N__66806;
    wire N__66805;
    wire N__66802;
    wire N__66799;
    wire N__66794;
    wire N__66789;
    wire N__66786;
    wire N__66785;
    wire N__66782;
    wire N__66779;
    wire N__66774;
    wire N__66771;
    wire N__66768;
    wire N__66765;
    wire N__66762;
    wire N__66761;
    wire N__66758;
    wire N__66755;
    wire N__66752;
    wire N__66749;
    wire N__66744;
    wire N__66741;
    wire N__66738;
    wire N__66735;
    wire N__66734;
    wire N__66733;
    wire N__66730;
    wire N__66725;
    wire N__66720;
    wire N__66717;
    wire N__66714;
    wire N__66711;
    wire N__66710;
    wire N__66707;
    wire N__66704;
    wire N__66701;
    wire N__66698;
    wire N__66693;
    wire N__66690;
    wire N__66687;
    wire N__66684;
    wire N__66681;
    wire N__66680;
    wire N__66679;
    wire N__66676;
    wire N__66671;
    wire N__66666;
    wire N__66663;
    wire N__66660;
    wire N__66657;
    wire N__66656;
    wire N__66653;
    wire N__66650;
    wire N__66647;
    wire N__66644;
    wire N__66641;
    wire N__66638;
    wire N__66633;
    wire N__66630;
    wire N__66627;
    wire N__66624;
    wire N__66621;
    wire N__66618;
    wire N__66615;
    wire N__66612;
    wire N__66609;
    wire N__66606;
    wire N__66605;
    wire N__66604;
    wire N__66601;
    wire N__66596;
    wire N__66593;
    wire N__66590;
    wire N__66585;
    wire N__66582;
    wire N__66581;
    wire N__66578;
    wire N__66575;
    wire N__66572;
    wire N__66569;
    wire N__66564;
    wire N__66563;
    wire N__66560;
    wire N__66557;
    wire N__66554;
    wire N__66553;
    wire N__66552;
    wire N__66551;
    wire N__66548;
    wire N__66545;
    wire N__66540;
    wire N__66537;
    wire N__66528;
    wire N__66525;
    wire N__66524;
    wire N__66523;
    wire N__66520;
    wire N__66519;
    wire N__66516;
    wire N__66515;
    wire N__66514;
    wire N__66511;
    wire N__66508;
    wire N__66505;
    wire N__66502;
    wire N__66497;
    wire N__66486;
    wire N__66483;
    wire N__66482;
    wire N__66481;
    wire N__66480;
    wire N__66477;
    wire N__66474;
    wire N__66471;
    wire N__66470;
    wire N__66469;
    wire N__66468;
    wire N__66465;
    wire N__66462;
    wire N__66457;
    wire N__66454;
    wire N__66447;
    wire N__66438;
    wire N__66437;
    wire N__66434;
    wire N__66433;
    wire N__66432;
    wire N__66429;
    wire N__66424;
    wire N__66421;
    wire N__66420;
    wire N__66419;
    wire N__66418;
    wire N__66415;
    wire N__66412;
    wire N__66407;
    wire N__66402;
    wire N__66397;
    wire N__66390;
    wire N__66389;
    wire N__66386;
    wire N__66385;
    wire N__66378;
    wire N__66377;
    wire N__66374;
    wire N__66371;
    wire N__66366;
    wire N__66363;
    wire N__66360;
    wire N__66357;
    wire N__66354;
    wire N__66351;
    wire N__66348;
    wire N__66347;
    wire N__66346;
    wire N__66343;
    wire N__66340;
    wire N__66337;
    wire N__66334;
    wire N__66327;
    wire N__66326;
    wire N__66323;
    wire N__66318;
    wire N__66315;
    wire N__66312;
    wire N__66309;
    wire N__66308;
    wire N__66307;
    wire N__66304;
    wire N__66301;
    wire N__66298;
    wire N__66295;
    wire N__66288;
    wire N__66285;
    wire N__66282;
    wire N__66279;
    wire N__66276;
    wire N__66273;
    wire N__66270;
    wire N__66267;
    wire N__66264;
    wire N__66261;
    wire N__66258;
    wire N__66255;
    wire N__66252;
    wire N__66251;
    wire N__66248;
    wire N__66245;
    wire N__66242;
    wire N__66239;
    wire N__66236;
    wire N__66231;
    wire N__66228;
    wire N__66227;
    wire N__66226;
    wire N__66219;
    wire N__66216;
    wire N__66213;
    wire N__66212;
    wire N__66209;
    wire N__66206;
    wire N__66203;
    wire N__66200;
    wire N__66197;
    wire N__66194;
    wire N__66189;
    wire N__66186;
    wire N__66183;
    wire N__66180;
    wire N__66177;
    wire N__66174;
    wire N__66171;
    wire N__66168;
    wire N__66167;
    wire N__66164;
    wire N__66161;
    wire N__66158;
    wire N__66155;
    wire N__66150;
    wire N__66149;
    wire N__66146;
    wire N__66143;
    wire N__66142;
    wire N__66139;
    wire N__66136;
    wire N__66133;
    wire N__66128;
    wire N__66123;
    wire N__66120;
    wire N__66117;
    wire N__66114;
    wire N__66111;
    wire N__66108;
    wire N__66105;
    wire N__66102;
    wire N__66099;
    wire N__66096;
    wire N__66093;
    wire N__66090;
    wire N__66087;
    wire N__66084;
    wire N__66081;
    wire N__66078;
    wire N__66075;
    wire N__66072;
    wire N__66069;
    wire N__66068;
    wire N__66067;
    wire N__66066;
    wire N__66065;
    wire N__66064;
    wire N__66063;
    wire N__66062;
    wire N__66061;
    wire N__66056;
    wire N__66049;
    wire N__66046;
    wire N__66045;
    wire N__66044;
    wire N__66043;
    wire N__66042;
    wire N__66041;
    wire N__66040;
    wire N__66039;
    wire N__66038;
    wire N__66035;
    wire N__66034;
    wire N__66031;
    wire N__66030;
    wire N__66029;
    wire N__66028;
    wire N__66027;
    wire N__66024;
    wire N__66019;
    wire N__66016;
    wire N__66013;
    wire N__66008;
    wire N__66005;
    wire N__66000;
    wire N__65999;
    wire N__65994;
    wire N__65991;
    wire N__65986;
    wire N__65985;
    wire N__65982;
    wire N__65979;
    wire N__65974;
    wire N__65971;
    wire N__65966;
    wire N__65963;
    wire N__65960;
    wire N__65957;
    wire N__65954;
    wire N__65951;
    wire N__65944;
    wire N__65941;
    wire N__65938;
    wire N__65933;
    wire N__65924;
    wire N__65919;
    wire N__65904;
    wire N__65901;
    wire N__65898;
    wire N__65895;
    wire N__65892;
    wire N__65889;
    wire N__65886;
    wire N__65883;
    wire N__65880;
    wire N__65877;
    wire N__65874;
    wire N__65873;
    wire N__65870;
    wire N__65867;
    wire N__65866;
    wire N__65865;
    wire N__65862;
    wire N__65859;
    wire N__65856;
    wire N__65855;
    wire N__65852;
    wire N__65847;
    wire N__65844;
    wire N__65841;
    wire N__65838;
    wire N__65835;
    wire N__65832;
    wire N__65827;
    wire N__65820;
    wire N__65817;
    wire N__65814;
    wire N__65813;
    wire N__65812;
    wire N__65809;
    wire N__65804;
    wire N__65799;
    wire N__65796;
    wire N__65793;
    wire N__65790;
    wire N__65787;
    wire N__65784;
    wire N__65781;
    wire N__65780;
    wire N__65779;
    wire N__65778;
    wire N__65773;
    wire N__65770;
    wire N__65767;
    wire N__65764;
    wire N__65759;
    wire N__65754;
    wire N__65751;
    wire N__65748;
    wire N__65747;
    wire N__65746;
    wire N__65745;
    wire N__65744;
    wire N__65743;
    wire N__65742;
    wire N__65741;
    wire N__65740;
    wire N__65739;
    wire N__65738;
    wire N__65737;
    wire N__65736;
    wire N__65735;
    wire N__65734;
    wire N__65733;
    wire N__65730;
    wire N__65727;
    wire N__65724;
    wire N__65719;
    wire N__65716;
    wire N__65707;
    wire N__65702;
    wire N__65699;
    wire N__65698;
    wire N__65697;
    wire N__65696;
    wire N__65689;
    wire N__65686;
    wire N__65683;
    wire N__65682;
    wire N__65681;
    wire N__65680;
    wire N__65679;
    wire N__65678;
    wire N__65673;
    wire N__65670;
    wire N__65665;
    wire N__65662;
    wire N__65659;
    wire N__65656;
    wire N__65653;
    wire N__65650;
    wire N__65645;
    wire N__65638;
    wire N__65633;
    wire N__65630;
    wire N__65623;
    wire N__65618;
    wire N__65601;
    wire N__65598;
    wire N__65595;
    wire N__65592;
    wire N__65589;
    wire N__65586;
    wire N__65583;
    wire N__65580;
    wire N__65577;
    wire N__65574;
    wire N__65571;
    wire N__65568;
    wire N__65565;
    wire N__65562;
    wire N__65559;
    wire N__65556;
    wire N__65553;
    wire N__65550;
    wire N__65547;
    wire N__65544;
    wire N__65541;
    wire N__65538;
    wire N__65535;
    wire N__65532;
    wire N__65529;
    wire N__65526;
    wire N__65523;
    wire N__65520;
    wire N__65517;
    wire N__65514;
    wire N__65511;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65490;
    wire N__65487;
    wire N__65484;
    wire N__65481;
    wire N__65480;
    wire N__65475;
    wire N__65472;
    wire N__65469;
    wire N__65466;
    wire N__65463;
    wire N__65460;
    wire N__65459;
    wire N__65458;
    wire N__65457;
    wire N__65456;
    wire N__65453;
    wire N__65452;
    wire N__65451;
    wire N__65450;
    wire N__65449;
    wire N__65448;
    wire N__65445;
    wire N__65442;
    wire N__65441;
    wire N__65438;
    wire N__65431;
    wire N__65430;
    wire N__65429;
    wire N__65426;
    wire N__65423;
    wire N__65420;
    wire N__65417;
    wire N__65414;
    wire N__65411;
    wire N__65408;
    wire N__65407;
    wire N__65406;
    wire N__65403;
    wire N__65400;
    wire N__65395;
    wire N__65390;
    wire N__65385;
    wire N__65384;
    wire N__65381;
    wire N__65376;
    wire N__65371;
    wire N__65360;
    wire N__65357;
    wire N__65350;
    wire N__65345;
    wire N__65342;
    wire N__65339;
    wire N__65336;
    wire N__65333;
    wire N__65328;
    wire N__65325;
    wire N__65322;
    wire N__65319;
    wire N__65318;
    wire N__65315;
    wire N__65312;
    wire N__65309;
    wire N__65304;
    wire N__65303;
    wire N__65298;
    wire N__65295;
    wire N__65292;
    wire N__65291;
    wire N__65288;
    wire N__65285;
    wire N__65280;
    wire N__65277;
    wire N__65274;
    wire N__65271;
    wire N__65268;
    wire N__65265;
    wire N__65262;
    wire N__65259;
    wire N__65258;
    wire N__65257;
    wire N__65250;
    wire N__65247;
    wire N__65244;
    wire N__65243;
    wire N__65238;
    wire N__65235;
    wire N__65232;
    wire N__65231;
    wire N__65228;
    wire N__65225;
    wire N__65222;
    wire N__65221;
    wire N__65218;
    wire N__65215;
    wire N__65212;
    wire N__65211;
    wire N__65210;
    wire N__65209;
    wire N__65202;
    wire N__65201;
    wire N__65200;
    wire N__65197;
    wire N__65194;
    wire N__65191;
    wire N__65188;
    wire N__65183;
    wire N__65180;
    wire N__65175;
    wire N__65172;
    wire N__65169;
    wire N__65166;
    wire N__65163;
    wire N__65160;
    wire N__65157;
    wire N__65148;
    wire N__65147;
    wire N__65146;
    wire N__65143;
    wire N__65142;
    wire N__65139;
    wire N__65132;
    wire N__65127;
    wire N__65126;
    wire N__65125;
    wire N__65124;
    wire N__65121;
    wire N__65118;
    wire N__65115;
    wire N__65112;
    wire N__65109;
    wire N__65106;
    wire N__65101;
    wire N__65096;
    wire N__65093;
    wire N__65090;
    wire N__65085;
    wire N__65084;
    wire N__65079;
    wire N__65076;
    wire N__65075;
    wire N__65070;
    wire N__65067;
    wire N__65066;
    wire N__65065;
    wire N__65062;
    wire N__65059;
    wire N__65056;
    wire N__65049;
    wire N__65048;
    wire N__65043;
    wire N__65040;
    wire N__65039;
    wire N__65036;
    wire N__65033;
    wire N__65028;
    wire N__65027;
    wire N__65024;
    wire N__65021;
    wire N__65018;
    wire N__65015;
    wire N__65012;
    wire N__65009;
    wire N__65006;
    wire N__65003;
    wire N__64998;
    wire N__64997;
    wire N__64996;
    wire N__64995;
    wire N__64994;
    wire N__64989;
    wire N__64986;
    wire N__64985;
    wire N__64980;
    wire N__64977;
    wire N__64974;
    wire N__64971;
    wire N__64968;
    wire N__64967;
    wire N__64966;
    wire N__64963;
    wire N__64960;
    wire N__64957;
    wire N__64954;
    wire N__64951;
    wire N__64948;
    wire N__64945;
    wire N__64942;
    wire N__64933;
    wire N__64930;
    wire N__64925;
    wire N__64920;
    wire N__64917;
    wire N__64914;
    wire N__64911;
    wire N__64908;
    wire N__64905;
    wire N__64902;
    wire N__64899;
    wire N__64896;
    wire N__64893;
    wire N__64890;
    wire N__64887;
    wire N__64884;
    wire N__64881;
    wire N__64878;
    wire N__64875;
    wire N__64872;
    wire N__64869;
    wire N__64866;
    wire N__64865;
    wire N__64862;
    wire N__64861;
    wire N__64858;
    wire N__64855;
    wire N__64852;
    wire N__64845;
    wire N__64842;
    wire N__64839;
    wire N__64836;
    wire N__64833;
    wire N__64832;
    wire N__64829;
    wire N__64828;
    wire N__64825;
    wire N__64822;
    wire N__64819;
    wire N__64814;
    wire N__64811;
    wire N__64806;
    wire N__64803;
    wire N__64802;
    wire N__64799;
    wire N__64796;
    wire N__64791;
    wire N__64790;
    wire N__64787;
    wire N__64784;
    wire N__64779;
    wire N__64778;
    wire N__64775;
    wire N__64772;
    wire N__64767;
    wire N__64764;
    wire N__64761;
    wire N__64758;
    wire N__64755;
    wire N__64754;
    wire N__64751;
    wire N__64748;
    wire N__64743;
    wire N__64740;
    wire N__64737;
    wire N__64736;
    wire N__64735;
    wire N__64734;
    wire N__64733;
    wire N__64732;
    wire N__64731;
    wire N__64730;
    wire N__64729;
    wire N__64728;
    wire N__64727;
    wire N__64726;
    wire N__64723;
    wire N__64722;
    wire N__64719;
    wire N__64716;
    wire N__64713;
    wire N__64710;
    wire N__64707;
    wire N__64704;
    wire N__64701;
    wire N__64698;
    wire N__64687;
    wire N__64682;
    wire N__64679;
    wire N__64676;
    wire N__64673;
    wire N__64668;
    wire N__64663;
    wire N__64650;
    wire N__64649;
    wire N__64644;
    wire N__64641;
    wire N__64638;
    wire N__64635;
    wire N__64632;
    wire N__64629;
    wire N__64626;
    wire N__64623;
    wire N__64620;
    wire N__64617;
    wire N__64614;
    wire N__64611;
    wire N__64608;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64590;
    wire N__64587;
    wire N__64584;
    wire N__64581;
    wire N__64578;
    wire N__64575;
    wire N__64572;
    wire N__64569;
    wire N__64566;
    wire N__64563;
    wire N__64560;
    wire N__64557;
    wire N__64554;
    wire N__64551;
    wire N__64548;
    wire N__64545;
    wire N__64542;
    wire N__64539;
    wire N__64536;
    wire N__64533;
    wire N__64530;
    wire N__64527;
    wire N__64524;
    wire N__64521;
    wire N__64518;
    wire N__64515;
    wire N__64512;
    wire N__64509;
    wire N__64506;
    wire N__64503;
    wire N__64500;
    wire N__64497;
    wire N__64494;
    wire N__64491;
    wire N__64488;
    wire N__64485;
    wire N__64482;
    wire N__64479;
    wire N__64476;
    wire N__64473;
    wire N__64470;
    wire N__64467;
    wire N__64464;
    wire N__64461;
    wire N__64458;
    wire N__64455;
    wire N__64452;
    wire N__64449;
    wire N__64446;
    wire N__64443;
    wire N__64440;
    wire N__64437;
    wire N__64434;
    wire N__64431;
    wire N__64428;
    wire N__64425;
    wire N__64422;
    wire N__64419;
    wire N__64416;
    wire N__64413;
    wire N__64410;
    wire N__64407;
    wire N__64404;
    wire N__64401;
    wire N__64398;
    wire N__64395;
    wire N__64392;
    wire N__64389;
    wire N__64386;
    wire N__64383;
    wire N__64380;
    wire N__64377;
    wire N__64376;
    wire N__64371;
    wire N__64368;
    wire N__64365;
    wire N__64362;
    wire N__64359;
    wire N__64356;
    wire N__64353;
    wire N__64350;
    wire N__64347;
    wire N__64346;
    wire N__64341;
    wire N__64338;
    wire N__64335;
    wire N__64332;
    wire N__64329;
    wire N__64326;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64316;
    wire N__64311;
    wire N__64308;
    wire N__64305;
    wire N__64302;
    wire N__64299;
    wire N__64296;
    wire N__64293;
    wire N__64292;
    wire N__64287;
    wire N__64284;
    wire N__64281;
    wire N__64278;
    wire N__64277;
    wire N__64274;
    wire N__64269;
    wire N__64266;
    wire N__64263;
    wire N__64260;
    wire N__64257;
    wire N__64254;
    wire N__64251;
    wire N__64248;
    wire N__64245;
    wire N__64242;
    wire N__64239;
    wire N__64236;
    wire N__64235;
    wire N__64232;
    wire N__64229;
    wire N__64226;
    wire N__64225;
    wire N__64222;
    wire N__64219;
    wire N__64216;
    wire N__64213;
    wire N__64212;
    wire N__64209;
    wire N__64206;
    wire N__64203;
    wire N__64200;
    wire N__64191;
    wire N__64188;
    wire N__64185;
    wire N__64184;
    wire N__64183;
    wire N__64180;
    wire N__64175;
    wire N__64170;
    wire N__64167;
    wire N__64164;
    wire N__64163;
    wire N__64160;
    wire N__64159;
    wire N__64156;
    wire N__64153;
    wire N__64148;
    wire N__64145;
    wire N__64142;
    wire N__64137;
    wire N__64134;
    wire N__64131;
    wire N__64128;
    wire N__64127;
    wire N__64126;
    wire N__64123;
    wire N__64118;
    wire N__64115;
    wire N__64112;
    wire N__64107;
    wire N__64104;
    wire N__64101;
    wire N__64100;
    wire N__64099;
    wire N__64096;
    wire N__64091;
    wire N__64088;
    wire N__64085;
    wire N__64082;
    wire N__64079;
    wire N__64074;
    wire N__64071;
    wire N__64068;
    wire N__64065;
    wire N__64062;
    wire N__64059;
    wire N__64056;
    wire N__64055;
    wire N__64054;
    wire N__64051;
    wire N__64048;
    wire N__64045;
    wire N__64042;
    wire N__64037;
    wire N__64034;
    wire N__64031;
    wire N__64026;
    wire N__64023;
    wire N__64022;
    wire N__64019;
    wire N__64018;
    wire N__64015;
    wire N__64012;
    wire N__64011;
    wire N__64010;
    wire N__64007;
    wire N__64002;
    wire N__63997;
    wire N__63994;
    wire N__63991;
    wire N__63986;
    wire N__63981;
    wire N__63978;
    wire N__63977;
    wire N__63976;
    wire N__63973;
    wire N__63968;
    wire N__63963;
    wire N__63960;
    wire N__63959;
    wire N__63956;
    wire N__63953;
    wire N__63950;
    wire N__63947;
    wire N__63944;
    wire N__63941;
    wire N__63936;
    wire N__63933;
    wire N__63930;
    wire N__63929;
    wire N__63928;
    wire N__63925;
    wire N__63920;
    wire N__63915;
    wire N__63912;
    wire N__63909;
    wire N__63906;
    wire N__63903;
    wire N__63900;
    wire N__63897;
    wire N__63894;
    wire N__63891;
    wire N__63888;
    wire N__63885;
    wire N__63884;
    wire N__63881;
    wire N__63878;
    wire N__63875;
    wire N__63870;
    wire N__63867;
    wire N__63866;
    wire N__63865;
    wire N__63862;
    wire N__63859;
    wire N__63856;
    wire N__63855;
    wire N__63850;
    wire N__63845;
    wire N__63840;
    wire N__63837;
    wire N__63834;
    wire N__63831;
    wire N__63828;
    wire N__63825;
    wire N__63822;
    wire N__63819;
    wire N__63816;
    wire N__63813;
    wire N__63810;
    wire N__63807;
    wire N__63804;
    wire N__63801;
    wire N__63798;
    wire N__63795;
    wire N__63792;
    wire N__63789;
    wire N__63786;
    wire N__63783;
    wire N__63780;
    wire N__63777;
    wire N__63774;
    wire N__63771;
    wire N__63768;
    wire N__63765;
    wire N__63762;
    wire N__63759;
    wire N__63756;
    wire N__63753;
    wire N__63750;
    wire N__63747;
    wire N__63744;
    wire N__63741;
    wire N__63738;
    wire N__63735;
    wire N__63732;
    wire N__63729;
    wire N__63726;
    wire N__63723;
    wire N__63720;
    wire N__63717;
    wire N__63714;
    wire N__63711;
    wire N__63708;
    wire N__63705;
    wire N__63702;
    wire N__63699;
    wire N__63696;
    wire N__63693;
    wire N__63690;
    wire N__63687;
    wire N__63684;
    wire N__63681;
    wire N__63678;
    wire N__63675;
    wire N__63672;
    wire N__63669;
    wire N__63666;
    wire N__63663;
    wire N__63660;
    wire N__63657;
    wire N__63654;
    wire N__63651;
    wire N__63648;
    wire N__63645;
    wire N__63642;
    wire N__63641;
    wire N__63638;
    wire N__63635;
    wire N__63632;
    wire N__63629;
    wire N__63626;
    wire N__63621;
    wire N__63618;
    wire N__63615;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63600;
    wire N__63597;
    wire N__63594;
    wire N__63591;
    wire N__63588;
    wire N__63585;
    wire N__63582;
    wire N__63579;
    wire N__63576;
    wire N__63573;
    wire N__63570;
    wire N__63567;
    wire N__63564;
    wire N__63561;
    wire N__63558;
    wire N__63555;
    wire N__63552;
    wire N__63549;
    wire N__63546;
    wire N__63543;
    wire N__63540;
    wire N__63537;
    wire N__63534;
    wire N__63533;
    wire N__63530;
    wire N__63527;
    wire N__63524;
    wire N__63521;
    wire N__63516;
    wire N__63513;
    wire N__63510;
    wire N__63507;
    wire N__63504;
    wire N__63503;
    wire N__63502;
    wire N__63501;
    wire N__63500;
    wire N__63499;
    wire N__63498;
    wire N__63495;
    wire N__63492;
    wire N__63491;
    wire N__63490;
    wire N__63489;
    wire N__63488;
    wire N__63485;
    wire N__63482;
    wire N__63479;
    wire N__63476;
    wire N__63473;
    wire N__63470;
    wire N__63467;
    wire N__63464;
    wire N__63463;
    wire N__63462;
    wire N__63459;
    wire N__63454;
    wire N__63447;
    wire N__63446;
    wire N__63445;
    wire N__63434;
    wire N__63433;
    wire N__63432;
    wire N__63429;
    wire N__63426;
    wire N__63421;
    wire N__63420;
    wire N__63419;
    wire N__63416;
    wire N__63413;
    wire N__63410;
    wire N__63407;
    wire N__63402;
    wire N__63395;
    wire N__63390;
    wire N__63385;
    wire N__63372;
    wire N__63371;
    wire N__63370;
    wire N__63369;
    wire N__63368;
    wire N__63365;
    wire N__63364;
    wire N__63363;
    wire N__63362;
    wire N__63361;
    wire N__63360;
    wire N__63357;
    wire N__63352;
    wire N__63349;
    wire N__63346;
    wire N__63343;
    wire N__63342;
    wire N__63339;
    wire N__63336;
    wire N__63333;
    wire N__63330;
    wire N__63329;
    wire N__63328;
    wire N__63327;
    wire N__63326;
    wire N__63321;
    wire N__63318;
    wire N__63313;
    wire N__63310;
    wire N__63307;
    wire N__63300;
    wire N__63295;
    wire N__63292;
    wire N__63289;
    wire N__63280;
    wire N__63267;
    wire N__63266;
    wire N__63265;
    wire N__63264;
    wire N__63263;
    wire N__63260;
    wire N__63259;
    wire N__63258;
    wire N__63257;
    wire N__63254;
    wire N__63251;
    wire N__63250;
    wire N__63249;
    wire N__63246;
    wire N__63243;
    wire N__63240;
    wire N__63235;
    wire N__63232;
    wire N__63227;
    wire N__63224;
    wire N__63223;
    wire N__63222;
    wire N__63219;
    wire N__63218;
    wire N__63217;
    wire N__63214;
    wire N__63205;
    wire N__63200;
    wire N__63197;
    wire N__63194;
    wire N__63191;
    wire N__63188;
    wire N__63185;
    wire N__63168;
    wire N__63165;
    wire N__63164;
    wire N__63163;
    wire N__63162;
    wire N__63161;
    wire N__63160;
    wire N__63157;
    wire N__63156;
    wire N__63155;
    wire N__63152;
    wire N__63149;
    wire N__63148;
    wire N__63145;
    wire N__63144;
    wire N__63143;
    wire N__63142;
    wire N__63141;
    wire N__63138;
    wire N__63135;
    wire N__63132;
    wire N__63129;
    wire N__63126;
    wire N__63121;
    wire N__63118;
    wire N__63117;
    wire N__63116;
    wire N__63113;
    wire N__63108;
    wire N__63103;
    wire N__63100;
    wire N__63091;
    wire N__63086;
    wire N__63081;
    wire N__63066;
    wire N__63063;
    wire N__63060;
    wire N__63059;
    wire N__63056;
    wire N__63055;
    wire N__63054;
    wire N__63051;
    wire N__63048;
    wire N__63047;
    wire N__63046;
    wire N__63045;
    wire N__63044;
    wire N__63041;
    wire N__63038;
    wire N__63037;
    wire N__63036;
    wire N__63035;
    wire N__63034;
    wire N__63029;
    wire N__63026;
    wire N__63023;
    wire N__63020;
    wire N__63017;
    wire N__63014;
    wire N__63011;
    wire N__63008;
    wire N__63003;
    wire N__63000;
    wire N__62999;
    wire N__62998;
    wire N__62997;
    wire N__62996;
    wire N__62995;
    wire N__62994;
    wire N__62991;
    wire N__62988;
    wire N__62981;
    wire N__62972;
    wire N__62969;
    wire N__62966;
    wire N__62963;
    wire N__62960;
    wire N__62957;
    wire N__62956;
    wire N__62953;
    wire N__62952;
    wire N__62949;
    wire N__62948;
    wire N__62943;
    wire N__62940;
    wire N__62937;
    wire N__62930;
    wire N__62927;
    wire N__62922;
    wire N__62913;
    wire N__62898;
    wire N__62895;
    wire N__62892;
    wire N__62889;
    wire N__62886;
    wire N__62883;
    wire N__62880;
    wire N__62879;
    wire N__62876;
    wire N__62873;
    wire N__62868;
    wire N__62865;
    wire N__62862;
    wire N__62859;
    wire N__62856;
    wire N__62853;
    wire N__62850;
    wire N__62847;
    wire N__62846;
    wire N__62845;
    wire N__62842;
    wire N__62837;
    wire N__62832;
    wire N__62829;
    wire N__62826;
    wire N__62823;
    wire N__62820;
    wire N__62817;
    wire N__62814;
    wire N__62811;
    wire N__62810;
    wire N__62807;
    wire N__62804;
    wire N__62799;
    wire N__62796;
    wire N__62793;
    wire N__62790;
    wire N__62789;
    wire N__62788;
    wire N__62785;
    wire N__62778;
    wire N__62775;
    wire N__62772;
    wire N__62769;
    wire N__62766;
    wire N__62765;
    wire N__62764;
    wire N__62761;
    wire N__62756;
    wire N__62751;
    wire N__62750;
    wire N__62749;
    wire N__62746;
    wire N__62743;
    wire N__62740;
    wire N__62739;
    wire N__62738;
    wire N__62737;
    wire N__62734;
    wire N__62727;
    wire N__62724;
    wire N__62721;
    wire N__62720;
    wire N__62719;
    wire N__62718;
    wire N__62717;
    wire N__62716;
    wire N__62715;
    wire N__62714;
    wire N__62713;
    wire N__62712;
    wire N__62711;
    wire N__62710;
    wire N__62709;
    wire N__62708;
    wire N__62707;
    wire N__62702;
    wire N__62695;
    wire N__62694;
    wire N__62693;
    wire N__62690;
    wire N__62687;
    wire N__62684;
    wire N__62683;
    wire N__62682;
    wire N__62679;
    wire N__62678;
    wire N__62677;
    wire N__62676;
    wire N__62675;
    wire N__62674;
    wire N__62673;
    wire N__62672;
    wire N__62671;
    wire N__62668;
    wire N__62665;
    wire N__62662;
    wire N__62659;
    wire N__62656;
    wire N__62655;
    wire N__62654;
    wire N__62653;
    wire N__62652;
    wire N__62649;
    wire N__62646;
    wire N__62643;
    wire N__62640;
    wire N__62639;
    wire N__62634;
    wire N__62633;
    wire N__62632;
    wire N__62629;
    wire N__62622;
    wire N__62619;
    wire N__62612;
    wire N__62605;
    wire N__62604;
    wire N__62601;
    wire N__62598;
    wire N__62597;
    wire N__62594;
    wire N__62593;
    wire N__62592;
    wire N__62591;
    wire N__62590;
    wire N__62583;
    wire N__62582;
    wire N__62581;
    wire N__62578;
    wire N__62571;
    wire N__62570;
    wire N__62569;
    wire N__62568;
    wire N__62565;
    wire N__62562;
    wire N__62559;
    wire N__62558;
    wire N__62545;
    wire N__62542;
    wire N__62535;
    wire N__62530;
    wire N__62525;
    wire N__62518;
    wire N__62509;
    wire N__62504;
    wire N__62501;
    wire N__62496;
    wire N__62491;
    wire N__62476;
    wire N__62471;
    wire N__62464;
    wire N__62453;
    wire N__62450;
    wire N__62443;
    wire N__62440;
    wire N__62437;
    wire N__62434;
    wire N__62431;
    wire N__62424;
    wire N__62421;
    wire N__62418;
    wire N__62415;
    wire N__62414;
    wire N__62411;
    wire N__62408;
    wire N__62403;
    wire N__62400;
    wire N__62397;
    wire N__62394;
    wire N__62391;
    wire N__62390;
    wire N__62389;
    wire N__62386;
    wire N__62383;
    wire N__62380;
    wire N__62377;
    wire N__62374;
    wire N__62367;
    wire N__62366;
    wire N__62365;
    wire N__62362;
    wire N__62359;
    wire N__62356;
    wire N__62353;
    wire N__62346;
    wire N__62343;
    wire N__62340;
    wire N__62337;
    wire N__62334;
    wire N__62331;
    wire N__62328;
    wire N__62325;
    wire N__62322;
    wire N__62319;
    wire N__62318;
    wire N__62315;
    wire N__62312;
    wire N__62307;
    wire N__62306;
    wire N__62303;
    wire N__62300;
    wire N__62297;
    wire N__62292;
    wire N__62291;
    wire N__62288;
    wire N__62285;
    wire N__62282;
    wire N__62279;
    wire N__62274;
    wire N__62271;
    wire N__62270;
    wire N__62267;
    wire N__62264;
    wire N__62259;
    wire N__62256;
    wire N__62253;
    wire N__62250;
    wire N__62247;
    wire N__62244;
    wire N__62241;
    wire N__62238;
    wire N__62235;
    wire N__62232;
    wire N__62229;
    wire N__62228;
    wire N__62223;
    wire N__62220;
    wire N__62217;
    wire N__62216;
    wire N__62213;
    wire N__62210;
    wire N__62205;
    wire N__62202;
    wire N__62199;
    wire N__62196;
    wire N__62193;
    wire N__62190;
    wire N__62187;
    wire N__62184;
    wire N__62181;
    wire N__62178;
    wire N__62175;
    wire N__62172;
    wire N__62169;
    wire N__62166;
    wire N__62165;
    wire N__62162;
    wire N__62159;
    wire N__62156;
    wire N__62153;
    wire N__62152;
    wire N__62151;
    wire N__62148;
    wire N__62145;
    wire N__62142;
    wire N__62141;
    wire N__62140;
    wire N__62139;
    wire N__62138;
    wire N__62137;
    wire N__62134;
    wire N__62127;
    wire N__62124;
    wire N__62121;
    wire N__62118;
    wire N__62115;
    wire N__62112;
    wire N__62109;
    wire N__62104;
    wire N__62103;
    wire N__62098;
    wire N__62093;
    wire N__62088;
    wire N__62085;
    wire N__62080;
    wire N__62077;
    wire N__62070;
    wire N__62067;
    wire N__62064;
    wire N__62061;
    wire N__62058;
    wire N__62055;
    wire N__62052;
    wire N__62049;
    wire N__62048;
    wire N__62045;
    wire N__62044;
    wire N__62041;
    wire N__62038;
    wire N__62035;
    wire N__62028;
    wire N__62025;
    wire N__62024;
    wire N__62023;
    wire N__62022;
    wire N__62019;
    wire N__62016;
    wire N__62013;
    wire N__62012;
    wire N__62009;
    wire N__62004;
    wire N__61999;
    wire N__61994;
    wire N__61989;
    wire N__61986;
    wire N__61983;
    wire N__61980;
    wire N__61977;
    wire N__61974;
    wire N__61971;
    wire N__61968;
    wire N__61965;
    wire N__61964;
    wire N__61963;
    wire N__61960;
    wire N__61955;
    wire N__61950;
    wire N__61947;
    wire N__61944;
    wire N__61941;
    wire N__61938;
    wire N__61937;
    wire N__61936;
    wire N__61933;
    wire N__61928;
    wire N__61923;
    wire N__61920;
    wire N__61917;
    wire N__61914;
    wire N__61913;
    wire N__61912;
    wire N__61911;
    wire N__61910;
    wire N__61907;
    wire N__61902;
    wire N__61899;
    wire N__61896;
    wire N__61893;
    wire N__61892;
    wire N__61891;
    wire N__61888;
    wire N__61885;
    wire N__61882;
    wire N__61879;
    wire N__61876;
    wire N__61873;
    wire N__61870;
    wire N__61863;
    wire N__61854;
    wire N__61851;
    wire N__61848;
    wire N__61845;
    wire N__61842;
    wire N__61839;
    wire N__61838;
    wire N__61835;
    wire N__61834;
    wire N__61833;
    wire N__61830;
    wire N__61827;
    wire N__61824;
    wire N__61821;
    wire N__61818;
    wire N__61815;
    wire N__61814;
    wire N__61811;
    wire N__61810;
    wire N__61809;
    wire N__61806;
    wire N__61805;
    wire N__61802;
    wire N__61799;
    wire N__61796;
    wire N__61793;
    wire N__61788;
    wire N__61785;
    wire N__61782;
    wire N__61779;
    wire N__61776;
    wire N__61773;
    wire N__61766;
    wire N__61761;
    wire N__61758;
    wire N__61749;
    wire N__61746;
    wire N__61745;
    wire N__61744;
    wire N__61739;
    wire N__61738;
    wire N__61735;
    wire N__61732;
    wire N__61729;
    wire N__61724;
    wire N__61721;
    wire N__61716;
    wire N__61713;
    wire N__61710;
    wire N__61709;
    wire N__61704;
    wire N__61701;
    wire N__61698;
    wire N__61695;
    wire N__61692;
    wire N__61691;
    wire N__61690;
    wire N__61685;
    wire N__61682;
    wire N__61679;
    wire N__61674;
    wire N__61673;
    wire N__61672;
    wire N__61671;
    wire N__61670;
    wire N__61669;
    wire N__61666;
    wire N__61665;
    wire N__61664;
    wire N__61661;
    wire N__61656;
    wire N__61655;
    wire N__61652;
    wire N__61649;
    wire N__61646;
    wire N__61643;
    wire N__61640;
    wire N__61639;
    wire N__61638;
    wire N__61637;
    wire N__61636;
    wire N__61635;
    wire N__61634;
    wire N__61629;
    wire N__61626;
    wire N__61623;
    wire N__61614;
    wire N__61609;
    wire N__61606;
    wire N__61605;
    wire N__61602;
    wire N__61597;
    wire N__61592;
    wire N__61591;
    wire N__61584;
    wire N__61581;
    wire N__61578;
    wire N__61573;
    wire N__61570;
    wire N__61567;
    wire N__61562;
    wire N__61559;
    wire N__61548;
    wire N__61545;
    wire N__61542;
    wire N__61541;
    wire N__61538;
    wire N__61535;
    wire N__61530;
    wire N__61527;
    wire N__61524;
    wire N__61521;
    wire N__61518;
    wire N__61515;
    wire N__61512;
    wire N__61509;
    wire N__61506;
    wire N__61503;
    wire N__61500;
    wire N__61497;
    wire N__61494;
    wire N__61491;
    wire N__61488;
    wire N__61485;
    wire N__61482;
    wire N__61479;
    wire N__61478;
    wire N__61477;
    wire N__61474;
    wire N__61471;
    wire N__61468;
    wire N__61461;
    wire N__61458;
    wire N__61455;
    wire N__61452;
    wire N__61449;
    wire N__61446;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61434;
    wire N__61431;
    wire N__61428;
    wire N__61425;
    wire N__61422;
    wire N__61419;
    wire N__61416;
    wire N__61413;
    wire N__61410;
    wire N__61407;
    wire N__61404;
    wire N__61401;
    wire N__61398;
    wire N__61395;
    wire N__61394;
    wire N__61391;
    wire N__61388;
    wire N__61383;
    wire N__61380;
    wire N__61379;
    wire N__61378;
    wire N__61375;
    wire N__61372;
    wire N__61369;
    wire N__61362;
    wire N__61361;
    wire N__61360;
    wire N__61359;
    wire N__61358;
    wire N__61353;
    wire N__61348;
    wire N__61345;
    wire N__61338;
    wire N__61335;
    wire N__61334;
    wire N__61331;
    wire N__61328;
    wire N__61323;
    wire N__61320;
    wire N__61317;
    wire N__61314;
    wire N__61311;
    wire N__61308;
    wire N__61305;
    wire N__61302;
    wire N__61299;
    wire N__61298;
    wire N__61295;
    wire N__61292;
    wire N__61287;
    wire N__61286;
    wire N__61281;
    wire N__61278;
    wire N__61275;
    wire N__61274;
    wire N__61271;
    wire N__61268;
    wire N__61267;
    wire N__61262;
    wire N__61259;
    wire N__61254;
    wire N__61253;
    wire N__61250;
    wire N__61249;
    wire N__61246;
    wire N__61241;
    wire N__61238;
    wire N__61233;
    wire N__61230;
    wire N__61229;
    wire N__61228;
    wire N__61225;
    wire N__61220;
    wire N__61215;
    wire N__61214;
    wire N__61213;
    wire N__61208;
    wire N__61205;
    wire N__61200;
    wire N__61199;
    wire N__61196;
    wire N__61193;
    wire N__61188;
    wire N__61185;
    wire N__61182;
    wire N__61181;
    wire N__61180;
    wire N__61177;
    wire N__61172;
    wire N__61167;
    wire N__61166;
    wire N__61163;
    wire N__61160;
    wire N__61155;
    wire N__61152;
    wire N__61151;
    wire N__61150;
    wire N__61147;
    wire N__61142;
    wire N__61137;
    wire N__61134;
    wire N__61133;
    wire N__61132;
    wire N__61129;
    wire N__61124;
    wire N__61119;
    wire N__61116;
    wire N__61115;
    wire N__61112;
    wire N__61109;
    wire N__61104;
    wire N__61101;
    wire N__61100;
    wire N__61099;
    wire N__61096;
    wire N__61091;
    wire N__61086;
    wire N__61085;
    wire N__61082;
    wire N__61079;
    wire N__61076;
    wire N__61073;
    wire N__61068;
    wire N__61065;
    wire N__61062;
    wire N__61059;
    wire N__61056;
    wire N__61055;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61038;
    wire N__61037;
    wire N__61034;
    wire N__61033;
    wire N__61030;
    wire N__61027;
    wire N__61024;
    wire N__61017;
    wire N__61014;
    wire N__61011;
    wire N__61010;
    wire N__61007;
    wire N__61004;
    wire N__60999;
    wire N__60996;
    wire N__60995;
    wire N__60992;
    wire N__60989;
    wire N__60984;
    wire N__60983;
    wire N__60980;
    wire N__60977;
    wire N__60972;
    wire N__60971;
    wire N__60968;
    wire N__60965;
    wire N__60960;
    wire N__60957;
    wire N__60954;
    wire N__60951;
    wire N__60948;
    wire N__60947;
    wire N__60942;
    wire N__60939;
    wire N__60936;
    wire N__60933;
    wire N__60932;
    wire N__60931;
    wire N__60928;
    wire N__60923;
    wire N__60920;
    wire N__60917;
    wire N__60912;
    wire N__60909;
    wire N__60906;
    wire N__60903;
    wire N__60900;
    wire N__60899;
    wire N__60894;
    wire N__60893;
    wire N__60890;
    wire N__60887;
    wire N__60884;
    wire N__60879;
    wire N__60876;
    wire N__60873;
    wire N__60872;
    wire N__60871;
    wire N__60868;
    wire N__60863;
    wire N__60858;
    wire N__60855;
    wire N__60852;
    wire N__60849;
    wire N__60846;
    wire N__60845;
    wire N__60842;
    wire N__60839;
    wire N__60834;
    wire N__60831;
    wire N__60828;
    wire N__60825;
    wire N__60824;
    wire N__60823;
    wire N__60820;
    wire N__60815;
    wire N__60812;
    wire N__60809;
    wire N__60804;
    wire N__60803;
    wire N__60800;
    wire N__60797;
    wire N__60794;
    wire N__60791;
    wire N__60786;
    wire N__60783;
    wire N__60780;
    wire N__60777;
    wire N__60774;
    wire N__60771;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60756;
    wire N__60753;
    wire N__60750;
    wire N__60747;
    wire N__60744;
    wire N__60741;
    wire N__60740;
    wire N__60737;
    wire N__60734;
    wire N__60729;
    wire N__60726;
    wire N__60725;
    wire N__60724;
    wire N__60723;
    wire N__60720;
    wire N__60717;
    wire N__60714;
    wire N__60713;
    wire N__60710;
    wire N__60707;
    wire N__60702;
    wire N__60699;
    wire N__60696;
    wire N__60693;
    wire N__60688;
    wire N__60685;
    wire N__60682;
    wire N__60679;
    wire N__60676;
    wire N__60669;
    wire N__60668;
    wire N__60665;
    wire N__60662;
    wire N__60657;
    wire N__60656;
    wire N__60655;
    wire N__60654;
    wire N__60653;
    wire N__60652;
    wire N__60649;
    wire N__60646;
    wire N__60643;
    wire N__60642;
    wire N__60639;
    wire N__60636;
    wire N__60635;
    wire N__60632;
    wire N__60631;
    wire N__60630;
    wire N__60629;
    wire N__60622;
    wire N__60621;
    wire N__60618;
    wire N__60613;
    wire N__60606;
    wire N__60603;
    wire N__60602;
    wire N__60599;
    wire N__60598;
    wire N__60597;
    wire N__60596;
    wire N__60595;
    wire N__60594;
    wire N__60593;
    wire N__60590;
    wire N__60587;
    wire N__60586;
    wire N__60583;
    wire N__60576;
    wire N__60573;
    wire N__60572;
    wire N__60571;
    wire N__60570;
    wire N__60567;
    wire N__60564;
    wire N__60561;
    wire N__60560;
    wire N__60557;
    wire N__60554;
    wire N__60551;
    wire N__60548;
    wire N__60547;
    wire N__60542;
    wire N__60539;
    wire N__60538;
    wire N__60537;
    wire N__60536;
    wire N__60533;
    wire N__60530;
    wire N__60527;
    wire N__60526;
    wire N__60523;
    wire N__60522;
    wire N__60521;
    wire N__60520;
    wire N__60517;
    wire N__60514;
    wire N__60511;
    wire N__60500;
    wire N__60495;
    wire N__60494;
    wire N__60491;
    wire N__60488;
    wire N__60485;
    wire N__60484;
    wire N__60481;
    wire N__60478;
    wire N__60475;
    wire N__60468;
    wire N__60465;
    wire N__60462;
    wire N__60459;
    wire N__60456;
    wire N__60455;
    wire N__60454;
    wire N__60453;
    wire N__60450;
    wire N__60449;
    wire N__60448;
    wire N__60447;
    wire N__60444;
    wire N__60441;
    wire N__60438;
    wire N__60433;
    wire N__60428;
    wire N__60425;
    wire N__60422;
    wire N__60415;
    wire N__60412;
    wire N__60409;
    wire N__60406;
    wire N__60401;
    wire N__60398;
    wire N__60395;
    wire N__60392;
    wire N__60389;
    wire N__60386;
    wire N__60383;
    wire N__60380;
    wire N__60377;
    wire N__60376;
    wire N__60375;
    wire N__60374;
    wire N__60373;
    wire N__60370;
    wire N__60367;
    wire N__60364;
    wire N__60359;
    wire N__60356;
    wire N__60349;
    wire N__60344;
    wire N__60335;
    wire N__60332;
    wire N__60329;
    wire N__60326;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60312;
    wire N__60309;
    wire N__60302;
    wire N__60299;
    wire N__60294;
    wire N__60291;
    wire N__60280;
    wire N__60277;
    wire N__60272;
    wire N__60269;
    wire N__60252;
    wire N__60249;
    wire N__60246;
    wire N__60243;
    wire N__60240;
    wire N__60237;
    wire N__60234;
    wire N__60231;
    wire N__60228;
    wire N__60225;
    wire N__60222;
    wire N__60219;
    wire N__60216;
    wire N__60213;
    wire N__60210;
    wire N__60207;
    wire N__60206;
    wire N__60203;
    wire N__60200;
    wire N__60197;
    wire N__60192;
    wire N__60189;
    wire N__60186;
    wire N__60183;
    wire N__60182;
    wire N__60179;
    wire N__60176;
    wire N__60173;
    wire N__60170;
    wire N__60167;
    wire N__60164;
    wire N__60159;
    wire N__60156;
    wire N__60153;
    wire N__60150;
    wire N__60147;
    wire N__60144;
    wire N__60143;
    wire N__60140;
    wire N__60137;
    wire N__60134;
    wire N__60131;
    wire N__60128;
    wire N__60125;
    wire N__60120;
    wire N__60117;
    wire N__60114;
    wire N__60111;
    wire N__60108;
    wire N__60105;
    wire N__60102;
    wire N__60101;
    wire N__60098;
    wire N__60095;
    wire N__60092;
    wire N__60089;
    wire N__60086;
    wire N__60083;
    wire N__60078;
    wire N__60075;
    wire N__60072;
    wire N__60069;
    wire N__60066;
    wire N__60063;
    wire N__60062;
    wire N__60059;
    wire N__60056;
    wire N__60053;
    wire N__60050;
    wire N__60047;
    wire N__60042;
    wire N__60039;
    wire N__60036;
    wire N__60033;
    wire N__60030;
    wire N__60027;
    wire N__60024;
    wire N__60021;
    wire N__60018;
    wire N__60015;
    wire N__60014;
    wire N__60011;
    wire N__60008;
    wire N__60003;
    wire N__60000;
    wire N__59997;
    wire N__59994;
    wire N__59991;
    wire N__59988;
    wire N__59985;
    wire N__59984;
    wire N__59981;
    wire N__59980;
    wire N__59977;
    wire N__59974;
    wire N__59971;
    wire N__59968;
    wire N__59965;
    wire N__59958;
    wire N__59957;
    wire N__59956;
    wire N__59953;
    wire N__59952;
    wire N__59951;
    wire N__59948;
    wire N__59947;
    wire N__59946;
    wire N__59943;
    wire N__59940;
    wire N__59937;
    wire N__59936;
    wire N__59935;
    wire N__59934;
    wire N__59933;
    wire N__59930;
    wire N__59927;
    wire N__59922;
    wire N__59919;
    wire N__59916;
    wire N__59913;
    wire N__59910;
    wire N__59907;
    wire N__59904;
    wire N__59901;
    wire N__59896;
    wire N__59877;
    wire N__59874;
    wire N__59871;
    wire N__59868;
    wire N__59867;
    wire N__59866;
    wire N__59863;
    wire N__59860;
    wire N__59855;
    wire N__59852;
    wire N__59849;
    wire N__59846;
    wire N__59843;
    wire N__59838;
    wire N__59837;
    wire N__59836;
    wire N__59833;
    wire N__59830;
    wire N__59825;
    wire N__59822;
    wire N__59819;
    wire N__59814;
    wire N__59811;
    wire N__59808;
    wire N__59805;
    wire N__59802;
    wire N__59799;
    wire N__59798;
    wire N__59797;
    wire N__59790;
    wire N__59787;
    wire N__59784;
    wire N__59783;
    wire N__59780;
    wire N__59777;
    wire N__59774;
    wire N__59771;
    wire N__59768;
    wire N__59765;
    wire N__59760;
    wire N__59757;
    wire N__59754;
    wire N__59751;
    wire N__59748;
    wire N__59745;
    wire N__59742;
    wire N__59739;
    wire N__59736;
    wire N__59733;
    wire N__59730;
    wire N__59727;
    wire N__59724;
    wire N__59721;
    wire N__59718;
    wire N__59715;
    wire N__59712;
    wire N__59711;
    wire N__59708;
    wire N__59705;
    wire N__59700;
    wire N__59697;
    wire N__59694;
    wire N__59693;
    wire N__59692;
    wire N__59685;
    wire N__59682;
    wire N__59679;
    wire N__59676;
    wire N__59673;
    wire N__59670;
    wire N__59667;
    wire N__59664;
    wire N__59663;
    wire N__59660;
    wire N__59657;
    wire N__59654;
    wire N__59651;
    wire N__59646;
    wire N__59643;
    wire N__59640;
    wire N__59639;
    wire N__59638;
    wire N__59635;
    wire N__59628;
    wire N__59625;
    wire N__59622;
    wire N__59621;
    wire N__59620;
    wire N__59617;
    wire N__59612;
    wire N__59607;
    wire N__59604;
    wire N__59603;
    wire N__59600;
    wire N__59597;
    wire N__59594;
    wire N__59589;
    wire N__59586;
    wire N__59583;
    wire N__59580;
    wire N__59577;
    wire N__59574;
    wire N__59571;
    wire N__59568;
    wire N__59565;
    wire N__59562;
    wire N__59559;
    wire N__59558;
    wire N__59555;
    wire N__59552;
    wire N__59547;
    wire N__59544;
    wire N__59541;
    wire N__59538;
    wire N__59537;
    wire N__59534;
    wire N__59531;
    wire N__59528;
    wire N__59525;
    wire N__59522;
    wire N__59519;
    wire N__59516;
    wire N__59513;
    wire N__59508;
    wire N__59507;
    wire N__59506;
    wire N__59503;
    wire N__59498;
    wire N__59493;
    wire N__59492;
    wire N__59491;
    wire N__59488;
    wire N__59485;
    wire N__59480;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59468;
    wire N__59467;
    wire N__59466;
    wire N__59463;
    wire N__59456;
    wire N__59451;
    wire N__59448;
    wire N__59445;
    wire N__59442;
    wire N__59439;
    wire N__59436;
    wire N__59433;
    wire N__59430;
    wire N__59427;
    wire N__59426;
    wire N__59425;
    wire N__59424;
    wire N__59423;
    wire N__59422;
    wire N__59419;
    wire N__59416;
    wire N__59413;
    wire N__59410;
    wire N__59407;
    wire N__59404;
    wire N__59403;
    wire N__59400;
    wire N__59397;
    wire N__59394;
    wire N__59391;
    wire N__59386;
    wire N__59383;
    wire N__59378;
    wire N__59377;
    wire N__59368;
    wire N__59367;
    wire N__59364;
    wire N__59363;
    wire N__59360;
    wire N__59357;
    wire N__59354;
    wire N__59351;
    wire N__59348;
    wire N__59347;
    wire N__59346;
    wire N__59345;
    wire N__59342;
    wire N__59337;
    wire N__59336;
    wire N__59331;
    wire N__59328;
    wire N__59327;
    wire N__59324;
    wire N__59321;
    wire N__59318;
    wire N__59315;
    wire N__59312;
    wire N__59309;
    wire N__59306;
    wire N__59303;
    wire N__59298;
    wire N__59295;
    wire N__59292;
    wire N__59289;
    wire N__59286;
    wire N__59283;
    wire N__59278;
    wire N__59275;
    wire N__59270;
    wire N__59267;
    wire N__59262;
    wire N__59259;
    wire N__59256;
    wire N__59253;
    wire N__59244;
    wire N__59241;
    wire N__59240;
    wire N__59239;
    wire N__59236;
    wire N__59233;
    wire N__59230;
    wire N__59225;
    wire N__59224;
    wire N__59221;
    wire N__59218;
    wire N__59215;
    wire N__59212;
    wire N__59207;
    wire N__59202;
    wire N__59201;
    wire N__59200;
    wire N__59199;
    wire N__59198;
    wire N__59195;
    wire N__59190;
    wire N__59187;
    wire N__59184;
    wire N__59179;
    wire N__59172;
    wire N__59169;
    wire N__59166;
    wire N__59163;
    wire N__59160;
    wire N__59159;
    wire N__59156;
    wire N__59153;
    wire N__59152;
    wire N__59149;
    wire N__59146;
    wire N__59143;
    wire N__59140;
    wire N__59137;
    wire N__59130;
    wire N__59129;
    wire N__59128;
    wire N__59125;
    wire N__59122;
    wire N__59119;
    wire N__59116;
    wire N__59113;
    wire N__59110;
    wire N__59107;
    wire N__59104;
    wire N__59097;
    wire N__59094;
    wire N__59091;
    wire N__59088;
    wire N__59085;
    wire N__59084;
    wire N__59083;
    wire N__59082;
    wire N__59079;
    wire N__59074;
    wire N__59071;
    wire N__59064;
    wire N__59063;
    wire N__59060;
    wire N__59057;
    wire N__59056;
    wire N__59053;
    wire N__59050;
    wire N__59047;
    wire N__59044;
    wire N__59041;
    wire N__59034;
    wire N__59031;
    wire N__59028;
    wire N__59025;
    wire N__59022;
    wire N__59021;
    wire N__59018;
    wire N__59015;
    wire N__59010;
    wire N__59007;
    wire N__59004;
    wire N__59001;
    wire N__58998;
    wire N__58995;
    wire N__58992;
    wire N__58989;
    wire N__58988;
    wire N__58987;
    wire N__58986;
    wire N__58983;
    wire N__58980;
    wire N__58975;
    wire N__58970;
    wire N__58965;
    wire N__58962;
    wire N__58959;
    wire N__58956;
    wire N__58953;
    wire N__58950;
    wire N__58949;
    wire N__58946;
    wire N__58943;
    wire N__58938;
    wire N__58935;
    wire N__58932;
    wire N__58929;
    wire N__58926;
    wire N__58923;
    wire N__58920;
    wire N__58917;
    wire N__58914;
    wire N__58913;
    wire N__58912;
    wire N__58911;
    wire N__58908;
    wire N__58903;
    wire N__58900;
    wire N__58893;
    wire N__58890;
    wire N__58887;
    wire N__58884;
    wire N__58881;
    wire N__58880;
    wire N__58879;
    wire N__58876;
    wire N__58871;
    wire N__58866;
    wire N__58865;
    wire N__58864;
    wire N__58863;
    wire N__58860;
    wire N__58857;
    wire N__58852;
    wire N__58845;
    wire N__58842;
    wire N__58839;
    wire N__58836;
    wire N__58833;
    wire N__58830;
    wire N__58827;
    wire N__58824;
    wire N__58821;
    wire N__58818;
    wire N__58815;
    wire N__58812;
    wire N__58809;
    wire N__58806;
    wire N__58803;
    wire N__58800;
    wire N__58797;
    wire N__58794;
    wire N__58791;
    wire N__58788;
    wire N__58785;
    wire N__58782;
    wire N__58779;
    wire N__58776;
    wire N__58773;
    wire N__58772;
    wire N__58769;
    wire N__58768;
    wire N__58767;
    wire N__58764;
    wire N__58761;
    wire N__58756;
    wire N__58755;
    wire N__58748;
    wire N__58745;
    wire N__58740;
    wire N__58737;
    wire N__58734;
    wire N__58731;
    wire N__58728;
    wire N__58725;
    wire N__58722;
    wire N__58719;
    wire N__58716;
    wire N__58713;
    wire N__58710;
    wire N__58707;
    wire N__58704;
    wire N__58701;
    wire N__58698;
    wire N__58695;
    wire N__58692;
    wire N__58689;
    wire N__58686;
    wire N__58683;
    wire N__58680;
    wire N__58679;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58659;
    wire N__58658;
    wire N__58655;
    wire N__58652;
    wire N__58649;
    wire N__58646;
    wire N__58643;
    wire N__58640;
    wire N__58635;
    wire N__58632;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58620;
    wire N__58617;
    wire N__58614;
    wire N__58611;
    wire N__58610;
    wire N__58605;
    wire N__58602;
    wire N__58599;
    wire N__58596;
    wire N__58593;
    wire N__58590;
    wire N__58587;
    wire N__58584;
    wire N__58581;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58569;
    wire N__58566;
    wire N__58563;
    wire N__58560;
    wire N__58559;
    wire N__58554;
    wire N__58551;
    wire N__58550;
    wire N__58547;
    wire N__58544;
    wire N__58541;
    wire N__58538;
    wire N__58535;
    wire N__58532;
    wire N__58529;
    wire N__58526;
    wire N__58521;
    wire N__58518;
    wire N__58517;
    wire N__58514;
    wire N__58513;
    wire N__58512;
    wire N__58511;
    wire N__58510;
    wire N__58509;
    wire N__58508;
    wire N__58507;
    wire N__58506;
    wire N__58505;
    wire N__58504;
    wire N__58499;
    wire N__58496;
    wire N__58495;
    wire N__58492;
    wire N__58489;
    wire N__58486;
    wire N__58485;
    wire N__58484;
    wire N__58483;
    wire N__58480;
    wire N__58477;
    wire N__58474;
    wire N__58471;
    wire N__58470;
    wire N__58467;
    wire N__58464;
    wire N__58461;
    wire N__58458;
    wire N__58449;
    wire N__58446;
    wire N__58443;
    wire N__58434;
    wire N__58425;
    wire N__58422;
    wire N__58419;
    wire N__58416;
    wire N__58411;
    wire N__58410;
    wire N__58405;
    wire N__58402;
    wire N__58401;
    wire N__58398;
    wire N__58393;
    wire N__58390;
    wire N__58389;
    wire N__58386;
    wire N__58383;
    wire N__58380;
    wire N__58373;
    wire N__58370;
    wire N__58367;
    wire N__58362;
    wire N__58359;
    wire N__58350;
    wire N__58349;
    wire N__58348;
    wire N__58347;
    wire N__58346;
    wire N__58343;
    wire N__58342;
    wire N__58341;
    wire N__58340;
    wire N__58339;
    wire N__58338;
    wire N__58335;
    wire N__58328;
    wire N__58325;
    wire N__58322;
    wire N__58313;
    wire N__58312;
    wire N__58311;
    wire N__58306;
    wire N__58305;
    wire N__58304;
    wire N__58303;
    wire N__58302;
    wire N__58301;
    wire N__58298;
    wire N__58295;
    wire N__58292;
    wire N__58287;
    wire N__58284;
    wire N__58281;
    wire N__58280;
    wire N__58277;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58269;
    wire N__58266;
    wire N__58265;
    wire N__58264;
    wire N__58261;
    wire N__58252;
    wire N__58249;
    wire N__58246;
    wire N__58243;
    wire N__58228;
    wire N__58225;
    wire N__58220;
    wire N__58217;
    wire N__58206;
    wire N__58203;
    wire N__58200;
    wire N__58197;
    wire N__58194;
    wire N__58193;
    wire N__58190;
    wire N__58187;
    wire N__58182;
    wire N__58179;
    wire N__58176;
    wire N__58173;
    wire N__58170;
    wire N__58167;
    wire N__58166;
    wire N__58163;
    wire N__58158;
    wire N__58155;
    wire N__58152;
    wire N__58149;
    wire N__58148;
    wire N__58147;
    wire N__58146;
    wire N__58143;
    wire N__58142;
    wire N__58139;
    wire N__58138;
    wire N__58137;
    wire N__58136;
    wire N__58135;
    wire N__58134;
    wire N__58123;
    wire N__58120;
    wire N__58119;
    wire N__58116;
    wire N__58115;
    wire N__58112;
    wire N__58111;
    wire N__58108;
    wire N__58107;
    wire N__58106;
    wire N__58103;
    wire N__58102;
    wire N__58099;
    wire N__58082;
    wire N__58075;
    wire N__58068;
    wire N__58065;
    wire N__58064;
    wire N__58059;
    wire N__58056;
    wire N__58055;
    wire N__58052;
    wire N__58047;
    wire N__58044;
    wire N__58041;
    wire N__58038;
    wire N__58037;
    wire N__58036;
    wire N__58033;
    wire N__58030;
    wire N__58029;
    wire N__58026;
    wire N__58023;
    wire N__58020;
    wire N__58015;
    wire N__58010;
    wire N__58005;
    wire N__58004;
    wire N__58001;
    wire N__57998;
    wire N__57997;
    wire N__57996;
    wire N__57995;
    wire N__57992;
    wire N__57991;
    wire N__57988;
    wire N__57985;
    wire N__57980;
    wire N__57979;
    wire N__57978;
    wire N__57975;
    wire N__57972;
    wire N__57969;
    wire N__57964;
    wire N__57959;
    wire N__57956;
    wire N__57953;
    wire N__57948;
    wire N__57945;
    wire N__57940;
    wire N__57937;
    wire N__57934;
    wire N__57927;
    wire N__57924;
    wire N__57921;
    wire N__57918;
    wire N__57915;
    wire N__57912;
    wire N__57909;
    wire N__57906;
    wire N__57903;
    wire N__57900;
    wire N__57897;
    wire N__57894;
    wire N__57891;
    wire N__57888;
    wire N__57885;
    wire N__57882;
    wire N__57879;
    wire N__57876;
    wire N__57873;
    wire N__57870;
    wire N__57867;
    wire N__57864;
    wire N__57861;
    wire N__57858;
    wire N__57855;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57843;
    wire N__57840;
    wire N__57837;
    wire N__57834;
    wire N__57831;
    wire N__57828;
    wire N__57825;
    wire N__57822;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57804;
    wire N__57801;
    wire N__57798;
    wire N__57795;
    wire N__57792;
    wire N__57789;
    wire N__57786;
    wire N__57783;
    wire N__57780;
    wire N__57777;
    wire N__57774;
    wire N__57771;
    wire N__57768;
    wire N__57765;
    wire N__57762;
    wire N__57759;
    wire N__57756;
    wire N__57753;
    wire N__57750;
    wire N__57747;
    wire N__57744;
    wire N__57741;
    wire N__57738;
    wire N__57735;
    wire N__57732;
    wire N__57729;
    wire N__57726;
    wire N__57723;
    wire N__57720;
    wire N__57717;
    wire N__57714;
    wire N__57711;
    wire N__57708;
    wire N__57705;
    wire N__57702;
    wire N__57699;
    wire N__57696;
    wire N__57693;
    wire N__57690;
    wire N__57687;
    wire N__57684;
    wire N__57681;
    wire N__57680;
    wire N__57677;
    wire N__57674;
    wire N__57673;
    wire N__57668;
    wire N__57665;
    wire N__57662;
    wire N__57657;
    wire N__57656;
    wire N__57653;
    wire N__57650;
    wire N__57647;
    wire N__57644;
    wire N__57643;
    wire N__57638;
    wire N__57635;
    wire N__57632;
    wire N__57627;
    wire N__57626;
    wire N__57623;
    wire N__57620;
    wire N__57617;
    wire N__57614;
    wire N__57611;
    wire N__57610;
    wire N__57605;
    wire N__57602;
    wire N__57599;
    wire N__57594;
    wire N__57593;
    wire N__57590;
    wire N__57587;
    wire N__57584;
    wire N__57579;
    wire N__57578;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57561;
    wire N__57558;
    wire N__57557;
    wire N__57556;
    wire N__57553;
    wire N__57550;
    wire N__57547;
    wire N__57540;
    wire N__57537;
    wire N__57536;
    wire N__57533;
    wire N__57530;
    wire N__57525;
    wire N__57522;
    wire N__57519;
    wire N__57516;
    wire N__57513;
    wire N__57510;
    wire N__57507;
    wire N__57504;
    wire N__57501;
    wire N__57498;
    wire N__57495;
    wire N__57492;
    wire N__57489;
    wire N__57486;
    wire N__57483;
    wire N__57482;
    wire N__57479;
    wire N__57476;
    wire N__57473;
    wire N__57470;
    wire N__57465;
    wire N__57462;
    wire N__57459;
    wire N__57456;
    wire N__57453;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57441;
    wire N__57440;
    wire N__57437;
    wire N__57434;
    wire N__57429;
    wire N__57426;
    wire N__57423;
    wire N__57420;
    wire N__57417;
    wire N__57414;
    wire N__57413;
    wire N__57410;
    wire N__57407;
    wire N__57404;
    wire N__57401;
    wire N__57398;
    wire N__57395;
    wire N__57390;
    wire N__57389;
    wire N__57386;
    wire N__57385;
    wire N__57380;
    wire N__57377;
    wire N__57374;
    wire N__57369;
    wire N__57366;
    wire N__57363;
    wire N__57360;
    wire N__57357;
    wire N__57354;
    wire N__57351;
    wire N__57350;
    wire N__57349;
    wire N__57342;
    wire N__57339;
    wire N__57336;
    wire N__57335;
    wire N__57332;
    wire N__57329;
    wire N__57326;
    wire N__57323;
    wire N__57318;
    wire N__57315;
    wire N__57312;
    wire N__57309;
    wire N__57306;
    wire N__57305;
    wire N__57304;
    wire N__57301;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57287;
    wire N__57284;
    wire N__57281;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57252;
    wire N__57251;
    wire N__57250;
    wire N__57247;
    wire N__57240;
    wire N__57237;
    wire N__57236;
    wire N__57235;
    wire N__57232;
    wire N__57227;
    wire N__57224;
    wire N__57219;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57204;
    wire N__57203;
    wire N__57202;
    wire N__57199;
    wire N__57194;
    wire N__57189;
    wire N__57186;
    wire N__57185;
    wire N__57182;
    wire N__57179;
    wire N__57176;
    wire N__57173;
    wire N__57168;
    wire N__57165;
    wire N__57162;
    wire N__57159;
    wire N__57156;
    wire N__57155;
    wire N__57154;
    wire N__57151;
    wire N__57148;
    wire N__57145;
    wire N__57142;
    wire N__57139;
    wire N__57132;
    wire N__57129;
    wire N__57128;
    wire N__57125;
    wire N__57120;
    wire N__57117;
    wire N__57114;
    wire N__57111;
    wire N__57108;
    wire N__57107;
    wire N__57104;
    wire N__57101;
    wire N__57100;
    wire N__57097;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57078;
    wire N__57075;
    wire N__57072;
    wire N__57069;
    wire N__57066;
    wire N__57063;
    wire N__57060;
    wire N__57059;
    wire N__57056;
    wire N__57053;
    wire N__57052;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57038;
    wire N__57033;
    wire N__57030;
    wire N__57027;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57015;
    wire N__57012;
    wire N__57009;
    wire N__57006;
    wire N__57005;
    wire N__57002;
    wire N__57001;
    wire N__56996;
    wire N__56993;
    wire N__56990;
    wire N__56987;
    wire N__56984;
    wire N__56979;
    wire N__56976;
    wire N__56973;
    wire N__56970;
    wire N__56967;
    wire N__56964;
    wire N__56963;
    wire N__56962;
    wire N__56955;
    wire N__56952;
    wire N__56951;
    wire N__56948;
    wire N__56945;
    wire N__56944;
    wire N__56941;
    wire N__56938;
    wire N__56935;
    wire N__56932;
    wire N__56925;
    wire N__56924;
    wire N__56921;
    wire N__56918;
    wire N__56915;
    wire N__56914;
    wire N__56911;
    wire N__56908;
    wire N__56905;
    wire N__56902;
    wire N__56899;
    wire N__56892;
    wire N__56889;
    wire N__56886;
    wire N__56883;
    wire N__56882;
    wire N__56879;
    wire N__56876;
    wire N__56871;
    wire N__56868;
    wire N__56865;
    wire N__56864;
    wire N__56861;
    wire N__56858;
    wire N__56853;
    wire N__56850;
    wire N__56849;
    wire N__56848;
    wire N__56841;
    wire N__56838;
    wire N__56835;
    wire N__56832;
    wire N__56829;
    wire N__56826;
    wire N__56823;
    wire N__56820;
    wire N__56817;
    wire N__56814;
    wire N__56811;
    wire N__56808;
    wire N__56807;
    wire N__56804;
    wire N__56803;
    wire N__56802;
    wire N__56799;
    wire N__56798;
    wire N__56795;
    wire N__56790;
    wire N__56787;
    wire N__56784;
    wire N__56779;
    wire N__56772;
    wire N__56769;
    wire N__56766;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56754;
    wire N__56751;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56739;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56727;
    wire N__56724;
    wire N__56721;
    wire N__56720;
    wire N__56717;
    wire N__56714;
    wire N__56713;
    wire N__56712;
    wire N__56709;
    wire N__56706;
    wire N__56701;
    wire N__56698;
    wire N__56695;
    wire N__56692;
    wire N__56685;
    wire N__56684;
    wire N__56683;
    wire N__56680;
    wire N__56677;
    wire N__56674;
    wire N__56667;
    wire N__56664;
    wire N__56661;
    wire N__56658;
    wire N__56655;
    wire N__56652;
    wire N__56649;
    wire N__56646;
    wire N__56643;
    wire N__56640;
    wire N__56637;
    wire N__56634;
    wire N__56631;
    wire N__56628;
    wire N__56625;
    wire N__56624;
    wire N__56623;
    wire N__56622;
    wire N__56619;
    wire N__56612;
    wire N__56607;
    wire N__56606;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56596;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56580;
    wire N__56577;
    wire N__56574;
    wire N__56571;
    wire N__56568;
    wire N__56565;
    wire N__56562;
    wire N__56559;
    wire N__56556;
    wire N__56553;
    wire N__56550;
    wire N__56547;
    wire N__56544;
    wire N__56541;
    wire N__56538;
    wire N__56535;
    wire N__56534;
    wire N__56531;
    wire N__56528;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56520;
    wire N__56519;
    wire N__56516;
    wire N__56515;
    wire N__56514;
    wire N__56513;
    wire N__56512;
    wire N__56509;
    wire N__56506;
    wire N__56505;
    wire N__56504;
    wire N__56501;
    wire N__56498;
    wire N__56497;
    wire N__56496;
    wire N__56495;
    wire N__56492;
    wire N__56489;
    wire N__56482;
    wire N__56481;
    wire N__56480;
    wire N__56477;
    wire N__56474;
    wire N__56473;
    wire N__56468;
    wire N__56467;
    wire N__56462;
    wire N__56455;
    wire N__56452;
    wire N__56447;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56437;
    wire N__56434;
    wire N__56431;
    wire N__56428;
    wire N__56425;
    wire N__56420;
    wire N__56413;
    wire N__56408;
    wire N__56403;
    wire N__56388;
    wire N__56385;
    wire N__56382;
    wire N__56379;
    wire N__56378;
    wire N__56377;
    wire N__56374;
    wire N__56371;
    wire N__56368;
    wire N__56363;
    wire N__56358;
    wire N__56355;
    wire N__56352;
    wire N__56349;
    wire N__56346;
    wire N__56343;
    wire N__56340;
    wire N__56337;
    wire N__56334;
    wire N__56331;
    wire N__56328;
    wire N__56325;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56315;
    wire N__56312;
    wire N__56309;
    wire N__56306;
    wire N__56303;
    wire N__56302;
    wire N__56299;
    wire N__56296;
    wire N__56293;
    wire N__56292;
    wire N__56289;
    wire N__56286;
    wire N__56281;
    wire N__56274;
    wire N__56271;
    wire N__56268;
    wire N__56265;
    wire N__56264;
    wire N__56263;
    wire N__56260;
    wire N__56257;
    wire N__56254;
    wire N__56251;
    wire N__56248;
    wire N__56245;
    wire N__56244;
    wire N__56243;
    wire N__56242;
    wire N__56241;
    wire N__56236;
    wire N__56233;
    wire N__56224;
    wire N__56217;
    wire N__56214;
    wire N__56211;
    wire N__56208;
    wire N__56207;
    wire N__56204;
    wire N__56203;
    wire N__56202;
    wire N__56199;
    wire N__56192;
    wire N__56187;
    wire N__56186;
    wire N__56185;
    wire N__56184;
    wire N__56181;
    wire N__56176;
    wire N__56173;
    wire N__56166;
    wire N__56163;
    wire N__56162;
    wire N__56159;
    wire N__56158;
    wire N__56157;
    wire N__56156;
    wire N__56153;
    wire N__56150;
    wire N__56147;
    wire N__56144;
    wire N__56141;
    wire N__56138;
    wire N__56135;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56123;
    wire N__56120;
    wire N__56117;
    wire N__56112;
    wire N__56103;
    wire N__56102;
    wire N__56099;
    wire N__56096;
    wire N__56093;
    wire N__56090;
    wire N__56089;
    wire N__56086;
    wire N__56083;
    wire N__56082;
    wire N__56079;
    wire N__56078;
    wire N__56075;
    wire N__56072;
    wire N__56069;
    wire N__56066;
    wire N__56063;
    wire N__56062;
    wire N__56059;
    wire N__56054;
    wire N__56049;
    wire N__56046;
    wire N__56041;
    wire N__56034;
    wire N__56033;
    wire N__56030;
    wire N__56029;
    wire N__56028;
    wire N__56025;
    wire N__56022;
    wire N__56019;
    wire N__56016;
    wire N__56007;
    wire N__56004;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55994;
    wire N__55991;
    wire N__55988;
    wire N__55985;
    wire N__55982;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55968;
    wire N__55965;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55953;
    wire N__55950;
    wire N__55947;
    wire N__55944;
    wire N__55941;
    wire N__55938;
    wire N__55935;
    wire N__55932;
    wire N__55929;
    wire N__55926;
    wire N__55923;
    wire N__55920;
    wire N__55917;
    wire N__55914;
    wire N__55911;
    wire N__55908;
    wire N__55907;
    wire N__55904;
    wire N__55903;
    wire N__55900;
    wire N__55895;
    wire N__55892;
    wire N__55887;
    wire N__55886;
    wire N__55881;
    wire N__55878;
    wire N__55875;
    wire N__55872;
    wire N__55869;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55857;
    wire N__55854;
    wire N__55853;
    wire N__55850;
    wire N__55847;
    wire N__55844;
    wire N__55839;
    wire N__55836;
    wire N__55833;
    wire N__55830;
    wire N__55829;
    wire N__55826;
    wire N__55823;
    wire N__55822;
    wire N__55819;
    wire N__55818;
    wire N__55815;
    wire N__55812;
    wire N__55809;
    wire N__55806;
    wire N__55805;
    wire N__55804;
    wire N__55801;
    wire N__55798;
    wire N__55797;
    wire N__55792;
    wire N__55789;
    wire N__55788;
    wire N__55785;
    wire N__55784;
    wire N__55781;
    wire N__55778;
    wire N__55775;
    wire N__55772;
    wire N__55767;
    wire N__55762;
    wire N__55749;
    wire N__55746;
    wire N__55745;
    wire N__55742;
    wire N__55741;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55731;
    wire N__55728;
    wire N__55727;
    wire N__55724;
    wire N__55723;
    wire N__55720;
    wire N__55717;
    wire N__55714;
    wire N__55711;
    wire N__55710;
    wire N__55707;
    wire N__55704;
    wire N__55701;
    wire N__55696;
    wire N__55691;
    wire N__55688;
    wire N__55683;
    wire N__55674;
    wire N__55671;
    wire N__55668;
    wire N__55665;
    wire N__55662;
    wire N__55661;
    wire N__55660;
    wire N__55653;
    wire N__55650;
    wire N__55649;
    wire N__55644;
    wire N__55641;
    wire N__55638;
    wire N__55635;
    wire N__55632;
    wire N__55629;
    wire N__55626;
    wire N__55623;
    wire N__55620;
    wire N__55617;
    wire N__55616;
    wire N__55613;
    wire N__55610;
    wire N__55607;
    wire N__55604;
    wire N__55601;
    wire N__55596;
    wire N__55593;
    wire N__55592;
    wire N__55589;
    wire N__55584;
    wire N__55583;
    wire N__55580;
    wire N__55577;
    wire N__55574;
    wire N__55571;
    wire N__55568;
    wire N__55565;
    wire N__55562;
    wire N__55559;
    wire N__55554;
    wire N__55551;
    wire N__55550;
    wire N__55547;
    wire N__55544;
    wire N__55539;
    wire N__55536;
    wire N__55533;
    wire N__55532;
    wire N__55529;
    wire N__55526;
    wire N__55523;
    wire N__55518;
    wire N__55515;
    wire N__55514;
    wire N__55511;
    wire N__55508;
    wire N__55507;
    wire N__55506;
    wire N__55501;
    wire N__55498;
    wire N__55495;
    wire N__55488;
    wire N__55485;
    wire N__55482;
    wire N__55479;
    wire N__55476;
    wire N__55473;
    wire N__55470;
    wire N__55467;
    wire N__55466;
    wire N__55463;
    wire N__55460;
    wire N__55457;
    wire N__55452;
    wire N__55449;
    wire N__55446;
    wire N__55443;
    wire N__55440;
    wire N__55437;
    wire N__55436;
    wire N__55433;
    wire N__55430;
    wire N__55429;
    wire N__55428;
    wire N__55423;
    wire N__55418;
    wire N__55413;
    wire N__55410;
    wire N__55407;
    wire N__55404;
    wire N__55401;
    wire N__55398;
    wire N__55395;
    wire N__55394;
    wire N__55391;
    wire N__55388;
    wire N__55387;
    wire N__55382;
    wire N__55379;
    wire N__55374;
    wire N__55373;
    wire N__55370;
    wire N__55367;
    wire N__55366;
    wire N__55361;
    wire N__55358;
    wire N__55353;
    wire N__55350;
    wire N__55347;
    wire N__55344;
    wire N__55343;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55330;
    wire N__55323;
    wire N__55320;
    wire N__55317;
    wire N__55314;
    wire N__55311;
    wire N__55308;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55298;
    wire N__55297;
    wire N__55294;
    wire N__55289;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55275;
    wire N__55272;
    wire N__55269;
    wire N__55268;
    wire N__55267;
    wire N__55264;
    wire N__55259;
    wire N__55254;
    wire N__55253;
    wire N__55250;
    wire N__55247;
    wire N__55242;
    wire N__55241;
    wire N__55238;
    wire N__55235;
    wire N__55230;
    wire N__55227;
    wire N__55226;
    wire N__55223;
    wire N__55220;
    wire N__55215;
    wire N__55212;
    wire N__55209;
    wire N__55208;
    wire N__55207;
    wire N__55204;
    wire N__55199;
    wire N__55194;
    wire N__55191;
    wire N__55190;
    wire N__55185;
    wire N__55182;
    wire N__55181;
    wire N__55176;
    wire N__55173;
    wire N__55172;
    wire N__55167;
    wire N__55164;
    wire N__55163;
    wire N__55162;
    wire N__55161;
    wire N__55160;
    wire N__55159;
    wire N__55146;
    wire N__55143;
    wire N__55142;
    wire N__55141;
    wire N__55140;
    wire N__55139;
    wire N__55128;
    wire N__55127;
    wire N__55126;
    wire N__55125;
    wire N__55124;
    wire N__55123;
    wire N__55122;
    wire N__55121;
    wire N__55120;
    wire N__55117;
    wire N__55110;
    wire N__55099;
    wire N__55092;
    wire N__55091;
    wire N__55088;
    wire N__55085;
    wire N__55084;
    wire N__55081;
    wire N__55078;
    wire N__55075;
    wire N__55072;
    wire N__55067;
    wire N__55062;
    wire N__55059;
    wire N__55056;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55044;
    wire N__55041;
    wire N__55038;
    wire N__55035;
    wire N__55032;
    wire N__55029;
    wire N__55028;
    wire N__55023;
    wire N__55020;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55007;
    wire N__55004;
    wire N__55003;
    wire N__55000;
    wire N__54999;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54987;
    wire N__54984;
    wire N__54983;
    wire N__54982;
    wire N__54979;
    wire N__54974;
    wire N__54973;
    wire N__54972;
    wire N__54969;
    wire N__54968;
    wire N__54967;
    wire N__54964;
    wire N__54961;
    wire N__54958;
    wire N__54955;
    wire N__54952;
    wire N__54949;
    wire N__54946;
    wire N__54941;
    wire N__54938;
    wire N__54933;
    wire N__54928;
    wire N__54925;
    wire N__54922;
    wire N__54919;
    wire N__54912;
    wire N__54909;
    wire N__54904;
    wire N__54901;
    wire N__54900;
    wire N__54895;
    wire N__54892;
    wire N__54889;
    wire N__54882;
    wire N__54879;
    wire N__54876;
    wire N__54873;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54865;
    wire N__54860;
    wire N__54855;
    wire N__54852;
    wire N__54849;
    wire N__54848;
    wire N__54847;
    wire N__54844;
    wire N__54839;
    wire N__54834;
    wire N__54831;
    wire N__54830;
    wire N__54827;
    wire N__54826;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54814;
    wire N__54807;
    wire N__54806;
    wire N__54801;
    wire N__54798;
    wire N__54795;
    wire N__54792;
    wire N__54791;
    wire N__54788;
    wire N__54785;
    wire N__54782;
    wire N__54777;
    wire N__54776;
    wire N__54771;
    wire N__54768;
    wire N__54765;
    wire N__54762;
    wire N__54759;
    wire N__54756;
    wire N__54753;
    wire N__54750;
    wire N__54747;
    wire N__54746;
    wire N__54745;
    wire N__54738;
    wire N__54735;
    wire N__54732;
    wire N__54729;
    wire N__54726;
    wire N__54723;
    wire N__54720;
    wire N__54719;
    wire N__54716;
    wire N__54713;
    wire N__54708;
    wire N__54705;
    wire N__54704;
    wire N__54703;
    wire N__54700;
    wire N__54693;
    wire N__54690;
    wire N__54687;
    wire N__54686;
    wire N__54683;
    wire N__54680;
    wire N__54675;
    wire N__54672;
    wire N__54669;
    wire N__54666;
    wire N__54663;
    wire N__54660;
    wire N__54657;
    wire N__54654;
    wire N__54653;
    wire N__54652;
    wire N__54649;
    wire N__54642;
    wire N__54639;
    wire N__54636;
    wire N__54633;
    wire N__54632;
    wire N__54631;
    wire N__54628;
    wire N__54625;
    wire N__54622;
    wire N__54619;
    wire N__54616;
    wire N__54609;
    wire N__54606;
    wire N__54603;
    wire N__54600;
    wire N__54597;
    wire N__54594;
    wire N__54591;
    wire N__54588;
    wire N__54587;
    wire N__54586;
    wire N__54583;
    wire N__54580;
    wire N__54577;
    wire N__54574;
    wire N__54567;
    wire N__54564;
    wire N__54561;
    wire N__54558;
    wire N__54557;
    wire N__54554;
    wire N__54553;
    wire N__54550;
    wire N__54547;
    wire N__54542;
    wire N__54537;
    wire N__54534;
    wire N__54533;
    wire N__54530;
    wire N__54529;
    wire N__54526;
    wire N__54523;
    wire N__54520;
    wire N__54513;
    wire N__54510;
    wire N__54507;
    wire N__54504;
    wire N__54501;
    wire N__54498;
    wire N__54495;
    wire N__54492;
    wire N__54489;
    wire N__54486;
    wire N__54483;
    wire N__54480;
    wire N__54479;
    wire N__54478;
    wire N__54471;
    wire N__54468;
    wire N__54465;
    wire N__54462;
    wire N__54459;
    wire N__54456;
    wire N__54453;
    wire N__54452;
    wire N__54449;
    wire N__54446;
    wire N__54441;
    wire N__54438;
    wire N__54437;
    wire N__54436;
    wire N__54433;
    wire N__54426;
    wire N__54423;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54408;
    wire N__54407;
    wire N__54404;
    wire N__54403;
    wire N__54400;
    wire N__54397;
    wire N__54394;
    wire N__54391;
    wire N__54386;
    wire N__54381;
    wire N__54380;
    wire N__54379;
    wire N__54376;
    wire N__54369;
    wire N__54366;
    wire N__54363;
    wire N__54360;
    wire N__54357;
    wire N__54354;
    wire N__54351;
    wire N__54350;
    wire N__54345;
    wire N__54342;
    wire N__54341;
    wire N__54338;
    wire N__54335;
    wire N__54332;
    wire N__54329;
    wire N__54326;
    wire N__54323;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54305;
    wire N__54300;
    wire N__54297;
    wire N__54294;
    wire N__54291;
    wire N__54288;
    wire N__54285;
    wire N__54282;
    wire N__54279;
    wire N__54276;
    wire N__54273;
    wire N__54270;
    wire N__54267;
    wire N__54264;
    wire N__54261;
    wire N__54258;
    wire N__54255;
    wire N__54252;
    wire N__54249;
    wire N__54246;
    wire N__54245;
    wire N__54244;
    wire N__54241;
    wire N__54238;
    wire N__54235;
    wire N__54232;
    wire N__54225;
    wire N__54222;
    wire N__54219;
    wire N__54216;
    wire N__54213;
    wire N__54210;
    wire N__54209;
    wire N__54208;
    wire N__54205;
    wire N__54202;
    wire N__54199;
    wire N__54196;
    wire N__54189;
    wire N__54188;
    wire N__54187;
    wire N__54184;
    wire N__54181;
    wire N__54178;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54162;
    wire N__54161;
    wire N__54160;
    wire N__54157;
    wire N__54154;
    wire N__54151;
    wire N__54148;
    wire N__54145;
    wire N__54142;
    wire N__54135;
    wire N__54132;
    wire N__54129;
    wire N__54126;
    wire N__54123;
    wire N__54120;
    wire N__54117;
    wire N__54114;
    wire N__54111;
    wire N__54108;
    wire N__54107;
    wire N__54104;
    wire N__54103;
    wire N__54100;
    wire N__54097;
    wire N__54094;
    wire N__54091;
    wire N__54088;
    wire N__54081;
    wire N__54078;
    wire N__54075;
    wire N__54072;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54060;
    wire N__54057;
    wire N__54054;
    wire N__54053;
    wire N__54050;
    wire N__54047;
    wire N__54042;
    wire N__54041;
    wire N__54038;
    wire N__54035;
    wire N__54030;
    wire N__54027;
    wire N__54026;
    wire N__54025;
    wire N__54022;
    wire N__54019;
    wire N__54016;
    wire N__54013;
    wire N__54006;
    wire N__54005;
    wire N__54004;
    wire N__54001;
    wire N__53998;
    wire N__53995;
    wire N__53992;
    wire N__53989;
    wire N__53982;
    wire N__53979;
    wire N__53976;
    wire N__53975;
    wire N__53974;
    wire N__53971;
    wire N__53968;
    wire N__53965;
    wire N__53962;
    wire N__53955;
    wire N__53952;
    wire N__53949;
    wire N__53948;
    wire N__53947;
    wire N__53944;
    wire N__53941;
    wire N__53938;
    wire N__53935;
    wire N__53928;
    wire N__53925;
    wire N__53922;
    wire N__53919;
    wire N__53916;
    wire N__53913;
    wire N__53912;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53899;
    wire N__53892;
    wire N__53889;
    wire N__53886;
    wire N__53885;
    wire N__53882;
    wire N__53879;
    wire N__53876;
    wire N__53873;
    wire N__53872;
    wire N__53867;
    wire N__53866;
    wire N__53865;
    wire N__53864;
    wire N__53861;
    wire N__53858;
    wire N__53855;
    wire N__53852;
    wire N__53849;
    wire N__53846;
    wire N__53835;
    wire N__53832;
    wire N__53831;
    wire N__53828;
    wire N__53825;
    wire N__53824;
    wire N__53821;
    wire N__53818;
    wire N__53815;
    wire N__53812;
    wire N__53811;
    wire N__53808;
    wire N__53805;
    wire N__53804;
    wire N__53803;
    wire N__53802;
    wire N__53799;
    wire N__53796;
    wire N__53793;
    wire N__53790;
    wire N__53787;
    wire N__53782;
    wire N__53777;
    wire N__53766;
    wire N__53763;
    wire N__53762;
    wire N__53761;
    wire N__53758;
    wire N__53753;
    wire N__53748;
    wire N__53747;
    wire N__53742;
    wire N__53739;
    wire N__53736;
    wire N__53733;
    wire N__53730;
    wire N__53727;
    wire N__53724;
    wire N__53721;
    wire N__53718;
    wire N__53715;
    wire N__53712;
    wire N__53709;
    wire N__53706;
    wire N__53703;
    wire N__53700;
    wire N__53697;
    wire N__53696;
    wire N__53693;
    wire N__53690;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53670;
    wire N__53667;
    wire N__53664;
    wire N__53661;
    wire N__53658;
    wire N__53655;
    wire N__53652;
    wire N__53649;
    wire N__53646;
    wire N__53643;
    wire N__53640;
    wire N__53637;
    wire N__53634;
    wire N__53631;
    wire N__53628;
    wire N__53625;
    wire N__53622;
    wire N__53619;
    wire N__53616;
    wire N__53613;
    wire N__53612;
    wire N__53609;
    wire N__53606;
    wire N__53601;
    wire N__53598;
    wire N__53597;
    wire N__53594;
    wire N__53591;
    wire N__53588;
    wire N__53585;
    wire N__53582;
    wire N__53579;
    wire N__53576;
    wire N__53573;
    wire N__53572;
    wire N__53569;
    wire N__53568;
    wire N__53567;
    wire N__53566;
    wire N__53563;
    wire N__53560;
    wire N__53559;
    wire N__53558;
    wire N__53555;
    wire N__53552;
    wire N__53549;
    wire N__53546;
    wire N__53541;
    wire N__53536;
    wire N__53523;
    wire N__53520;
    wire N__53519;
    wire N__53516;
    wire N__53515;
    wire N__53512;
    wire N__53509;
    wire N__53508;
    wire N__53507;
    wire N__53504;
    wire N__53503;
    wire N__53500;
    wire N__53497;
    wire N__53494;
    wire N__53493;
    wire N__53492;
    wire N__53489;
    wire N__53484;
    wire N__53481;
    wire N__53478;
    wire N__53475;
    wire N__53470;
    wire N__53465;
    wire N__53462;
    wire N__53459;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53434;
    wire N__53429;
    wire N__53424;
    wire N__53421;
    wire N__53418;
    wire N__53417;
    wire N__53412;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53402;
    wire N__53397;
    wire N__53394;
    wire N__53391;
    wire N__53388;
    wire N__53387;
    wire N__53384;
    wire N__53383;
    wire N__53378;
    wire N__53375;
    wire N__53372;
    wire N__53367;
    wire N__53364;
    wire N__53361;
    wire N__53360;
    wire N__53359;
    wire N__53356;
    wire N__53355;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53341;
    wire N__53338;
    wire N__53335;
    wire N__53328;
    wire N__53327;
    wire N__53326;
    wire N__53325;
    wire N__53322;
    wire N__53319;
    wire N__53316;
    wire N__53315;
    wire N__53312;
    wire N__53311;
    wire N__53310;
    wire N__53309;
    wire N__53308;
    wire N__53307;
    wire N__53306;
    wire N__53305;
    wire N__53304;
    wire N__53303;
    wire N__53302;
    wire N__53295;
    wire N__53292;
    wire N__53285;
    wire N__53278;
    wire N__53271;
    wire N__53266;
    wire N__53265;
    wire N__53262;
    wire N__53257;
    wire N__53252;
    wire N__53249;
    wire N__53246;
    wire N__53241;
    wire N__53236;
    wire N__53235;
    wire N__53234;
    wire N__53231;
    wire N__53226;
    wire N__53221;
    wire N__53216;
    wire N__53211;
    wire N__53210;
    wire N__53209;
    wire N__53208;
    wire N__53205;
    wire N__53202;
    wire N__53201;
    wire N__53200;
    wire N__53197;
    wire N__53196;
    wire N__53193;
    wire N__53184;
    wire N__53177;
    wire N__53176;
    wire N__53175;
    wire N__53174;
    wire N__53173;
    wire N__53168;
    wire N__53165;
    wire N__53162;
    wire N__53159;
    wire N__53156;
    wire N__53153;
    wire N__53144;
    wire N__53139;
    wire N__53138;
    wire N__53133;
    wire N__53130;
    wire N__53127;
    wire N__53124;
    wire N__53121;
    wire N__53118;
    wire N__53115;
    wire N__53112;
    wire N__53111;
    wire N__53110;
    wire N__53105;
    wire N__53102;
    wire N__53099;
    wire N__53096;
    wire N__53093;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53081;
    wire N__53080;
    wire N__53077;
    wire N__53074;
    wire N__53071;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53052;
    wire N__53049;
    wire N__53046;
    wire N__53043;
    wire N__53040;
    wire N__53037;
    wire N__53036;
    wire N__53033;
    wire N__53030;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53013;
    wire N__53010;
    wire N__53007;
    wire N__53006;
    wire N__53001;
    wire N__53000;
    wire N__52999;
    wire N__52998;
    wire N__52997;
    wire N__52994;
    wire N__52991;
    wire N__52984;
    wire N__52977;
    wire N__52976;
    wire N__52973;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52961;
    wire N__52958;
    wire N__52955;
    wire N__52952;
    wire N__52947;
    wire N__52946;
    wire N__52945;
    wire N__52944;
    wire N__52939;
    wire N__52934;
    wire N__52929;
    wire N__52926;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52902;
    wire N__52901;
    wire N__52900;
    wire N__52899;
    wire N__52898;
    wire N__52893;
    wire N__52886;
    wire N__52881;
    wire N__52880;
    wire N__52877;
    wire N__52874;
    wire N__52873;
    wire N__52868;
    wire N__52865;
    wire N__52862;
    wire N__52857;
    wire N__52856;
    wire N__52855;
    wire N__52854;
    wire N__52853;
    wire N__52852;
    wire N__52851;
    wire N__52850;
    wire N__52841;
    wire N__52840;
    wire N__52839;
    wire N__52830;
    wire N__52827;
    wire N__52826;
    wire N__52825;
    wire N__52824;
    wire N__52819;
    wire N__52814;
    wire N__52809;
    wire N__52806;
    wire N__52805;
    wire N__52804;
    wire N__52803;
    wire N__52800;
    wire N__52795;
    wire N__52786;
    wire N__52783;
    wire N__52780;
    wire N__52777;
    wire N__52770;
    wire N__52767;
    wire N__52764;
    wire N__52761;
    wire N__52758;
    wire N__52757;
    wire N__52756;
    wire N__52753;
    wire N__52748;
    wire N__52743;
    wire N__52740;
    wire N__52737;
    wire N__52734;
    wire N__52731;
    wire N__52728;
    wire N__52727;
    wire N__52724;
    wire N__52721;
    wire N__52718;
    wire N__52715;
    wire N__52712;
    wire N__52707;
    wire N__52706;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52692;
    wire N__52689;
    wire N__52686;
    wire N__52685;
    wire N__52682;
    wire N__52679;
    wire N__52676;
    wire N__52671;
    wire N__52670;
    wire N__52665;
    wire N__52662;
    wire N__52659;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52649;
    wire N__52644;
    wire N__52641;
    wire N__52640;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52626;
    wire N__52623;
    wire N__52622;
    wire N__52619;
    wire N__52616;
    wire N__52611;
    wire N__52608;
    wire N__52605;
    wire N__52602;
    wire N__52599;
    wire N__52596;
    wire N__52595;
    wire N__52592;
    wire N__52589;
    wire N__52584;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52572;
    wire N__52571;
    wire N__52570;
    wire N__52569;
    wire N__52566;
    wire N__52563;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52555;
    wire N__52552;
    wire N__52547;
    wire N__52544;
    wire N__52543;
    wire N__52542;
    wire N__52541;
    wire N__52540;
    wire N__52537;
    wire N__52528;
    wire N__52527;
    wire N__52524;
    wire N__52521;
    wire N__52518;
    wire N__52515;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52492;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52476;
    wire N__52467;
    wire N__52466;
    wire N__52465;
    wire N__52462;
    wire N__52461;
    wire N__52458;
    wire N__52455;
    wire N__52452;
    wire N__52449;
    wire N__52448;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52433;
    wire N__52430;
    wire N__52429;
    wire N__52428;
    wire N__52425;
    wire N__52422;
    wire N__52419;
    wire N__52416;
    wire N__52411;
    wire N__52406;
    wire N__52403;
    wire N__52400;
    wire N__52397;
    wire N__52394;
    wire N__52391;
    wire N__52388;
    wire N__52379;
    wire N__52378;
    wire N__52375;
    wire N__52370;
    wire N__52367;
    wire N__52364;
    wire N__52361;
    wire N__52358;
    wire N__52355;
    wire N__52352;
    wire N__52347;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52319;
    wire N__52316;
    wire N__52315;
    wire N__52314;
    wire N__52311;
    wire N__52304;
    wire N__52299;
    wire N__52298;
    wire N__52297;
    wire N__52294;
    wire N__52291;
    wire N__52288;
    wire N__52283;
    wire N__52278;
    wire N__52277;
    wire N__52274;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52247;
    wire N__52244;
    wire N__52239;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52212;
    wire N__52209;
    wire N__52206;
    wire N__52205;
    wire N__52200;
    wire N__52197;
    wire N__52196;
    wire N__52195;
    wire N__52194;
    wire N__52193;
    wire N__52186;
    wire N__52185;
    wire N__52184;
    wire N__52179;
    wire N__52176;
    wire N__52173;
    wire N__52170;
    wire N__52169;
    wire N__52166;
    wire N__52163;
    wire N__52160;
    wire N__52155;
    wire N__52152;
    wire N__52149;
    wire N__52146;
    wire N__52137;
    wire N__52136;
    wire N__52135;
    wire N__52134;
    wire N__52133;
    wire N__52132;
    wire N__52131;
    wire N__52130;
    wire N__52127;
    wire N__52126;
    wire N__52111;
    wire N__52110;
    wire N__52109;
    wire N__52106;
    wire N__52105;
    wire N__52104;
    wire N__52101;
    wire N__52098;
    wire N__52095;
    wire N__52092;
    wire N__52089;
    wire N__52082;
    wire N__52081;
    wire N__52080;
    wire N__52077;
    wire N__52072;
    wire N__52067;
    wire N__52062;
    wire N__52057;
    wire N__52054;
    wire N__52047;
    wire N__52044;
    wire N__52041;
    wire N__52038;
    wire N__52035;
    wire N__52032;
    wire N__52031;
    wire N__52026;
    wire N__52023;
    wire N__52020;
    wire N__52019;
    wire N__52014;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51998;
    wire N__51993;
    wire N__51990;
    wire N__51987;
    wire N__51986;
    wire N__51983;
    wire N__51980;
    wire N__51977;
    wire N__51972;
    wire N__51969;
    wire N__51968;
    wire N__51965;
    wire N__51962;
    wire N__51957;
    wire N__51954;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51942;
    wire N__51939;
    wire N__51938;
    wire N__51933;
    wire N__51930;
    wire N__51927;
    wire N__51926;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51911;
    wire N__51908;
    wire N__51905;
    wire N__51900;
    wire N__51899;
    wire N__51896;
    wire N__51893;
    wire N__51892;
    wire N__51891;
    wire N__51888;
    wire N__51883;
    wire N__51880;
    wire N__51875;
    wire N__51872;
    wire N__51869;
    wire N__51864;
    wire N__51861;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51843;
    wire N__51842;
    wire N__51837;
    wire N__51834;
    wire N__51833;
    wire N__51832;
    wire N__51829;
    wire N__51828;
    wire N__51825;
    wire N__51818;
    wire N__51813;
    wire N__51810;
    wire N__51807;
    wire N__51806;
    wire N__51805;
    wire N__51802;
    wire N__51797;
    wire N__51792;
    wire N__51789;
    wire N__51788;
    wire N__51787;
    wire N__51786;
    wire N__51781;
    wire N__51776;
    wire N__51771;
    wire N__51770;
    wire N__51767;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51755;
    wire N__51752;
    wire N__51749;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51732;
    wire N__51729;
    wire N__51726;
    wire N__51725;
    wire N__51722;
    wire N__51719;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51707;
    wire N__51706;
    wire N__51705;
    wire N__51704;
    wire N__51703;
    wire N__51702;
    wire N__51701;
    wire N__51700;
    wire N__51699;
    wire N__51698;
    wire N__51697;
    wire N__51696;
    wire N__51693;
    wire N__51678;
    wire N__51667;
    wire N__51660;
    wire N__51657;
    wire N__51654;
    wire N__51651;
    wire N__51648;
    wire N__51647;
    wire N__51644;
    wire N__51641;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51628;
    wire N__51623;
    wire N__51618;
    wire N__51617;
    wire N__51614;
    wire N__51613;
    wire N__51612;
    wire N__51611;
    wire N__51610;
    wire N__51609;
    wire N__51606;
    wire N__51603;
    wire N__51596;
    wire N__51593;
    wire N__51590;
    wire N__51581;
    wire N__51576;
    wire N__51575;
    wire N__51570;
    wire N__51567;
    wire N__51564;
    wire N__51561;
    wire N__51558;
    wire N__51555;
    wire N__51554;
    wire N__51549;
    wire N__51546;
    wire N__51543;
    wire N__51540;
    wire N__51537;
    wire N__51534;
    wire N__51531;
    wire N__51530;
    wire N__51527;
    wire N__51524;
    wire N__51521;
    wire N__51518;
    wire N__51515;
    wire N__51510;
    wire N__51507;
    wire N__51506;
    wire N__51503;
    wire N__51500;
    wire N__51497;
    wire N__51494;
    wire N__51491;
    wire N__51488;
    wire N__51485;
    wire N__51482;
    wire N__51479;
    wire N__51476;
    wire N__51471;
    wire N__51470;
    wire N__51467;
    wire N__51464;
    wire N__51461;
    wire N__51458;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51438;
    wire N__51435;
    wire N__51432;
    wire N__51429;
    wire N__51426;
    wire N__51423;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51411;
    wire N__51408;
    wire N__51407;
    wire N__51406;
    wire N__51405;
    wire N__51404;
    wire N__51403;
    wire N__51402;
    wire N__51399;
    wire N__51386;
    wire N__51381;
    wire N__51380;
    wire N__51379;
    wire N__51376;
    wire N__51373;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51357;
    wire N__51354;
    wire N__51351;
    wire N__51350;
    wire N__51347;
    wire N__51344;
    wire N__51341;
    wire N__51338;
    wire N__51333;
    wire N__51330;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51312;
    wire N__51311;
    wire N__51308;
    wire N__51305;
    wire N__51302;
    wire N__51299;
    wire N__51296;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51284;
    wire N__51281;
    wire N__51276;
    wire N__51273;
    wire N__51272;
    wire N__51269;
    wire N__51266;
    wire N__51263;
    wire N__51260;
    wire N__51257;
    wire N__51254;
    wire N__51251;
    wire N__51248;
    wire N__51245;
    wire N__51240;
    wire N__51237;
    wire N__51236;
    wire N__51233;
    wire N__51230;
    wire N__51227;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51215;
    wire N__51212;
    wire N__51209;
    wire N__51204;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51179;
    wire N__51176;
    wire N__51171;
    wire N__51168;
    wire N__51165;
    wire N__51162;
    wire N__51159;
    wire N__51156;
    wire N__51155;
    wire N__51152;
    wire N__51149;
    wire N__51146;
    wire N__51143;
    wire N__51138;
    wire N__51135;
    wire N__51132;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51099;
    wire N__51096;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51078;
    wire N__51075;
    wire N__51074;
    wire N__51071;
    wire N__51068;
    wire N__51065;
    wire N__51062;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51042;
    wire N__51039;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51017;
    wire N__51014;
    wire N__51013;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__50997;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50985;
    wire N__50982;
    wire N__50979;
    wire N__50978;
    wire N__50975;
    wire N__50972;
    wire N__50967;
    wire N__50964;
    wire N__50961;
    wire N__50960;
    wire N__50957;
    wire N__50954;
    wire N__50949;
    wire N__50946;
    wire N__50943;
    wire N__50940;
    wire N__50937;
    wire N__50934;
    wire N__50931;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50910;
    wire N__50907;
    wire N__50904;
    wire N__50903;
    wire N__50900;
    wire N__50897;
    wire N__50894;
    wire N__50891;
    wire N__50888;
    wire N__50885;
    wire N__50882;
    wire N__50877;
    wire N__50876;
    wire N__50873;
    wire N__50870;
    wire N__50869;
    wire N__50864;
    wire N__50861;
    wire N__50858;
    wire N__50855;
    wire N__50852;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50838;
    wire N__50835;
    wire N__50834;
    wire N__50831;
    wire N__50828;
    wire N__50827;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50805;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50774;
    wire N__50773;
    wire N__50770;
    wire N__50765;
    wire N__50760;
    wire N__50759;
    wire N__50758;
    wire N__50755;
    wire N__50748;
    wire N__50745;
    wire N__50742;
    wire N__50741;
    wire N__50738;
    wire N__50735;
    wire N__50734;
    wire N__50731;
    wire N__50728;
    wire N__50725;
    wire N__50720;
    wire N__50715;
    wire N__50712;
    wire N__50709;
    wire N__50708;
    wire N__50705;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50693;
    wire N__50688;
    wire N__50687;
    wire N__50686;
    wire N__50679;
    wire N__50676;
    wire N__50675;
    wire N__50674;
    wire N__50671;
    wire N__50664;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50652;
    wire N__50649;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50636;
    wire N__50635;
    wire N__50632;
    wire N__50629;
    wire N__50626;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50610;
    wire N__50609;
    wire N__50608;
    wire N__50605;
    wire N__50598;
    wire N__50595;
    wire N__50594;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50561;
    wire N__50560;
    wire N__50553;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50531;
    wire N__50528;
    wire N__50525;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50508;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50472;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50459;
    wire N__50456;
    wire N__50453;
    wire N__50448;
    wire N__50445;
    wire N__50444;
    wire N__50441;
    wire N__50438;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50418;
    wire N__50415;
    wire N__50412;
    wire N__50409;
    wire N__50406;
    wire N__50403;
    wire N__50400;
    wire N__50399;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50381;
    wire N__50376;
    wire N__50373;
    wire N__50370;
    wire N__50369;
    wire N__50366;
    wire N__50363;
    wire N__50360;
    wire N__50357;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50350;
    wire N__50347;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50319;
    wire N__50310;
    wire N__50307;
    wire N__50306;
    wire N__50303;
    wire N__50300;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50270;
    wire N__50265;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50238;
    wire N__50235;
    wire N__50232;
    wire N__50229;
    wire N__50226;
    wire N__50223;
    wire N__50222;
    wire N__50219;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50207;
    wire N__50204;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50196;
    wire N__50195;
    wire N__50194;
    wire N__50193;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50175;
    wire N__50172;
    wire N__50165;
    wire N__50158;
    wire N__50151;
    wire N__50150;
    wire N__50147;
    wire N__50144;
    wire N__50141;
    wire N__50138;
    wire N__50135;
    wire N__50134;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50108;
    wire N__50105;
    wire N__50098;
    wire N__50091;
    wire N__50088;
    wire N__50087;
    wire N__50084;
    wire N__50081;
    wire N__50078;
    wire N__50073;
    wire N__50072;
    wire N__50069;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50061;
    wire N__50058;
    wire N__50057;
    wire N__50054;
    wire N__50051;
    wire N__50046;
    wire N__50043;
    wire N__50042;
    wire N__50039;
    wire N__50036;
    wire N__50033;
    wire N__50030;
    wire N__50027;
    wire N__50024;
    wire N__50019;
    wire N__50016;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49997;
    wire N__49994;
    wire N__49991;
    wire N__49988;
    wire N__49985;
    wire N__49984;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49974;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49961;
    wire N__49960;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49945;
    wire N__49942;
    wire N__49939;
    wire N__49932;
    wire N__49927;
    wire N__49920;
    wire N__49917;
    wire N__49914;
    wire N__49911;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49839;
    wire N__49836;
    wire N__49833;
    wire N__49830;
    wire N__49827;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49731;
    wire N__49728;
    wire N__49727;
    wire N__49724;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49706;
    wire N__49701;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49686;
    wire N__49683;
    wire N__49682;
    wire N__49677;
    wire N__49674;
    wire N__49673;
    wire N__49670;
    wire N__49667;
    wire N__49662;
    wire N__49659;
    wire N__49656;
    wire N__49653;
    wire N__49650;
    wire N__49647;
    wire N__49646;
    wire N__49643;
    wire N__49640;
    wire N__49637;
    wire N__49634;
    wire N__49631;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49620;
    wire N__49617;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49609;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49595;
    wire N__49592;
    wire N__49589;
    wire N__49578;
    wire N__49575;
    wire N__49572;
    wire N__49569;
    wire N__49566;
    wire N__49563;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49472;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49449;
    wire N__49446;
    wire N__49443;
    wire N__49440;
    wire N__49437;
    wire N__49434;
    wire N__49433;
    wire N__49428;
    wire N__49425;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49413;
    wire N__49412;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49391;
    wire N__49386;
    wire N__49383;
    wire N__49380;
    wire N__49379;
    wire N__49376;
    wire N__49373;
    wire N__49370;
    wire N__49365;
    wire N__49362;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49333;
    wire N__49330;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49308;
    wire N__49307;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49284;
    wire N__49281;
    wire N__49280;
    wire N__49277;
    wire N__49274;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49247;
    wire N__49246;
    wire N__49243;
    wire N__49238;
    wire N__49233;
    wire N__49232;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49208;
    wire N__49205;
    wire N__49202;
    wire N__49197;
    wire N__49194;
    wire N__49193;
    wire N__49192;
    wire N__49189;
    wire N__49184;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49169;
    wire N__49168;
    wire N__49167;
    wire N__49166;
    wire N__49163;
    wire N__49162;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49152;
    wire N__49149;
    wire N__49148;
    wire N__49147;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49137;
    wire N__49126;
    wire N__49123;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49104;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49074;
    wire N__49071;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49055;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49045;
    wire N__49040;
    wire N__49037;
    wire N__49032;
    wire N__49029;
    wire N__49026;
    wire N__49025;
    wire N__49022;
    wire N__49019;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48996;
    wire N__48993;
    wire N__48990;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48980;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48966;
    wire N__48963;
    wire N__48960;
    wire N__48959;
    wire N__48956;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48936;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48917;
    wire N__48916;
    wire N__48913;
    wire N__48908;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48896;
    wire N__48895;
    wire N__48892;
    wire N__48887;
    wire N__48882;
    wire N__48879;
    wire N__48878;
    wire N__48875;
    wire N__48872;
    wire N__48871;
    wire N__48868;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48854;
    wire N__48849;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48837;
    wire N__48836;
    wire N__48831;
    wire N__48830;
    wire N__48827;
    wire N__48824;
    wire N__48821;
    wire N__48816;
    wire N__48815;
    wire N__48814;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48793;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48756;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48744;
    wire N__48741;
    wire N__48738;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48728;
    wire N__48727;
    wire N__48724;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48698;
    wire N__48697;
    wire N__48694;
    wire N__48689;
    wire N__48684;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48674;
    wire N__48671;
    wire N__48668;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48656;
    wire N__48655;
    wire N__48652;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48636;
    wire N__48633;
    wire N__48632;
    wire N__48631;
    wire N__48630;
    wire N__48629;
    wire N__48628;
    wire N__48623;
    wire N__48622;
    wire N__48619;
    wire N__48612;
    wire N__48611;
    wire N__48610;
    wire N__48609;
    wire N__48608;
    wire N__48605;
    wire N__48604;
    wire N__48603;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48582;
    wire N__48579;
    wire N__48568;
    wire N__48565;
    wire N__48560;
    wire N__48553;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48533;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48509;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48491;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48470;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48455;
    wire N__48454;
    wire N__48451;
    wire N__48446;
    wire N__48443;
    wire N__48440;
    wire N__48437;
    wire N__48434;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48420;
    wire N__48417;
    wire N__48416;
    wire N__48411;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48395;
    wire N__48390;
    wire N__48387;
    wire N__48384;
    wire N__48381;
    wire N__48380;
    wire N__48377;
    wire N__48374;
    wire N__48369;
    wire N__48366;
    wire N__48365;
    wire N__48362;
    wire N__48359;
    wire N__48356;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48341;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48321;
    wire N__48320;
    wire N__48317;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48287;
    wire N__48284;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48269;
    wire N__48268;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48256;
    wire N__48249;
    wire N__48248;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48237;
    wire N__48236;
    wire N__48227;
    wire N__48222;
    wire N__48211;
    wire N__48208;
    wire N__48205;
    wire N__48200;
    wire N__48197;
    wire N__48192;
    wire N__48187;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48159;
    wire N__48156;
    wire N__48153;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48122;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48108;
    wire N__48107;
    wire N__48104;
    wire N__48101;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48077;
    wire N__48074;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48064;
    wire N__48057;
    wire N__48056;
    wire N__48055;
    wire N__48054;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48029;
    wire N__48024;
    wire N__48021;
    wire N__48020;
    wire N__48019;
    wire N__48016;
    wire N__48015;
    wire N__48012;
    wire N__48009;
    wire N__48006;
    wire N__48005;
    wire N__48002;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47986;
    wire N__47979;
    wire N__47976;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47918;
    wire N__47917;
    wire N__47914;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47892;
    wire N__47889;
    wire N__47886;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47871;
    wire N__47868;
    wire N__47867;
    wire N__47862;
    wire N__47859;
    wire N__47858;
    wire N__47853;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47837;
    wire N__47832;
    wire N__47829;
    wire N__47828;
    wire N__47825;
    wire N__47822;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47804;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47790;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47765;
    wire N__47764;
    wire N__47761;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47732;
    wire N__47731;
    wire N__47730;
    wire N__47727;
    wire N__47726;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47721;
    wire N__47720;
    wire N__47717;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47698;
    wire N__47697;
    wire N__47696;
    wire N__47689;
    wire N__47688;
    wire N__47687;
    wire N__47686;
    wire N__47685;
    wire N__47684;
    wire N__47683;
    wire N__47680;
    wire N__47677;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47580;
    wire N__47577;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47558;
    wire N__47557;
    wire N__47554;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47532;
    wire N__47529;
    wire N__47526;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47508;
    wire N__47507;
    wire N__47502;
    wire N__47499;
    wire N__47498;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47483;
    wire N__47478;
    wire N__47475;
    wire N__47474;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47462;
    wire N__47457;
    wire N__47454;
    wire N__47453;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47427;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47417;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47403;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47379;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47359;
    wire N__47358;
    wire N__47355;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47335;
    wire N__47332;
    wire N__47329;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47304;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47285;
    wire N__47284;
    wire N__47279;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47264;
    wire N__47261;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47198;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47186;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47166;
    wire N__47165;
    wire N__47162;
    wire N__47159;
    wire N__47156;
    wire N__47153;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47111;
    wire N__47108;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47090;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47076;
    wire N__47073;
    wire N__47070;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47027;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46986;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46922;
    wire N__46917;
    wire N__46914;
    wire N__46913;
    wire N__46908;
    wire N__46905;
    wire N__46904;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46827;
    wire N__46824;
    wire N__46823;
    wire N__46818;
    wire N__46815;
    wire N__46814;
    wire N__46809;
    wire N__46806;
    wire N__46803;
    wire N__46800;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46745;
    wire N__46740;
    wire N__46737;
    wire N__46736;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46721;
    wire N__46718;
    wire N__46715;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46694;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46673;
    wire N__46672;
    wire N__46669;
    wire N__46664;
    wire N__46659;
    wire N__46656;
    wire N__46655;
    wire N__46654;
    wire N__46651;
    wire N__46646;
    wire N__46641;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46627;
    wire N__46626;
    wire N__46625;
    wire N__46624;
    wire N__46621;
    wire N__46618;
    wire N__46609;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46595;
    wire N__46592;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46576;
    wire N__46573;
    wire N__46572;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46555;
    wire N__46550;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46518;
    wire N__46515;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46507;
    wire N__46504;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46490;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46473;
    wire N__46466;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46431;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46423;
    wire N__46418;
    wire N__46415;
    wire N__46410;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46359;
    wire N__46358;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46314;
    wire N__46311;
    wire N__46310;
    wire N__46309;
    wire N__46306;
    wire N__46301;
    wire N__46296;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46157;
    wire N__46156;
    wire N__46155;
    wire N__46154;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46150;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46126;
    wire N__46125;
    wire N__46124;
    wire N__46123;
    wire N__46122;
    wire N__46119;
    wire N__46118;
    wire N__46109;
    wire N__46106;
    wire N__46097;
    wire N__46092;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46069;
    wire N__46068;
    wire N__46067;
    wire N__46066;
    wire N__46065;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45997;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45944;
    wire N__45941;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45773;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45763;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45747;
    wire N__45744;
    wire N__45743;
    wire N__45742;
    wire N__45741;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45720;
    wire N__45717;
    wire N__45712;
    wire N__45709;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45686;
    wire N__45683;
    wire N__45678;
    wire N__45675;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45659;
    wire N__45654;
    wire N__45651;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45623;
    wire N__45620;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45602;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45578;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45545;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45524;
    wire N__45521;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45509;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45485;
    wire N__45484;
    wire N__45481;
    wire N__45480;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45462;
    wire N__45459;
    wire N__45458;
    wire N__45455;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45443;
    wire N__45438;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45426;
    wire N__45423;
    wire N__45422;
    wire N__45421;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45362;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45296;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45258;
    wire N__45257;
    wire N__45256;
    wire N__45253;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45237;
    wire N__45234;
    wire N__45233;
    wire N__45232;
    wire N__45229;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45213;
    wire N__45210;
    wire N__45209;
    wire N__45208;
    wire N__45205;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45189;
    wire N__45186;
    wire N__45185;
    wire N__45180;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45125;
    wire N__45124;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45116;
    wire N__45115;
    wire N__45114;
    wire N__45113;
    wire N__45112;
    wire N__45111;
    wire N__45110;
    wire N__45109;
    wire N__45100;
    wire N__45095;
    wire N__45082;
    wire N__45079;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45063;
    wire N__45062;
    wire N__45061;
    wire N__45058;
    wire N__45057;
    wire N__45056;
    wire N__45051;
    wire N__45048;
    wire N__45043;
    wire N__45040;
    wire N__45033;
    wire N__45030;
    wire N__45029;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45006;
    wire N__45003;
    wire N__45002;
    wire N__45001;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44984;
    wire N__44983;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44966;
    wire N__44965;
    wire N__44958;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44908;
    wire N__44907;
    wire N__44906;
    wire N__44905;
    wire N__44904;
    wire N__44899;
    wire N__44896;
    wire N__44887;
    wire N__44886;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44880;
    wire N__44875;
    wire N__44866;
    wire N__44859;
    wire N__44858;
    wire N__44857;
    wire N__44856;
    wire N__44855;
    wire N__44852;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44841;
    wire N__44838;
    wire N__44833;
    wire N__44830;
    wire N__44821;
    wire N__44820;
    wire N__44819;
    wire N__44816;
    wire N__44811;
    wire N__44806;
    wire N__44799;
    wire N__44798;
    wire N__44797;
    wire N__44796;
    wire N__44795;
    wire N__44794;
    wire N__44793;
    wire N__44788;
    wire N__44785;
    wire N__44776;
    wire N__44775;
    wire N__44774;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44758;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44741;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44717;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44693;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44660;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44645;
    wire N__44642;
    wire N__44639;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44538;
    wire N__44535;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44527;
    wire N__44522;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44498;
    wire N__44495;
    wire N__44494;
    wire N__44493;
    wire N__44490;
    wire N__44485;
    wire N__44482;
    wire N__44477;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44459;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44435;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44408;
    wire N__44405;
    wire N__44404;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44392;
    wire N__44389;
    wire N__44384;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44307;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44192;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44150;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44119;
    wire N__44116;
    wire N__44111;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44093;
    wire N__44092;
    wire N__44089;
    wire N__44088;
    wire N__44085;
    wire N__44084;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44068;
    wire N__44065;
    wire N__44064;
    wire N__44061;
    wire N__44060;
    wire N__44057;
    wire N__44056;
    wire N__44053;
    wire N__44052;
    wire N__44051;
    wire N__44048;
    wire N__44047;
    wire N__44044;
    wire N__44027;
    wire N__44020;
    wire N__44013;
    wire N__44010;
    wire N__44009;
    wire N__44008;
    wire N__44005;
    wire N__44000;
    wire N__43995;
    wire N__43994;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43982;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43961;
    wire N__43960;
    wire N__43957;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43925;
    wire N__43924;
    wire N__43921;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43883;
    wire N__43882;
    wire N__43879;
    wire N__43874;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43848;
    wire N__43845;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43829;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43811;
    wire N__43810;
    wire N__43807;
    wire N__43802;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43781;
    wire N__43780;
    wire N__43777;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43745;
    wire N__43744;
    wire N__43741;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43670;
    wire N__43669;
    wire N__43666;
    wire N__43661;
    wire N__43656;
    wire N__43653;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43619;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43596;
    wire N__43595;
    wire N__43594;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43559;
    wire N__43556;
    wire N__43555;
    wire N__43554;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43523;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43449;
    wire N__43448;
    wire N__43447;
    wire N__43442;
    wire N__43439;
    wire N__43434;
    wire N__43433;
    wire N__43432;
    wire N__43427;
    wire N__43424;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43359;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43344;
    wire N__43343;
    wire N__43340;
    wire N__43337;
    wire N__43332;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43317;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43307;
    wire N__43302;
    wire N__43301;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43235;
    wire N__43234;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43229;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43202;
    wire N__43201;
    wire N__43198;
    wire N__43193;
    wire N__43188;
    wire N__43185;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43179;
    wire N__43178;
    wire N__43177;
    wire N__43176;
    wire N__43175;
    wire N__43174;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43156;
    wire N__43143;
    wire N__43142;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43134;
    wire N__43133;
    wire N__43128;
    wire N__43123;
    wire N__43118;
    wire N__43113;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43080;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43065;
    wire N__43064;
    wire N__43063;
    wire N__43062;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43054;
    wire N__43051;
    wire N__43050;
    wire N__43049;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43014;
    wire N__43013;
    wire N__43010;
    wire N__43009;
    wire N__43002;
    wire N__42999;
    wire N__42998;
    wire N__42997;
    wire N__42996;
    wire N__42995;
    wire N__42990;
    wire N__42989;
    wire N__42988;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42968;
    wire N__42957;
    wire N__42956;
    wire N__42955;
    wire N__42952;
    wire N__42951;
    wire N__42950;
    wire N__42949;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42933;
    wire N__42932;
    wire N__42931;
    wire N__42930;
    wire N__42927;
    wire N__42920;
    wire N__42913;
    wire N__42910;
    wire N__42903;
    wire N__42902;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42833;
    wire N__42832;
    wire N__42831;
    wire N__42830;
    wire N__42827;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42770;
    wire N__42769;
    wire N__42766;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42746;
    wire N__42743;
    wire N__42742;
    wire N__42739;
    wire N__42732;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42720;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42708;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42696;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42681;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42623;
    wire N__42622;
    wire N__42619;
    wire N__42614;
    wire N__42609;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42581;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42558;
    wire N__42557;
    wire N__42556;
    wire N__42553;
    wire N__42550;
    wire N__42547;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42513;
    wire N__42512;
    wire N__42511;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42499;
    wire N__42492;
    wire N__42491;
    wire N__42490;
    wire N__42489;
    wire N__42486;
    wire N__42481;
    wire N__42478;
    wire N__42471;
    wire N__42470;
    wire N__42469;
    wire N__42468;
    wire N__42465;
    wire N__42460;
    wire N__42457;
    wire N__42450;
    wire N__42449;
    wire N__42448;
    wire N__42447;
    wire N__42442;
    wire N__42437;
    wire N__42432;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42423;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42396;
    wire N__42393;
    wire N__42392;
    wire N__42391;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42369;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42353;
    wire N__42352;
    wire N__42349;
    wire N__42348;
    wire N__42343;
    wire N__42342;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42324;
    wire N__42323;
    wire N__42320;
    wire N__42319;
    wire N__42318;
    wire N__42313;
    wire N__42308;
    wire N__42307;
    wire N__42302;
    wire N__42299;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42272;
    wire N__42271;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42242;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42210;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42170;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42153;
    wire N__42152;
    wire N__42151;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42135;
    wire N__42134;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42124;
    wire N__42121;
    wire N__42118;
    wire N__42111;
    wire N__42110;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42066;
    wire N__42065;
    wire N__42062;
    wire N__42059;
    wire N__42056;
    wire N__42053;
    wire N__42048;
    wire N__42045;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42033;
    wire N__42032;
    wire N__42027;
    wire N__42024;
    wire N__42023;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42011;
    wire N__42006;
    wire N__42003;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41991;
    wire N__41990;
    wire N__41987;
    wire N__41982;
    wire N__41979;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41959;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41922;
    wire N__41919;
    wire N__41918;
    wire N__41917;
    wire N__41916;
    wire N__41915;
    wire N__41906;
    wire N__41903;
    wire N__41898;
    wire N__41897;
    wire N__41894;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41871;
    wire N__41870;
    wire N__41869;
    wire N__41866;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41850;
    wire N__41849;
    wire N__41848;
    wire N__41845;
    wire N__41844;
    wire N__41841;
    wire N__41840;
    wire N__41839;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41813;
    wire N__41812;
    wire N__41809;
    wire N__41804;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41792;
    wire N__41787;
    wire N__41784;
    wire N__41783;
    wire N__41782;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41765;
    wire N__41764;
    wire N__41761;
    wire N__41756;
    wire N__41751;
    wire N__41748;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41736;
    wire N__41733;
    wire N__41732;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41693;
    wire N__41690;
    wire N__41689;
    wire N__41686;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41670;
    wire N__41667;
    wire N__41666;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41646;
    wire N__41645;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41627;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41613;
    wire N__41610;
    wire N__41605;
    wire N__41602;
    wire N__41595;
    wire N__41594;
    wire N__41593;
    wire N__41590;
    wire N__41585;
    wire N__41580;
    wire N__41577;
    wire N__41574;
    wire N__41573;
    wire N__41572;
    wire N__41569;
    wire N__41564;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41552;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41542;
    wire N__41539;
    wire N__41534;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41504;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41489;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41432;
    wire N__41429;
    wire N__41428;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41416;
    wire N__41409;
    wire N__41408;
    wire N__41407;
    wire N__41402;
    wire N__41399;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41376;
    wire N__41373;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41361;
    wire N__41358;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41346;
    wire N__41343;
    wire N__41342;
    wire N__41339;
    wire N__41338;
    wire N__41335;
    wire N__41330;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41320;
    wire N__41319;
    wire N__41316;
    wire N__41309;
    wire N__41304;
    wire N__41301;
    wire N__41300;
    wire N__41299;
    wire N__41296;
    wire N__41295;
    wire N__41292;
    wire N__41285;
    wire N__41280;
    wire N__41277;
    wire N__41276;
    wire N__41273;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41258;
    wire N__41255;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41231;
    wire N__41228;
    wire N__41227;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41215;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41193;
    wire N__41192;
    wire N__41189;
    wire N__41188;
    wire N__41185;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41163;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41103;
    wire N__41100;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41088;
    wire N__41085;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40986;
    wire N__40983;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40947;
    wire N__40944;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40914;
    wire N__40911;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40860;
    wire N__40857;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40842;
    wire N__40839;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40812;
    wire N__40811;
    wire N__40810;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40798;
    wire N__40795;
    wire N__40788;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40755;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40676;
    wire N__40673;
    wire N__40672;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40641;
    wire N__40638;
    wire N__40637;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40625;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40491;
    wire N__40488;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40476;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40464;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40452;
    wire N__40449;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40409;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40374;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40319;
    wire N__40318;
    wire N__40317;
    wire N__40314;
    wire N__40309;
    wire N__40306;
    wire N__40299;
    wire N__40298;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40290;
    wire N__40287;
    wire N__40280;
    wire N__40275;
    wire N__40274;
    wire N__40271;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40223;
    wire N__40222;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40210;
    wire N__40209;
    wire N__40208;
    wire N__40207;
    wire N__40206;
    wire N__40205;
    wire N__40204;
    wire N__40203;
    wire N__40202;
    wire N__40199;
    wire N__40194;
    wire N__40179;
    wire N__40178;
    wire N__40177;
    wire N__40174;
    wire N__40167;
    wire N__40162;
    wire N__40155;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40140;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40068;
    wire N__40067;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40049;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40037;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40010;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39989;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39968;
    wire N__39963;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39951;
    wire N__39948;
    wire N__39947;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39896;
    wire N__39895;
    wire N__39894;
    wire N__39889;
    wire N__39884;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39773;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39752;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39722;
    wire N__39719;
    wire N__39718;
    wire N__39713;
    wire N__39710;
    wire N__39705;
    wire N__39704;
    wire N__39703;
    wire N__39698;
    wire N__39695;
    wire N__39690;
    wire N__39689;
    wire N__39686;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39665;
    wire N__39662;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39591;
    wire N__39590;
    wire N__39589;
    wire N__39588;
    wire N__39587;
    wire N__39586;
    wire N__39585;
    wire N__39584;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39572;
    wire N__39569;
    wire N__39562;
    wire N__39559;
    wire N__39546;
    wire N__39545;
    wire N__39544;
    wire N__39543;
    wire N__39542;
    wire N__39539;
    wire N__39538;
    wire N__39537;
    wire N__39534;
    wire N__39533;
    wire N__39530;
    wire N__39529;
    wire N__39528;
    wire N__39523;
    wire N__39518;
    wire N__39507;
    wire N__39504;
    wire N__39495;
    wire N__39494;
    wire N__39493;
    wire N__39492;
    wire N__39491;
    wire N__39490;
    wire N__39489;
    wire N__39488;
    wire N__39487;
    wire N__39486;
    wire N__39485;
    wire N__39480;
    wire N__39475;
    wire N__39462;
    wire N__39459;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39423;
    wire N__39422;
    wire N__39421;
    wire N__39420;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39409;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39402;
    wire N__39401;
    wire N__39396;
    wire N__39387;
    wire N__39382;
    wire N__39379;
    wire N__39378;
    wire N__39377;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39362;
    wire N__39359;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39341;
    wire N__39336;
    wire N__39333;
    wire N__39328;
    wire N__39325;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39313;
    wire N__39312;
    wire N__39311;
    wire N__39306;
    wire N__39293;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39281;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39258;
    wire N__39255;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39237;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39219;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39207;
    wire N__39204;
    wire N__39203;
    wire N__39202;
    wire N__39201;
    wire N__39200;
    wire N__39199;
    wire N__39198;
    wire N__39197;
    wire N__39188;
    wire N__39181;
    wire N__39178;
    wire N__39171;
    wire N__39170;
    wire N__39169;
    wire N__39168;
    wire N__39167;
    wire N__39166;
    wire N__39157;
    wire N__39152;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39042;
    wire N__39041;
    wire N__39038;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39014;
    wire N__39011;
    wire N__39010;
    wire N__39007;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38982;
    wire N__38979;
    wire N__38978;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38951;
    wire N__38950;
    wire N__38949;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38931;
    wire N__38930;
    wire N__38927;
    wire N__38922;
    wire N__38917;
    wire N__38910;
    wire N__38907;
    wire N__38906;
    wire N__38905;
    wire N__38904;
    wire N__38903;
    wire N__38902;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38885;
    wire N__38880;
    wire N__38875;
    wire N__38868;
    wire N__38865;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38832;
    wire N__38831;
    wire N__38830;
    wire N__38829;
    wire N__38826;
    wire N__38821;
    wire N__38816;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38774;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38750;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38715;
    wire N__38714;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38660;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38601;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38593;
    wire N__38590;
    wire N__38585;
    wire N__38582;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38549;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38537;
    wire N__38536;
    wire N__38535;
    wire N__38534;
    wire N__38531;
    wire N__38522;
    wire N__38517;
    wire N__38514;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38490;
    wire N__38489;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38481;
    wire N__38478;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38462;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38381;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38341;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38309;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38261;
    wire N__38258;
    wire N__38257;
    wire N__38250;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38238;
    wire N__38237;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38211;
    wire N__38210;
    wire N__38209;
    wire N__38206;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38192;
    wire N__38189;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38172;
    wire N__38169;
    wire N__38168;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38145;
    wire N__38144;
    wire N__38143;
    wire N__38140;
    wire N__38135;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38115;
    wire N__38114;
    wire N__38113;
    wire N__38112;
    wire N__38111;
    wire N__38104;
    wire N__38103;
    wire N__38102;
    wire N__38101;
    wire N__38096;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38033;
    wire N__38032;
    wire N__38031;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38017;
    wire N__38014;
    wire N__38007;
    wire N__38006;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37988;
    wire N__37985;
    wire N__37984;
    wire N__37981;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37960;
    wire N__37955;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37922;
    wire N__37919;
    wire N__37918;
    wire N__37917;
    wire N__37914;
    wire N__37913;
    wire N__37910;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37890;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37880;
    wire N__37877;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37854;
    wire N__37853;
    wire N__37848;
    wire N__37847;
    wire N__37846;
    wire N__37843;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37827;
    wire N__37824;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37783;
    wire N__37780;
    wire N__37775;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37716;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37668;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37640;
    wire N__37637;
    wire N__37632;
    wire N__37631;
    wire N__37626;
    wire N__37623;
    wire N__37622;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37568;
    wire N__37567;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37541;
    wire N__37536;
    wire N__37533;
    wire N__37532;
    wire N__37531;
    wire N__37530;
    wire N__37529;
    wire N__37528;
    wire N__37527;
    wire N__37526;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37521;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37517;
    wire N__37516;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37466;
    wire N__37461;
    wire N__37458;
    wire N__37457;
    wire N__37456;
    wire N__37453;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37431;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37410;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37359;
    wire N__37358;
    wire N__37355;
    wire N__37350;
    wire N__37347;
    wire N__37346;
    wire N__37345;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37323;
    wire N__37320;
    wire N__37319;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37259;
    wire N__37258;
    wire N__37257;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37248;
    wire N__37247;
    wire N__37246;
    wire N__37245;
    wire N__37236;
    wire N__37231;
    wire N__37230;
    wire N__37221;
    wire N__37216;
    wire N__37213;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37201;
    wire N__37200;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37192;
    wire N__37189;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37161;
    wire N__37160;
    wire N__37159;
    wire N__37156;
    wire N__37155;
    wire N__37154;
    wire N__37151;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37126;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37081;
    wire N__37078;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37056;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37037;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37029;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37013;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36989;
    wire N__36988;
    wire N__36987;
    wire N__36986;
    wire N__36985;
    wire N__36984;
    wire N__36983;
    wire N__36982;
    wire N__36979;
    wire N__36966;
    wire N__36961;
    wire N__36958;
    wire N__36953;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36887;
    wire N__36886;
    wire N__36883;
    wire N__36878;
    wire N__36873;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36865;
    wire N__36862;
    wire N__36857;
    wire N__36852;
    wire N__36851;
    wire N__36848;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36836;
    wire N__36831;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36821;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36809;
    wire N__36808;
    wire N__36805;
    wire N__36800;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36788;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36658;
    wire N__36655;
    wire N__36650;
    wire N__36645;
    wire N__36644;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36547;
    wire N__36542;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36489;
    wire N__36488;
    wire N__36487;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36472;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36451;
    wire N__36446;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36425;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36415;
    wire N__36412;
    wire N__36407;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36374;
    wire N__36373;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36347;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36293;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36281;
    wire N__36280;
    wire N__36279;
    wire N__36278;
    wire N__36277;
    wire N__36276;
    wire N__36275;
    wire N__36274;
    wire N__36273;
    wire N__36272;
    wire N__36271;
    wire N__36270;
    wire N__36269;
    wire N__36268;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36227;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36212;
    wire N__36211;
    wire N__36210;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36192;
    wire N__36191;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36177;
    wire N__36174;
    wire N__36173;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36141;
    wire N__36138;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36057;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36038;
    wire N__36035;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36005;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35967;
    wire N__35964;
    wire N__35963;
    wire N__35958;
    wire N__35955;
    wire N__35954;
    wire N__35953;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35933;
    wire N__35928;
    wire N__35925;
    wire N__35924;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35867;
    wire N__35866;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35844;
    wire N__35841;
    wire N__35840;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35828;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35796;
    wire N__35795;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35753;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35714;
    wire N__35709;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35670;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35624;
    wire N__35621;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35592;
    wire N__35589;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35537;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35516;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35481;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35457;
    wire N__35454;
    wire N__35453;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35404;
    wire N__35399;
    wire N__35394;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35358;
    wire N__35357;
    wire N__35356;
    wire N__35351;
    wire N__35348;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35232;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35019;
    wire N__35016;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34857;
    wire N__34854;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34806;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34760;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34719;
    wire N__34716;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34625;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34508;
    wire N__34507;
    wire N__34504;
    wire N__34499;
    wire N__34494;
    wire N__34493;
    wire N__34490;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34463;
    wire N__34460;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34426;
    wire N__34421;
    wire N__34416;
    wire N__34415;
    wire N__34412;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34376;
    wire N__34371;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34333;
    wire N__34328;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34316;
    wire N__34315;
    wire N__34312;
    wire N__34307;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34295;
    wire N__34294;
    wire N__34291;
    wire N__34286;
    wire N__34281;
    wire N__34280;
    wire N__34279;
    wire N__34276;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34245;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34233;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34200;
    wire N__34199;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34181;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34152;
    wire N__34149;
    wire N__34148;
    wire N__34147;
    wire N__34144;
    wire N__34139;
    wire N__34134;
    wire N__34133;
    wire N__34132;
    wire N__34129;
    wire N__34124;
    wire N__34119;
    wire N__34118;
    wire N__34115;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34055;
    wire N__34054;
    wire N__34051;
    wire N__34046;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34031;
    wire N__34028;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34004;
    wire N__34001;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33959;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33916;
    wire N__33911;
    wire N__33908;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33872;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33851;
    wire N__33850;
    wire N__33847;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33831;
    wire N__33828;
    wire N__33827;
    wire N__33822;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33779;
    wire N__33778;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33756;
    wire N__33755;
    wire N__33750;
    wire N__33747;
    wire N__33746;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33725;
    wire N__33724;
    wire N__33719;
    wire N__33716;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33689;
    wire N__33688;
    wire N__33685;
    wire N__33680;
    wire N__33675;
    wire N__33672;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33653;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33641;
    wire N__33636;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33572;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33548;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33524;
    wire N__33523;
    wire N__33520;
    wire N__33515;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33494;
    wire N__33493;
    wire N__33490;
    wire N__33485;
    wire N__33480;
    wire N__33479;
    wire N__33474;
    wire N__33471;
    wire N__33470;
    wire N__33465;
    wire N__33462;
    wire N__33461;
    wire N__33460;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33440;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33419;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33395;
    wire N__33394;
    wire N__33391;
    wire N__33386;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33365;
    wire N__33364;
    wire N__33361;
    wire N__33356;
    wire N__33351;
    wire N__33350;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33335;
    wire N__33334;
    wire N__33331;
    wire N__33326;
    wire N__33321;
    wire N__33320;
    wire N__33315;
    wire N__33312;
    wire N__33311;
    wire N__33306;
    wire N__33303;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33254;
    wire N__33253;
    wire N__33250;
    wire N__33245;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33217;
    wire N__33212;
    wire N__33207;
    wire N__33206;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33189;
    wire N__33188;
    wire N__33187;
    wire N__33184;
    wire N__33179;
    wire N__33174;
    wire N__33173;
    wire N__33170;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33153;
    wire N__33152;
    wire N__33151;
    wire N__33148;
    wire N__33143;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33117;
    wire N__33114;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33089;
    wire N__33088;
    wire N__33085;
    wire N__33080;
    wire N__33075;
    wire N__33074;
    wire N__33071;
    wire N__33070;
    wire N__33067;
    wire N__33062;
    wire N__33059;
    wire N__33054;
    wire N__33053;
    wire N__33052;
    wire N__33049;
    wire N__33044;
    wire N__33039;
    wire N__33038;
    wire N__33035;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32937;
    wire N__32934;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32857;
    wire N__32852;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32717;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32674;
    wire N__32667;
    wire N__32664;
    wire N__32663;
    wire N__32662;
    wire N__32661;
    wire N__32656;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32648;
    wire N__32645;
    wire N__32638;
    wire N__32635;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32616;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32604;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32584;
    wire N__32579;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32567;
    wire N__32560;
    wire N__32559;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32036;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31868;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31847;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31748;
    wire N__31745;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31730;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31706;
    wire N__31703;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31688;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31661;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31646;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31607;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31578;
    wire N__31575;
    wire N__31574;
    wire N__31571;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31532;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31442;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31413;
    wire N__31410;
    wire N__31409;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31376;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31364;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31328;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31292;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31277;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31238;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31142;
    wire N__31137;
    wire N__31134;
    wire N__31133;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31064;
    wire N__31061;
    wire N__31056;
    wire N__31053;
    wire N__31052;
    wire N__31051;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31031;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire \Pc2drone_pll_inst.clk_system_pll ;
    wire GNDG0;
    wire VCCG0;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.O_3_21 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_3_15 ;
    wire \pid_alt.O_3_19 ;
    wire \pid_alt.O_3_17 ;
    wire \pid_alt.O_3_18 ;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_3_24 ;
    wire \pid_alt.O_3_22 ;
    wire \pid_alt.O_3_23 ;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.O_3_8 ;
    wire \pid_alt.O_3_16 ;
    wire \pid_alt.O_3_20 ;
    wire \pid_alt.O_3_9 ;
    wire \pid_alt.O_3_13 ;
    wire alt_ki_0;
    wire alt_ki_1;
    wire alt_ki_2;
    wire alt_ki_3;
    wire alt_ki_4;
    wire alt_ki_5;
    wire alt_ki_6;
    wire alt_ki_7;
    wire \pid_alt.O_4_24 ;
    wire \pid_alt.O_4_11 ;
    wire \pid_alt.O_4_18 ;
    wire \pid_alt.O_4_13 ;
    wire \pid_alt.O_4_16 ;
    wire \pid_alt.O_4_22 ;
    wire \pid_alt.O_4_17 ;
    wire \pid_alt.O_4_14 ;
    wire \pid_alt.O_4_9 ;
    wire \pid_alt.O_4_23 ;
    wire \pid_alt.O_4_19 ;
    wire \pid_alt.O_4_12 ;
    wire \pid_alt.O_4_20 ;
    wire \pid_alt.O_4_15 ;
    wire \pid_alt.O_4_6 ;
    wire \pid_alt.O_4_5 ;
    wire \pid_alt.O_4_8 ;
    wire \pid_alt.O_4_7 ;
    wire \pid_alt.O_4_10 ;
    wire \pid_alt.O_4_4 ;
    wire \pid_alt.O_4_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6_cascade_ ;
    wire \pid_alt.un1_pid_prereg_236_1_cascade_ ;
    wire \pid_alt.un1_pid_prereg_236_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_front.O_0_23 ;
    wire \pid_front.O_0_24 ;
    wire \pid_front.O_0_12 ;
    wire \pid_front.O_0_7 ;
    wire \pid_front.O_0_8 ;
    wire \pid_front.O_0_5 ;
    wire \pid_front.O_0_10 ;
    wire \pid_front.O_0_11 ;
    wire \pid_front.O_0_16 ;
    wire \pid_front.O_0_17 ;
    wire \pid_front.O_0_18 ;
    wire \pid_front.O_0_19 ;
    wire \pid_front.O_0_20 ;
    wire \pid_front.O_0_21 ;
    wire \pid_front.O_0_22 ;
    wire \pid_front.O_0_9 ;
    wire bfn_1_17_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_1_18_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire drone_altitude_i_5;
    wire drone_altitude_i_6;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire \pid_alt.O_5_9 ;
    wire \pid_alt.O_5_14 ;
    wire \pid_alt.O_5_24 ;
    wire \pid_alt.O_5_17 ;
    wire \pid_alt.O_5_18 ;
    wire \pid_alt.O_5_19 ;
    wire \pid_alt.O_5_20 ;
    wire \pid_alt.O_5_21 ;
    wire \pid_alt.O_5_22 ;
    wire \pid_alt.O_5_23 ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.O_5_16 ;
    wire \pid_alt.O_5_8 ;
    wire \pid_alt.O_5_15 ;
    wire \pid_alt.O_5_10 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire alt_kd_1;
    wire alt_kd_2;
    wire alt_kd_0;
    wire alt_kd_5;
    wire alt_kd_7;
    wire alt_kd_4;
    wire alt_kd_6;
    wire alt_kd_3;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.N_62_mux_cascade_ ;
    wire \pid_alt.N_94_cascade_ ;
    wire \pid_alt.N_94 ;
    wire bfn_2_12_0_;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.un2_pid_prereg_cry_0 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.un2_pid_prereg_cry_1 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.un2_pid_prereg_cry_2 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.un2_pid_prereg_cry_3 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.un2_pid_prereg_cry_4 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.un2_pid_prereg_cry_5 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.un2_pid_prereg_cry_6 ;
    wire \pid_alt.un2_pid_prereg_cry_7 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire bfn_2_13_0_;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.un2_pid_prereg_cry_8 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.un2_pid_prereg_cry_9 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.un2_pid_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.un2_pid_prereg_cry_11 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.un2_pid_prereg_cry_12 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.un2_pid_prereg_cry_13 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.un2_pid_prereg_cry_14 ;
    wire \pid_alt.un2_pid_prereg_cry_15 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire bfn_2_14_0_;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.un2_pid_prereg_cry_16 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.un2_pid_prereg_cry_17 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.un2_pid_prereg_cry_18 ;
    wire \pid_alt.un2_pid_prereg_cry_19 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.un2_pid_prereg_cry_20 ;
    wire \pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.drone_altitude_i_0 ;
    wire drone_altitude_i_8;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire drone_altitude_i_10;
    wire drone_altitude_i_11;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire drone_altitude_i_4;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire alt_kp_6;
    wire alt_kp_2;
    wire alt_kp_7;
    wire alt_kp_1;
    wire alt_kp_3;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.m7_e_4_cascade_ ;
    wire \pid_alt.N_222_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.un2_pid_prereg_cry_19_c_RNIO4IA ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.m21_e_8_cascade_ ;
    wire \pid_alt.m21_e_2 ;
    wire \pid_alt.un2_pid_prereg_cry_5_c_RNIKEAS ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_4_c_RNIHA9S ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.un2_pid_prereg_cry_3_c_RNIN46R ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_12_c_RNI7SBD ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_11_c_RNIRGEG ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_10_c_RNIOCDG ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_9_c_RNIEPOG ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_17_c_RNIT6FA ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_16_c_RNIR3EA ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_15_c_RNIP0DA ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.un2_pid_prereg_cry_6_c_RNINIBS ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_18_c_RNIV9GA ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.un2_pid_prereg_cry_8_c_RNITQDS ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire drone_altitude_0;
    wire bfn_3_17_0_;
    wire \pid_alt.error_i_acumm_prereg6_cry_0 ;
    wire drone_altitude_2;
    wire \pid_alt.error_i_acumm_prereg6_cry_1 ;
    wire drone_altitude_3;
    wire \pid_alt.error_i_acumm_prereg6_cry_2 ;
    wire drone_altitude_4;
    wire alt_command_0;
    wire \pid_alt.alt_command_i_0 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_3 ;
    wire alt_command_1;
    wire drone_altitude_5;
    wire \pid_alt.alt_command_i_1 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_4 ;
    wire drone_altitude_6;
    wire alt_command_2;
    wire \pid_alt.alt_command_i_2 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_5 ;
    wire alt_command_3;
    wire \pid_alt.alt_command_i_3 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_6 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_7 ;
    wire drone_altitude_8;
    wire alt_command_4;
    wire \pid_alt.alt_command_i_4 ;
    wire bfn_3_18_0_;
    wire alt_command_5;
    wire \pid_alt.alt_command_i_5 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_8 ;
    wire drone_altitude_10;
    wire alt_command_6;
    wire \pid_alt.alt_command_i_6 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_9 ;
    wire drone_altitude_11;
    wire alt_command_7;
    wire \pid_alt.alt_command_i_7 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_10 ;
    wire drone_altitude_12;
    wire \pid_alt.error_i_acumm_prereg6_cry_11 ;
    wire drone_altitude_13;
    wire \pid_alt.error_i_acumm_prereg6_cry_12 ;
    wire drone_altitude_14;
    wire \pid_alt.error_i_acumm_prereg6_cry_13 ;
    wire \pid_alt.drone_altitude_i_15 ;
    wire \pid_alt.error_i_acumm_prereg6_cry_14 ;
    wire \pid_alt.error_i_acumm_prereg6 ;
    wire \pid_alt.error_i_acumm_prereg15lt7 ;
    wire \pid_alt.error_i_acumm_prereg15lto7Z0Z_2 ;
    wire bfn_3_19_0_;
    wire \pid_alt.error_i_acumm_prereg_1_sqmuxa ;
    wire \pid_alt.error_i_acumm_prereg_1_sqmuxa_0 ;
    wire \pid_alt.state_1_0_0 ;
    wire \pid_alt.O_5_12 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.O_5_11 ;
    wire \pid_alt.O_3_5 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.m21_e_0_cascade_ ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.m21_e_10 ;
    wire \pid_alt.N_117_cascade_ ;
    wire \pid_alt.un1_reset_1_0_i_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.N_222 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.un1_reset_1_cascade_ ;
    wire bfn_4_11_0_;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL2IS8Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0K6S5Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0KHT2Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9ABT5Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI00LU2Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIRUDT5Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9AMU2Z0Z_5 ;
    wire bfn_4_12_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIV7JT5Z0Z_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKLA75Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI49QU2Z0Z_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI5H064Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGCG82Z0Z_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL4GT1Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJJ1R3Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIEF0O3Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUEHT1Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire bfn_4_13_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNI060F3Z0Z_15 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGO2F3Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKNGN1Z0Z_15 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0B5F3Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0IN1Z0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGT7F3Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI4AJN1Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISEDF3Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICJKN1Z0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI06021_0Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGRON1Z0Z_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI06021_1Z0Z_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI06021Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI06021_2Z0Z_20 ;
    wire bfn_4_14_0_;
    wire \pid_alt.un1_pid_prereg_0_axb_24 ;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.un2_pid_prereg_cry_0_c_RNIEO2R ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3RCL2Z0Z_1 ;
    wire \pid_alt.O_5_4 ;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.O_3_4 ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.un2_pid_prereg_cry_2_c_RNIK05R ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9F5Q6Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIKNU2Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDJGT5Z0Z_7 ;
    wire \pid_alt.un2_pid_prereg_cry_7_c_RNIQMCS ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIRUOU2Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_16_0_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_1_c_RNIHS3R ;
    wire \pid_alt.error_d_reg_prev_esr_RNI32PN4Z0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire drone_altitude_1;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire drone_H_disp_side_1;
    wire drone_altitude_9;
    wire drone_altitude_i_9;
    wire \pid_alt.O_5_5 ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.O_5_7 ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.O_5_6 ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.O_5_13 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.N_579_0_g ;
    wire \pid_alt.N_579_0 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire bfn_5_7_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.timer_Count_0_sqmuxa_cascade_ ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \pid_alt.source_pid_9_0_tz_6_cascade_ ;
    wire \pid_alt.N_44_cascade_ ;
    wire \pid_alt.N_46_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.N_46 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ;
    wire \pid_alt.N_90_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ;
    wire \pid_alt.N_43 ;
    wire \pid_alt.N_48 ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.N_90 ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.source_pid_9_0_0_4_cascade_ ;
    wire \pid_alt.N_44 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ;
    wire \pid_alt.N_216 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.N_216_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.N_76_i_1 ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.N_93 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire \pid_alt.N_76_i_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGJTE3Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ;
    wire \pid_alt.un2_pid_prereg_cry_14_c_RNINTBA ;
    wire \pid_alt.error_d_reg_prev_esr_RNICEFN1Z0Z_14 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIG0FQ1Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK5TH3Z0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.state_0_g_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.un2_pid_prereg_cry_13_c_RNILQAA ;
    wire \pid_alt.error_d_reg_prev_esr_RNI45EN1Z0Z_13 ;
    wire \Commands_frame_decoder.source_CH1data_1_sqmuxa_0 ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.N_369_2_cascade_ ;
    wire \Commands_frame_decoder.N_370_cascade_ ;
    wire \Commands_frame_decoder.N_369_2 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_i_0_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_1_1_0_cascade_ ;
    wire \Commands_frame_decoder.N_405 ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ;
    wire \Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ;
    wire \Commands_frame_decoder.N_409 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_3_2_cascade_ ;
    wire \Commands_frame_decoder.N_371 ;
    wire \Commands_frame_decoder.stateZ0Z_14 ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.data_rdyc_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ;
    wire \uart_pc.N_152_cascade_ ;
    wire \uart_pc.CO0_cascade_ ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \Commands_frame_decoder.source_CH1data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_CH1data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ;
    wire xy_kp_4;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \Commands_frame_decoder.state_RNIRSI31Z0Z_11 ;
    wire \Commands_frame_decoder.stateZ0Z_13 ;
    wire \pid_alt.source_pid_9_0_tz_6 ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \pid_front.O_0_3 ;
    wire \pid_front.O_0_6 ;
    wire \dron_frame_decoder_1.WDT10_0_cascade_ ;
    wire \dron_frame_decoder_1.N_371_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.N_10_0 ;
    wire \pid_front.N_1662_i ;
    wire \pid_front.error_p_regZ0Z_6 ;
    wire \pid_front.N_1662_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ;
    wire \pid_front.un1_pid_prereg_66_0_cascade_ ;
    wire alt_kp_0;
    wire alt_kp_5;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \Commands_frame_decoder.N_364_0 ;
    wire \Commands_frame_decoder.WDT_RNIET8A1Z0Z_4 ;
    wire \Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire bfn_8_7_0_;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \uart_pc.data_rdyc_1 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.reset6_11 ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_Auxce_0_5_cascade_ ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire \dron_frame_decoder_1.WDT10lt13 ;
    wire \dron_frame_decoder_1.WDT10_0_icf0_1_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_icf0_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_icf1_1_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_icf1 ;
    wire \dron_frame_decoder_1.WDT10lto9_3_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lt10 ;
    wire \dron_frame_decoder_1.m34Z0Z_2 ;
    wire \dron_frame_decoder_1.N_123_mux ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.N_123_mux_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_3Z0Z_1 ;
    wire \dron_frame_decoder_1.state_ns_i_i_a2_1_0 ;
    wire \dron_frame_decoder_1.N_186_cascade_ ;
    wire \dron_frame_decoder_1.N_127_mux ;
    wire \dron_frame_decoder_1.state_ns_i_i_0_0 ;
    wire \reset_module_System.reset6_3 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire \pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ;
    wire \pid_front.N_1668_i ;
    wire \pid_front.error_p_regZ0Z_7 ;
    wire \pid_front.error_d_reg_prevZ0Z_6 ;
    wire \pid_front.N_1668_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ;
    wire \pid_front.O_7 ;
    wire \pid_front.O_8 ;
    wire \pid_front.error_d_regZ0Z_6 ;
    wire \pid_front.O_9 ;
    wire \pid_front.O_0_13 ;
    wire \pid_front.O_0_14 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ;
    wire \pid_front.error_p_regZ0Z_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_5 ;
    wire \pid_front.error_d_regZ0Z_5 ;
    wire \pid_front.error_p_regZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \Commands_frame_decoder.N_402 ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ;
    wire \pid_front.un10lt9_1_cascade_ ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ;
    wire \pid_front.error_i_acumm16lt9_0_cascade_ ;
    wire \pid_front.un10lt9_1 ;
    wire \pid_front.un10lt9_cascade_ ;
    wire \pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ;
    wire \pid_front.error_i_acumm16lto27_7_cascade_ ;
    wire \pid_front.error_i_acumm16lto27_8 ;
    wire \pid_front.error_i_acumm16lto27_9 ;
    wire \pid_front.error_i_acumm16lto27_10 ;
    wire \pid_front.un10lto27_8_cascade_ ;
    wire \pid_front.error_i_acumm_preregZ0Z_26 ;
    wire \pid_front.un10lto27_9_cascade_ ;
    wire \pid_front.un10lto27_11 ;
    wire \pid_front.un10lto27_10 ;
    wire \pid_front.error_i_acumm_preregZ0Z_18 ;
    wire \pid_front.error_i_acumm_preregZ0Z_19 ;
    wire \pid_front.error_i_acumm_preregZ0Z_14 ;
    wire \pid_front.error_i_acumm_preregZ0Z_20 ;
    wire \pid_front.error_i_acumm_preregZ0Z_15 ;
    wire drone_H_disp_side_3;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire uart_input_drone_c;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_9_5_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire bfn_9_6_0_;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.un1_state57_iZ0 ;
    wire \reset_module_System.count_1_1 ;
    wire \reset_module_System.reset6_15 ;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire \uart_drone.N_143_cascade_ ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire bfn_9_8_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire bfn_9_9_0_;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_9_10_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_9_13_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire bfn_9_14_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \pid_front.pid_preregZ0Z_14 ;
    wire \pid_front.pid_prereg_esr_RNIQ6EVZ0Z_17_cascade_ ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a2_0_0_cascade_ ;
    wire \pid_front.N_1698_i_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIUO6U_0Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIROQ33Z0Z_12 ;
    wire \pid_front.error_p_regZ0Z_14 ;
    wire \pid_front.error_d_reg_prevZ0Z_14 ;
    wire \pid_front.N_1674_i ;
    wire \pid_front.error_p_regZ0Z_8 ;
    wire \pid_front.N_1674_i_cascade_ ;
    wire \pid_front.un1_pid_prereg_79_cascade_ ;
    wire \pid_front.error_d_regZ0Z_7 ;
    wire \pid_front.error_d_reg_prevZ0Z_7 ;
    wire \pid_front.error_i_acumm_preregZ0Z_7 ;
    wire \pid_front.error_i_acumm_3_sqmuxa_cascade_ ;
    wire \pid_front.error_i_acumm_preregZ0Z_8 ;
    wire \pid_front.error_i_acumm_3_sqmuxa ;
    wire \pid_front.error_i_acumm_preregZ0Z_9 ;
    wire \pid_front.error_i_acumm_preregZ0Z_1 ;
    wire \pid_front.error_i_acumm_preregZ0Z_2 ;
    wire \pid_front.error_i_acumm16lto27_13 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ;
    wire \pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ;
    wire \pid_front.error_i_acumm_2_sqmuxa_cascade_ ;
    wire \pid_front.error_i_acumm_preregZ0Z_11 ;
    wire \pid_front.error_i_acumm_preregZ0Z_4 ;
    wire \pid_front.error_i_acumm_preregZ0Z_5 ;
    wire \pid_front.error_i_acumm_preregZ0Z_6 ;
    wire \pid_front.error_i_acumm_preregZ0Z_13 ;
    wire \pid_front.error_i_acumm_2_sqmuxa_1 ;
    wire \pid_front.error_i_acumm_preregZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_0_24_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_16_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_16 ;
    wire \pid_front.un1_pid_prereg_0_19_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_17 ;
    wire \pid_front.un1_pid_prereg_0_25_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_24 ;
    wire \pid_front.un1_pid_prereg_0_26_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_26 ;
    wire \pid_front.un1_pid_prereg_0_25 ;
    wire \pid_front.error_i_acumm_preregZ0Z_0 ;
    wire \pid_front.error_i_acumm_preregZ0Z_21 ;
    wire \pid_front.error_i_acumm_preregZ0Z_17 ;
    wire \pid_front.error_i_acumm_preregZ0Z_22 ;
    wire \pid_front.error_i_acumm_preregZ0Z_23 ;
    wire \pid_front.error_i_acumm_preregZ0Z_24 ;
    wire \pid_front.error_i_acumm_preregZ0Z_16 ;
    wire \pid_front.error_i_acumm_preregZ0Z_25 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_4 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10 ;
    wire \pid_front.un10lt11_0 ;
    wire \pid_front.un10lto12 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ;
    wire drone_H_disp_front_1;
    wire drone_H_disp_front_3;
    wire \pid_front.state_RNIPKTDZ0Z_0 ;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire \Commands_frame_decoder.WDT8lto9_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf1 ;
    wire \Commands_frame_decoder.WDT8lt12_0_cascade_ ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.N_145 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.reset6_13 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \uart_drone.N_152_cascade_ ;
    wire \uart_drone.un1_state_7_0_cascade_ ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.un1_state_4_0_cascade_ ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.CO0_cascade_ ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.N_144_1 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \uart_drone.un1_state_2_0 ;
    wire \uart_drone.N_152 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire bfn_10_13_0_;
    wire \pid_front.un11lto30_i_a2 ;
    wire \pid_front.un11lto30_i_a2_0 ;
    wire \pid_front.un11lto30_i_a2_2_and ;
    wire \pid_front.un11lto30_i_a2_1 ;
    wire \pid_front.un11lto30_i_a2_3_and ;
    wire \pid_front.un11lto30_i_a2_2 ;
    wire \pid_front.un11lto30_i_a2_3 ;
    wire \pid_front.un11lto30_i_a2_4 ;
    wire \pid_front.un11lto30_i_a2_5 ;
    wire \pid_front.un11lto30_i_a2_6 ;
    wire bfn_10_14_0_;
    wire \pid_front.un11lto30_i_a2_0_and ;
    wire \pid_front.N_1698_i ;
    wire \pid_front.O_0_15 ;
    wire \pid_front.pid_prereg_esr_RNIBQKJ3Z0Z_20 ;
    wire \pid_front.un11lto30_i_a2_4_and ;
    wire \pid_front.un11lto30_i_a2_6_and ;
    wire \pid_front.un11lto30_i_a2_5_and ;
    wire \pid_front.un11lto30_i_a2_4_and_cascade_ ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ;
    wire \pid_front.N_98_cascade_ ;
    wire \pid_front.N_389_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12_cascade_ ;
    wire \pid_front.un1_pid_prereg_79 ;
    wire \pid_front.un1_pid_prereg_135_0 ;
    wire \pid_front.error_p_reg_esr_RNIJ1FT1Z0Z_12_cascade_ ;
    wire \pid_front.un1_pid_prereg_167_0_1 ;
    wire \pid_front.error_p_regZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIBQB61Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12 ;
    wire \pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12 ;
    wire \pid_front.un1_pid_prereg_0_3_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_3 ;
    wire \pid_front.un1_pid_prereg_0_4_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_5_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_2 ;
    wire \pid_front.error_i_acummZ0Z_0 ;
    wire bfn_10_18_0_;
    wire \pid_front.error_i_acummZ0Z_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_front.error_i_acummZ0Z_2 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_front.error_i_acummZ0Z_4 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_front.error_i_acummZ0Z_5 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4_c_RNILQKE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_front.error_i_acummZ0Z_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_front.error_i_acummZ0Z_7 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_front.error_i_acummZ0Z_8 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ;
    wire bfn_10_19_0_;
    wire \pid_front.error_i_acummZ0Z_9 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_front.error_i_acummZ0Z_10 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_front.error_i_acummZ0Z_11 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_front.error_i_acummZ0Z_12 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_15 ;
    wire bfn_10_20_0_;
    wire \pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_23 ;
    wire \pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ;
    wire bfn_10_21_0_;
    wire \pid_front.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_front.error_i_acummZ0Z_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ;
    wire \pid_front.error_i_acumm_preregZ0Z_28 ;
    wire \pid_front.error_i_acumm_preregZ0Z_27 ;
    wire \pid_front.g0_8_1_cascade_ ;
    wire \pid_front.N_88_0_0_cascade_ ;
    wire \pid_front.g1_cascade_ ;
    wire \pid_front.error_i_regZ0Z_21 ;
    wire \pid_front.N_126_0 ;
    wire \pid_front.g3 ;
    wire \pid_front.error_i_regZ0Z_27 ;
    wire \pid_front.error_i_regZ0Z_23 ;
    wire \pid_front.N_11_0_cascade_ ;
    wire \pid_front.N_12_1_cascade_ ;
    wire \pid_front.error_i_regZ0Z_1 ;
    wire \pid_front.N_9_1 ;
    wire \pid_front.N_9_1_cascade_ ;
    wire \pid_front.N_39_0_cascade_ ;
    wire \pid_front.m7_2_03_cascade_ ;
    wire \pid_front.N_126_cascade_ ;
    wire \pid_front.N_12_1 ;
    wire \pid_front.m1_0_03_cascade_ ;
    wire \pid_front.N_93_0_cascade_ ;
    wire \pid_front.m29_2_03_0 ;
    wire \pid_front.error_i_reg_9_rn_0_25_cascade_ ;
    wire \pid_front.error_i_regZ0Z_25 ;
    wire \pid_front.N_93_0 ;
    wire \pid_front.error_i_regZ0Z_9 ;
    wire \pid_front.error_i_regZ0Z_0 ;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_0_16_cascade_ ;
    wire \pid_front.error_i_regZ0Z_16 ;
    wire \pid_front.m4_2_03 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_16 ;
    wire \pid_front.error_i_regZ0Z_2 ;
    wire debug_CH3_20A_c;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_11_8_0_;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire bfn_11_9_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire \scaler_4.debug_CH3_20A_c_0 ;
    wire frame_decoder_CH4data_0;
    wire bfn_11_10_0_;
    wire frame_decoder_CH4data_1;
    wire \scaler_4.un2_source_data_0 ;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire bfn_11_11_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.N_2232_i_l_ofxZ0 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a4_4 ;
    wire \pid_front.source_pid10lt4_0 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a4_3 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ;
    wire \pid_front.N_99_cascade_ ;
    wire \pid_front.N_98 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_o2_sx ;
    wire \pid_front.N_75_cascade_ ;
    wire \pid_front.N_102 ;
    wire \pid_front.N_99 ;
    wire \pid_front.N_11_i ;
    wire \pid_front.N_76 ;
    wire \pid_front.N_75 ;
    wire \pid_front.error_p_regZ0Z_0 ;
    wire bfn_11_15_0_;
    wire \pid_front.pid_preregZ0Z_0 ;
    wire \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_front.pid_preregZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_0_cry_0 ;
    wire \pid_front.pid_preregZ0Z_2 ;
    wire \pid_front.un1_pid_prereg_0_cry_1 ;
    wire \pid_front.pid_preregZ0Z_3 ;
    wire \pid_front.un1_pid_prereg_0_cry_2 ;
    wire \pid_front.error_p_reg_esr_RNI4U472Z0Z_3 ;
    wire \pid_front.pid_preregZ0Z_4 ;
    wire \pid_front.un1_pid_prereg_0_cry_3 ;
    wire \pid_front.error_p_reg_esr_RNIKJHV_0Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ;
    wire \pid_front.pid_preregZ0Z_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_4 ;
    wire \pid_front.error_p_reg_esr_RNIHMAE2Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIKJHVZ0Z_5 ;
    wire \pid_front.pid_preregZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_0_cry_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_6 ;
    wire \pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ;
    wire \pid_front.pid_preregZ0Z_7 ;
    wire bfn_11_16_0_;
    wire \pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ;
    wire \pid_front.pid_preregZ0Z_8 ;
    wire \pid_front.un1_pid_prereg_0_cry_7 ;
    wire \pid_front.pid_preregZ0Z_9 ;
    wire \pid_front.un1_pid_prereg_0_cry_8 ;
    wire \pid_front.pid_preregZ0Z_10 ;
    wire \pid_front.un1_pid_prereg_0_cry_9 ;
    wire \pid_front.pid_preregZ0Z_11 ;
    wire \pid_front.un1_pid_prereg_0_cry_10 ;
    wire \pid_front.pid_preregZ0Z_12 ;
    wire \pid_front.un1_pid_prereg_0_cry_11 ;
    wire \pid_front.pid_preregZ0Z_13 ;
    wire \pid_front.un1_pid_prereg_0_cry_12 ;
    wire \pid_front.un1_pid_prereg_0_axb_14 ;
    wire \pid_front.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_front.un1_pid_prereg_0_cry_13 ;
    wire \pid_front.un1_pid_prereg_0_cry_14 ;
    wire \pid_front.pid_preregZ0Z_15 ;
    wire bfn_11_17_0_;
    wire \pid_front.pid_preregZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_cry_15 ;
    wire \pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ;
    wire \pid_front.pid_preregZ0Z_17 ;
    wire \pid_front.un1_pid_prereg_0_cry_16 ;
    wire \pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ;
    wire \pid_front.pid_preregZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_cry_17 ;
    wire \pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ;
    wire \pid_front.pid_preregZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_cry_18 ;
    wire \pid_front.pid_preregZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_0_cry_19 ;
    wire \pid_front.pid_preregZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_20 ;
    wire \pid_front.pid_preregZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_cry_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_22 ;
    wire \pid_front.pid_preregZ0Z_23 ;
    wire bfn_11_18_0_;
    wire \pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_24 ;
    wire \pid_front.un1_pid_prereg_0_cry_23 ;
    wire \pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ;
    wire \pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_25 ;
    wire \pid_front.un1_pid_prereg_0_cry_24 ;
    wire \pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_26 ;
    wire \pid_front.un1_pid_prereg_0_cry_25 ;
    wire \pid_front.pid_preregZ0Z_27 ;
    wire \pid_front.un1_pid_prereg_0_cry_26 ;
    wire \pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_28 ;
    wire \pid_front.un1_pid_prereg_0_cry_27 ;
    wire \pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ;
    wire \pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_29 ;
    wire \pid_front.un1_pid_prereg_0_cry_28 ;
    wire \pid_front.un1_pid_prereg_0_axb_30 ;
    wire \pid_front.un1_pid_prereg_0_cry_29 ;
    wire \pid_front.pid_preregZ0Z_30 ;
    wire \pid_front.N_404_g ;
    wire \pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ;
    wire \pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ;
    wire \pid_front.un1_pid_prereg_0_15 ;
    wire \pid_front.un1_pid_prereg_0_15_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ;
    wire \pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_8_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ;
    wire \pid_front.un1_pid_prereg_0_13 ;
    wire \pid_front.un1_pid_prereg_0_13_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_0_9 ;
    wire \pid_front.un1_pid_prereg_0_8 ;
    wire \pid_front.un1_pid_prereg_0_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_11 ;
    wire \pid_front.un1_pid_prereg_0_11_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_10 ;
    wire \pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ;
    wire \pid_front.un1_pid_prereg_370_1 ;
    wire \pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_14 ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_12 ;
    wire \pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ;
    wire \pid_front.error_p_regZ0Z_20 ;
    wire \pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ;
    wire \pid_front.m14_0_ns_1_cascade_ ;
    wire \pid_front.N_15_1_cascade_ ;
    wire \pid_front.m104_1_cascade_ ;
    wire \pid_front.m11_2_03_3_i_0 ;
    wire \pid_front.m11_2_03_3_i_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_7 ;
    wire \pid_front.m53_0_ns_1_cascade_ ;
    wire \pid_front.m5_2_03 ;
    wire \pid_front.error_i_reg_9_rn_0_17_cascade_ ;
    wire \pid_front.error_i_regZ0Z_17 ;
    wire \pid_front.N_44_1_cascade_ ;
    wire \pid_front.N_46_1_cascade_ ;
    wire \pid_front.m27_2_03_0 ;
    wire \pid_front.N_44_1 ;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_17 ;
    wire \pid_front.N_50_1_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_0_19 ;
    wire \pid_front.error_i_regZ0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_17 ;
    wire \pid_front.N_51_1 ;
    wire \pid_front.N_51_1_cascade_ ;
    wire \pid_front.N_47_1_cascade_ ;
    wire \pid_front.N_45_1 ;
    wire \pid_front.N_126 ;
    wire \pid_front.N_88_0_cascade_ ;
    wire \pid_front.N_89_0 ;
    wire \pid_front.N_88_0 ;
    wire \pid_front.N_90_0 ;
    wire \pid_front.g0_6_1 ;
    wire \pid_front.g0_7_1_cascade_ ;
    wire \pid_front.N_89_0_1_cascade_ ;
    wire \pid_front.N_12_1_1 ;
    wire \pid_front.N_116_0_cascade_ ;
    wire \pid_front.un4_error_i_reg_23_ns_1 ;
    wire \pid_front.error_i_reg_9_1_13_cascade_ ;
    wire \pid_front.N_127 ;
    wire \pid_front.error_i_regZ0Z_13 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.N_134_0 ;
    wire bfn_12_7_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire scaler_4_data_14;
    wire bfn_12_8_0_;
    wire bfn_12_9_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire throttle_order_4;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire throttle_order_5;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_12_10_0_;
    wire throttle_order_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_OFF4data_1;
    wire frame_decoder_OFF4data_2;
    wire frame_decoder_OFF4data_3;
    wire frame_decoder_OFF4data_4;
    wire frame_decoder_OFF4data_5;
    wire frame_decoder_OFF4data_6;
    wire frame_decoder_OFF4data_7;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire scaler_4_data_4;
    wire scaler_4_data_5;
    wire \pid_front.state_ns_0_cascade_ ;
    wire \pid_front.un1_reset_0_i ;
    wire \pid_front.state_0_1 ;
    wire \pid_alt.N_76_i ;
    wire \pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ;
    wire \pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ;
    wire \pid_front.error_p_regZ0Z_2 ;
    wire \pid_front.error_d_reg_prevZ0Z_2 ;
    wire \pid_front.error_p_regZ0Z_3 ;
    wire \pid_front.error_d_reg_prevZ0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ;
    wire \pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ;
    wire \pid_front.N_1680_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ;
    wire \pid_front.error_p_regZ0Z_9 ;
    wire \pid_front.error_d_reg_prevZ0Z_8 ;
    wire \pid_front.N_1680_i ;
    wire \pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ;
    wire \pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa ;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ;
    wire front_command_7;
    wire drone_H_disp_front_11;
    wire \pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ;
    wire \pid_front.N_1686_i ;
    wire \pid_front.error_p_reg_esr_RNI6J6A4Z0Z_12 ;
    wire \pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ;
    wire \pid_front.error_d_reg_prev_esr_RNI4CD85Z0Z_12_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ;
    wire \pid_front.un1_pid_prereg_167_0 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ;
    wire \pid_front.un1_pid_prereg_97 ;
    wire \pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIUBM0GZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNI3TJH01Z0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNI5HTGGZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13 ;
    wire \pid_front.un1_pid_prereg_0_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI31A7NZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ;
    wire \pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ;
    wire \pid_front.error_p_regZ0Z_19 ;
    wire \pid_front.error_d_reg_prevZ0Z_19 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ;
    wire \pid_front.error_p_regZ0Z_11 ;
    wire \pid_front.error_d_reg_prevZ0Z_11 ;
    wire \pid_front.error_p_regZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIETB61Z0Z_13 ;
    wire \pid_front.error_d_reg_prevZ0Z_13 ;
    wire \pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_1 ;
    wire \pid_front.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_0 ;
    wire \pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ;
    wire \pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ;
    wire \pid_front.un1_pid_prereg_0_18 ;
    wire \pid_front.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_19 ;
    wire \pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ;
    wire \pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ;
    wire \pid_front.error_p_regZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_22_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_21 ;
    wire \pid_front.un1_pid_prereg_0_20 ;
    wire \pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_22 ;
    wire \pid_front.un1_pid_prereg_0_23 ;
    wire \pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ;
    wire \pid_front.error_d_reg_prevZ0Z_22 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_5 ;
    wire \pid_front.un1_pid_prereg_0_4 ;
    wire \pid_front.un1_pid_prereg_0_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ;
    wire \pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_7 ;
    wire \pid_front.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_6 ;
    wire \pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ;
    wire \pid_front.error_p_regZ0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ;
    wire \pid_front.error_d_reg_prevZ0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ;
    wire \pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ;
    wire \pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ;
    wire \pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ;
    wire \pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ;
    wire \pid_front.g2_cascade_ ;
    wire \dron_frame_decoder_1.drone_H_disp_front_8 ;
    wire drone_H_disp_front_2;
    wire dron_frame_decoder_1_source_H_disp_front_fast_0;
    wire \pid_front.error_axb_0 ;
    wire bfn_12_23_0_;
    wire \pid_front.error_axbZ0Z_1 ;
    wire \pid_front.error_1 ;
    wire \pid_front.error_cry_0 ;
    wire \pid_front.error_axbZ0Z_2 ;
    wire \pid_front.error_cry_1 ;
    wire \pid_front.error_axbZ0Z_3 ;
    wire \pid_front.error_cry_2 ;
    wire drone_H_disp_front_i_4;
    wire front_command_0;
    wire \pid_front.error_cry_3 ;
    wire front_command_1;
    wire \pid_front.error_cry_0_0 ;
    wire front_command_2;
    wire \pid_front.error_cry_1_0 ;
    wire front_command_3;
    wire \pid_front.error_cry_2_0 ;
    wire \pid_front.error_cry_3_0 ;
    wire drone_H_disp_front_i_8;
    wire front_command_4;
    wire bfn_12_24_0_;
    wire drone_H_disp_front_i_9;
    wire front_command_5;
    wire \pid_front.error_cry_4 ;
    wire front_command_6;
    wire \pid_front.error_cry_5 ;
    wire \pid_front.error_axbZ0Z_7 ;
    wire \pid_front.error_cry_6 ;
    wire \pid_front.error_axb_8_l_ofx_0 ;
    wire drone_H_disp_front_12;
    wire \pid_front.error_cry_7 ;
    wire drone_H_disp_front_i_12;
    wire \pid_front.error_cry_8 ;
    wire \pid_front.error_cry_9 ;
    wire \pid_front.error_cry_10 ;
    wire \pid_front.error_2 ;
    wire \pid_front.g0_11_1_cascade_ ;
    wire \pid_front.N_12_1_0_cascade_ ;
    wire \pid_front.N_116_0_0_cascade_ ;
    wire \pid_front.N_117_0 ;
    wire \pid_front.un4_error_i_reg_31_ns_1_0 ;
    wire \pid_front.g0_3_1 ;
    wire \pid_front.N_89_0_0 ;
    wire \pid_front.m6_2_03_cascade_ ;
    wire \pid_front.error_5 ;
    wire \pid_front.error_6 ;
    wire \pid_front.N_27_1_cascade_ ;
    wire \pid_front.N_63_cascade_ ;
    wire \pid_front.N_41_0 ;
    wire \pid_front.N_41_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_10 ;
    wire \pid_front.error_3 ;
    wire \pid_front.error_4 ;
    wire \pid_front.N_30_1 ;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.state_0_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ;
    wire \ppm_encoder_1.N_232_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ;
    wire \ppm_encoder_1.N_139_17 ;
    wire \ppm_encoder_1.N_139 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \ppm_encoder_1.N_313_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire scaler_4_data_10;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire scaler_4_data_7;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire \ppm_encoder_1.N_292_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire throttle_order_6;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire throttle_order_7;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire throttle_order_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire scaler_4_data_12;
    wire scaler_4_data_8;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire scaler_4_data_9;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_order_1;
    wire throttle_order_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire bfn_13_11_0_;
    wire \ppm_encoder_1.un1_elevator_cry_0 ;
    wire \ppm_encoder_1.un1_elevator_cry_1 ;
    wire \ppm_encoder_1.un1_elevator_cry_2 ;
    wire \ppm_encoder_1.un1_elevator_cry_3 ;
    wire \ppm_encoder_1.un1_elevator_cry_4 ;
    wire front_order_6;
    wire \ppm_encoder_1.un1_elevator_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_5 ;
    wire front_order_7;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire bfn_13_12_0_;
    wire front_order_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire front_order_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire xy_kp_0;
    wire xy_kp_1;
    wire xy_kp_2;
    wire xy_kp_3;
    wire xy_kp_5;
    wire xy_kp_6;
    wire xy_kp_7;
    wire \Commands_frame_decoder.state_RNIG48SZ0Z_7 ;
    wire \dron_frame_decoder_1.N_186 ;
    wire \dron_frame_decoder_1.WDT10_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \pid_front.error_d_reg_prevZ0Z_12 ;
    wire \pid_front.error_d_reg_prevZ0Z_20 ;
    wire \pid_front.error_d_reg_prevZ0Z_21 ;
    wire \pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIKI4D7Z0Z_12 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIJ35VFZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIROQ33_0Z0Z_12 ;
    wire \pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ;
    wire \pid_front.un1_pid_prereg_153_0_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNINH0UDZ0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ;
    wire \pid_front.error_d_reg_prevZ0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ;
    wire \pid_front.error_d_reg_prevZ0Z_9 ;
    wire \pid_front.error_p_regZ0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ;
    wire \pid_front.N_196_mux_cascade_ ;
    wire \pid_front.error_i_acumm16lto3 ;
    wire \pid_front.error_i_acumm_2_sqmuxa ;
    wire \pid_front.error_i_acummZ0Z_3 ;
    wire \pid_front.error_i_acumm_1_sqmuxa_1_i ;
    wire pid_side_m153_e_5;
    wire pid_side_m153_e_5_cascade_;
    wire \pid_side.N_196_mux_cascade_ ;
    wire pid_side_m153_e_4;
    wire \pid_front.stateZ0Z_0 ;
    wire \pid_front.stateZ0Z_1 ;
    wire \pid_front.state_RNIVIRQZ0Z_0 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ;
    wire \pid_front.error_p_regZ0Z_15 ;
    wire \pid_front.error_d_reg_prevZ0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ;
    wire \pid_front.error_p_regZ0Z_16 ;
    wire \pid_front.error_d_reg_prevZ0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ;
    wire \pid_front.error_p_regZ0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ;
    wire \pid_front.error_d_reg_prevZ0Z_18 ;
    wire \pid_front.N_404_0 ;
    wire \pid_front.state_RNIM14NZ0Z_0 ;
    wire \pid_front.O_0_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_1 ;
    wire \pid_front.error_p_regZ0Z_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ;
    wire \pid_front.un1_pid_prereg_9_0_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ;
    wire \pid_front.O_3 ;
    wire \pid_front.error_d_regZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_0 ;
    wire \pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ;
    wire \pid_front.O_2 ;
    wire \pid_front.error_d_regZ0Z_0 ;
    wire drone_altitude_15;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_0 ;
    wire drone_altitude_7;
    wire drone_altitude_i_7;
    wire drone_H_disp_front_15;
    wire \dron_frame_decoder_1.drone_H_disp_front_7 ;
    wire drone_H_disp_front_i_7;
    wire \dron_frame_decoder_1.drone_H_disp_front_10 ;
    wire drone_H_disp_front_i_10;
    wire \pid_front.error_cry_5_c_RNIUOTVZ0Z1_cascade_ ;
    wire \pid_front.error_cry_5_c_RNIUOTV1Z0Z_0 ;
    wire \pid_front.N_49_0 ;
    wire \pid_front.N_49_0_cascade_ ;
    wire \pid_front.N_46_1 ;
    wire \pid_front.m134_0_ns_1_cascade_ ;
    wire \pid_front.m19_2_03_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_15 ;
    wire \pid_front.N_48_1 ;
    wire drone_H_disp_front_13;
    wire drone_H_disp_front_i_13;
    wire \dron_frame_decoder_1.drone_H_disp_front_5 ;
    wire drone_H_disp_front_i_5;
    wire \dron_frame_decoder_1.drone_H_disp_front_6 ;
    wire drone_H_disp_front_i_6;
    wire drone_H_disp_front_14;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \dron_frame_decoder_1.N_122_mux_i ;
    wire \pid_front.error_i_reg_esr_RNO_1_0_24_cascade_ ;
    wire \pid_front.error_i_regZ0Z_24 ;
    wire \pid_front.error_cry_7_c_RNI1ADUZ0Z1 ;
    wire \pid_front.error_cry_7_c_RNI1ADU1Z0Z_0 ;
    wire \pid_front.N_22_0_cascade_ ;
    wire \pid_front.N_27_1 ;
    wire \pid_front.error_cry_2_0_c_RNI198HZ0Z2_cascade_ ;
    wire \pid_front.error_cry_2_0_c_RNI198H2Z0Z_0 ;
    wire \pid_front.N_28_1 ;
    wire \pid_front.N_28_1_cascade_ ;
    wire \pid_front.error_8 ;
    wire \pid_front.error_7 ;
    wire \pid_front.N_25_0_cascade_ ;
    wire \pid_front.error_9 ;
    wire \pid_front.error_10 ;
    wire \pid_front.N_21_1_cascade_ ;
    wire \pid_front.N_21_1 ;
    wire \pid_front.N_25_0 ;
    wire \pid_front.m38_1_ns_1 ;
    wire \pid_front.N_39_1_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_1_18 ;
    wire \pid_front.error_i_regZ0Z_18 ;
    wire \pid_front.error_i_reg_9_rn_1_26 ;
    wire \pid_front.N_39_1 ;
    wire \pid_front.error_i_regZ0Z_26 ;
    wire bfn_14_2_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_14_3_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_14_4_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.N_293 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.N_314_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ;
    wire \ppm_encoder_1.N_232 ;
    wire \ppm_encoder_1.PPM_STATE_53_d_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_6_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8 ;
    wire \ppm_encoder_1.N_294_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire front_order_8;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire throttle_order_8;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.N_295_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire front_order_12;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire throttle_order_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \pid_side.un1_reset_0_i_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_1 ;
    wire \pid_side.error_i_acumm16lto3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_2 ;
    wire \pid_side.un10lt9_1 ;
    wire \pid_side.un10lt9_1_cascade_ ;
    wire \pid_side.un10lt9_cascade_ ;
    wire \pid_side.un10lt11_0_cascade_ ;
    wire reset_system;
    wire \pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ;
    wire \pid_side.error_i_acumm_2_sqmuxa_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_4 ;
    wire \pid_side.error_i_acumm_preregZ0Z_5 ;
    wire \pid_side.error_i_acumm_preregZ0Z_6 ;
    wire \pid_side.error_i_acumm_2_sqmuxa_1 ;
    wire \pid_side.error_i_acumm_2_sqmuxa ;
    wire \pid_side.error_i_acumm_1_sqmuxa_1_i ;
    wire \pid_side.error_i_acumm16lto27_10 ;
    wire \pid_side.error_i_acumm16lto27_8 ;
    wire \pid_side.error_i_acumm16lto27_9_cascade_ ;
    wire \pid_side.error_i_acumm16lto27_7 ;
    wire \pid_side.error_i_acumm16lto27_13 ;
    wire \pid_side.un10lto27_8_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_26 ;
    wire \pid_side.error_i_acumm_preregZ0Z_0 ;
    wire \pid_side.error_i_acumm_preregZ0Z_13 ;
    wire \pid_side.error_i_acumm_preregZ0Z_23 ;
    wire \pid_side.error_i_acumm_preregZ0Z_22 ;
    wire \pid_side.error_i_acumm_preregZ0Z_24 ;
    wire \pid_side.error_i_acumm_preregZ0Z_9 ;
    wire \pid_side.error_i_acumm_preregZ0Z_7 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ;
    wire \pid_side.un10lto12 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ;
    wire \pid_side.error_i_acumm16lt9_0 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ;
    wire \pid_side.error_i_acumm_preregZ0Z_10 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ;
    wire \pid_side.error_i_acumm_preregZ0Z_11 ;
    wire \pid_side.error_i_acumm_preregZ0Z_8 ;
    wire \ppm_encoder_1.N_2569_i ;
    wire pid_front_N_331_cascade_;
    wire pid_side_N_166_mux_cascade_;
    wire \pid_front.N_39_0 ;
    wire \pid_front.error_i_regZ0Z_3 ;
    wire \pid_side.N_41_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_26 ;
    wire \pid_front.m8_2_03_3_i_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_4 ;
    wire \pid_front.state_ns_0 ;
    wire \pid_front.N_54_0 ;
    wire \pid_front.error_i_regZ0Z_11 ;
    wire \pid_front.N_15_1 ;
    wire \pid_front.m3_2_03 ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_7 ;
    wire \pid_side.N_49_0_cascade_ ;
    wire \pid_side.m134_0_ns_1_cascade_ ;
    wire \pid_side.N_11_0_cascade_ ;
    wire \pid_side.N_14_1 ;
    wire \pid_side.N_11_0 ;
    wire \pid_side.N_104_cascade_ ;
    wire \pid_side.error_i_reg_9_1_15_cascade_ ;
    wire \pid_side.m19_2_03_0 ;
    wire \pid_front.m24_2_03_0_cascade_ ;
    wire \pid_front.m8_2_03_3_i_0 ;
    wire \pid_front.error_i_regZ0Z_20 ;
    wire \pid_front.N_57_0_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_0_0_24 ;
    wire \pid_front.m138_0_1 ;
    wire \pid_front.N_22_0 ;
    wire \pid_front.N_57_0 ;
    wire \pid_front.N_129_cascade_ ;
    wire \pid_front.error_i_regZ0Z_12 ;
    wire \pid_front.N_60_0 ;
    wire \pid_front.error_i_reg_9_1_12 ;
    wire \pid_front.error_11 ;
    wire \pid_front.error_12 ;
    wire \pid_front.N_18_1 ;
    wire \pid_front.N_18_1_cascade_ ;
    wire \pid_front.N_37_1_cascade_ ;
    wire \pid_front.error_13 ;
    wire \pid_front.error_14 ;
    wire \pid_front.N_36_0 ;
    wire \pid_side.m18_2_03_4_cascade_ ;
    wire \pid_side.m2_2_03 ;
    wire \pid_front.N_3 ;
    wire \pid_front.m2_0_03_3_i_0_cascade_ ;
    wire \pid_front.m2_2_03_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_1_14_cascade_ ;
    wire \pid_front.error_i_regZ0Z_14 ;
    wire \pid_front.N_37_1 ;
    wire \pid_front.error_15 ;
    wire \pid_front.N_136 ;
    wire \pid_front.N_63 ;
    wire \pid_front.error_cry_2_0_c_RNI1CZ0Z944 ;
    wire \pid_front.error_cry_2_0_c_RNI1C944Z0Z_0 ;
    wire \pid_front.N_110_cascade_ ;
    wire \pid_front.m10_2_03_3_i_0_cascade_ ;
    wire \pid_front.m26_2_03_0 ;
    wire \pid_front.error_i_regZ0Z_22 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_15_4_0_;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_15_5_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.N_286_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.N_221_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.N_291_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.N_300_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire \ppm_encoder_1.N_287 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13 ;
    wire \ppm_encoder_1.N_299_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire front_order_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire throttle_order_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire front_order_1;
    wire \ppm_encoder_1.un1_elevator_cry_0_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_1 ;
    wire front_order_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_3_THRU_CO ;
    wire front_order_4;
    wire \ppm_encoder_1.un1_elevator_cry_4_THRU_CO ;
    wire front_order_5;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire bfn_15_12_0_;
    wire \pid_side.un11lto30_i_a2 ;
    wire \pid_side.un11lto30_i_a2_0 ;
    wire \pid_side.un11lto30_i_a2_1 ;
    wire \pid_side.un11lto30_i_a2_2 ;
    wire \pid_side.un11lto30_i_a2_3 ;
    wire \pid_side.un11lto30_i_a2_4 ;
    wire \pid_side.un11lto30_i_a2_5 ;
    wire \pid_side.un11lto30_i_a2_6 ;
    wire bfn_15_13_0_;
    wire \pid_side.source_pid_1_sqmuxa_1_0_o2_sx ;
    wire \pid_side.N_102 ;
    wire \pid_side.N_389 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \pid_side.pid_prereg_esr_RNIVRQ8Z0Z_20_cascade_ ;
    wire xy_ki_5;
    wire xy_ki_6;
    wire xy_ki_7;
    wire \pid_side.un11lto30_i_a2_5_and ;
    wire \pid_side.un11lto30_i_a2_6_and ;
    wire \pid_side.un11lto30_i_a2_5_and_cascade_ ;
    wire \pid_side.un11lto30_i_a2_4_and ;
    wire \pid_side.error_i_acummZ0Z_0 ;
    wire bfn_15_15_0_;
    wire \pid_side.error_i_acummZ0Z_1 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_side.error_i_acummZ0Z_2 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_side.error_i_acummZ0Z_3 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_side.error_i_acummZ0Z_4 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_side.error_i_acummZ0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_side.error_i_acummZ0Z_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_side.error_i_regZ0Z_7 ;
    wire \pid_side.error_i_acummZ0Z_7 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_side.error_i_acummZ0Z_8 ;
    wire bfn_15_16_0_;
    wire \pid_side.error_i_acummZ0Z_9 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_side.error_i_acummZ0Z_10 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_side.error_i_acummZ0Z_11 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_side.error_i_acummZ0Z_12 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_side.error_i_regZ0Z_13 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_side.error_i_regZ0Z_14 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_side.error_i_regZ0Z_15 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_15 ;
    wire bfn_15_17_0_;
    wire \pid_side.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_23 ;
    wire bfn_15_18_0_;
    wire \pid_side.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_side.error_i_regZ0Z_26 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_side.error_i_acummZ0Z_13 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_side.error_i_acumm_preregZ0Z_27 ;
    wire \pid_side.error_i_acumm_preregZ0Z_25 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire uart_drone_data_1;
    wire \dron_frame_decoder_1.un1_sink_data_valid_1_0_cascade_ ;
    wire \dron_frame_decoder_1.drone_H_disp_side_4 ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire uart_drone_data_rdy;
    wire \pid_side.m45_0_ns_1_cascade_ ;
    wire \pid_side.N_46_1_cascade_ ;
    wire \pid_side.N_46_1 ;
    wire \pid_side.N_50_1_cascade_ ;
    wire \pid_side.error_i_regZ0Z_11 ;
    wire \pid_side.error_i_regZ0Z_27 ;
    wire \pid_side.N_50_1 ;
    wire \pid_side.error_i_regZ0Z_19 ;
    wire \pid_side.error_i_regZ0Z_18 ;
    wire \pid_side.N_3_cascade_ ;
    wire \pid_side.m2_0_03_3_i_0_cascade_ ;
    wire \pid_side.m6_2_03_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_18 ;
    wire \pid_side.m51_0_ns_1_cascade_ ;
    wire \pid_side.N_39_0_cascade_ ;
    wire \pid_side.m7_2_03 ;
    wire \pid_side.error_i_reg_9_rn_0_19 ;
    wire \pid_side.N_53_0 ;
    wire \pid_side.N_53_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_27 ;
    wire \pid_side.error_cry_0_c_RNI9I2AZ0Z2 ;
    wire \pid_side.m104_ns_sx ;
    wire \pid_side.m104_ns_sx_cascade_ ;
    wire \pid_side.N_49_0 ;
    wire \pid_side.error_i_regZ0Z_0 ;
    wire \pid_side.error_i_regZ0Z_1 ;
    wire \pid_side.error_i_regZ0Z_2 ;
    wire \pid_side.N_15_1 ;
    wire \pid_side.N_39_0 ;
    wire \pid_side.error_i_regZ0Z_3 ;
    wire \pid_side.m5_2_03_cascade_ ;
    wire \pid_side.error_i_regZ0Z_17 ;
    wire \pid_side.m27_2_03_0 ;
    wire \pid_side.m11_2_03_3_i_0 ;
    wire \pid_side.error_i_regZ0Z_23 ;
    wire \pid_side.error_i_regZ0Z_24 ;
    wire \pid_side.m136_ns_1 ;
    wire \pid_side.N_110_cascade_ ;
    wire \pid_side.m2_0_03_3_i_0 ;
    wire \pid_front.N_110 ;
    wire \pid_front.error_i_regZ0Z_6 ;
    wire \pid_front.N_15_0 ;
    wire \pid_front.N_32_0 ;
    wire \pid_front.N_32_0_cascade_ ;
    wire \pid_front.N_29_1 ;
    wire \pid_front.error_i_regZ0Z_8 ;
    wire \pid_front.m1_0_03 ;
    wire \pid_front.N_117_cascade_ ;
    wire \pid_front.N_116_0 ;
    wire \pid_front.error_i_regZ0Z_5 ;
    wire \pid_front.state_ns_0_0 ;
    wire pid_side_error_i_reg_9_sn_27;
    wire \pid_front.m2_0_03_3_i_0 ;
    wire \pid_front.N_55_0 ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.N_290 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGAZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.throttle_m_1_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire front_order_0;
    wire throttle_order_0;
    wire \ppm_encoder_1.elevatorZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0 ;
    wire \ppm_encoder_1.aileronZ0Z_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_0_cascade_ ;
    wire \ppm_encoder_1.N_289 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ;
    wire \ppm_encoder_1.un1_elevator_cry_2_THRU_CO ;
    wire front_order_3;
    wire \ppm_encoder_1.elevatorZ0Z_3 ;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire throttle_order_3;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.aileronZ0Z_3 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.N_296_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire side_order_0;
    wire bfn_16_10_0_;
    wire \ppm_encoder_1.un1_aileron_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_0 ;
    wire \ppm_encoder_1.un1_aileron_cry_1 ;
    wire \ppm_encoder_1.un1_aileron_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_2 ;
    wire side_order_4;
    wire \ppm_encoder_1.un1_aileron_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_3 ;
    wire side_order_5;
    wire \ppm_encoder_1.un1_aileron_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_4 ;
    wire side_order_6;
    wire \ppm_encoder_1.un1_aileron_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_5 ;
    wire side_order_7;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire side_order_8;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire bfn_16_11_0_;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire side_order_10;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire side_order_11;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire CONSTANT_ONE_NET;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a4_4 ;
    wire \pid_side.source_pid10lt4_0 ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a4_3 ;
    wire \pid_side.un11lto30_i_a2_0_and ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ;
    wire \pid_side.N_99 ;
    wire \pid_side.N_11_i ;
    wire side_order_12;
    wire \pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ;
    wire \pid_side.error_d_reg_prevZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ;
    wire \pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_2_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_3_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_0 ;
    wire \pid_side.un1_pid_prereg_0_0_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIG7B43Z0Z_12_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_19_cascade_ ;
    wire \pid_side.un1_pid_prereg_97 ;
    wire \pid_side.un1_pid_prereg_0_18_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_14_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ;
    wire \pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_10_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ;
    wire \pid_side.un1_pid_prereg_0_14 ;
    wire \pid_side.un1_pid_prereg_0_15 ;
    wire \pid_side.un1_pid_prereg_0_16_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_17 ;
    wire \pid_side.un1_pid_prereg_0_16 ;
    wire \pid_side.un1_pid_prereg_0_11_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_12 ;
    wire \pid_side.un1_pid_prereg_0_11 ;
    wire \pid_side.un1_pid_prereg_0_10 ;
    wire \pid_side.un1_pid_prereg_0_12_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_13 ;
    wire \pid_side.un1_pid_prereg_0_26 ;
    wire \pid_side.un1_pid_prereg_0_23_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ;
    wire \pid_side.un1_pid_prereg_0_22 ;
    wire \pid_side.un1_pid_prereg_0_23 ;
    wire \pid_side.un1_pid_prereg_0_24_cascade_ ;
    wire \pid_side.un1_pid_prereg_370_1 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ;
    wire \pid_side.un1_pid_prereg_0_25 ;
    wire \pid_side.un1_pid_prereg_0_25_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_24 ;
    wire \pid_side.m11_0_ns_1 ;
    wire \pid_side.m88_0_ns_1_cascade_ ;
    wire \pid_side.N_89_0_cascade_ ;
    wire \pid_side.N_116_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_2_13 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_9 ;
    wire \pid_side.m29_2_03_0_cascade_ ;
    wire \pid_side.error_i_regZ0Z_25 ;
    wire \pid_side.N_117_cascade_ ;
    wire \pid_side.N_116_0 ;
    wire \pid_side.error_i_regZ0Z_5 ;
    wire \pid_side.N_41_0 ;
    wire \pid_side.N_39_1 ;
    wire \pid_side.error_i_regZ0Z_10 ;
    wire \pid_side.error_i_regZ0Z_4 ;
    wire \pid_side.N_55_0 ;
    wire \pid_side.N_110 ;
    wire \pid_side.error_i_regZ0Z_6 ;
    wire drone_H_disp_front_0;
    wire \pid_front.m0_0_03 ;
    wire \pid_front.m0_0_03_cascade_ ;
    wire \pid_front.un4_error_i_reg_22_nsZ0Z_1 ;
    wire \pid_side.m0_0_03 ;
    wire xy_ki_fast_2;
    wire \pid_side.m0_0_03_cascade_ ;
    wire \pid_side.N_32_0_cascade_ ;
    wire \pid_side.N_15_0 ;
    wire \pid_side.N_27_1_cascade_ ;
    wire \pid_side.N_63 ;
    wire \pid_side.error_i_reg_esr_RNO_3Z0Z_24 ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_24 ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_24 ;
    wire \pid_side.N_27_1 ;
    wire \pid_side.N_28_1 ;
    wire \pid_side.N_25_0 ;
    wire \pid_side.N_25_0_cascade_ ;
    wire \pid_side.N_38_1 ;
    wire \pid_side.m4_2_03 ;
    wire \pid_side.error_i_reg_9_rn_0_16_cascade_ ;
    wire pid_front_error_i_reg_9_sn_19;
    wire \pid_side.error_i_regZ0Z_16 ;
    wire \pid_side.N_58_0 ;
    wire \pid_side.N_36_0 ;
    wire \pid_side.N_36_0_cascade_ ;
    wire \pid_side.N_57_0_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_24 ;
    wire \pid_side.N_29_1 ;
    wire \pid_side.N_32_0 ;
    wire \pid_side.error_i_regZ0Z_8 ;
    wire \pid_side.N_60_0 ;
    wire \pid_side.m0_2_03 ;
    wire \pid_side.N_60_0_cascade_ ;
    wire pid_side_N_166_mux;
    wire \pid_side.error_i_reg_9_rn_1_12_cascade_ ;
    wire \pid_side.error_i_regZ0Z_12 ;
    wire \pid_side.N_57_0 ;
    wire \pid_side.N_129 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \pid_side.state_RNIL5IFZ0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire xy_kd_1;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.N_288 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire front_order_2;
    wire \ppm_encoder_1.un1_elevator_cry_1_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_order_2;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.un1_aileron_cry_1_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_2 ;
    wire pid_altitude_dv;
    wire scaler_4_data_6;
    wire \ppm_encoder_1.aileron_RNI2Q3U4Z0Z_0 ;
    wire bfn_17_8_0_;
    wire \ppm_encoder_1.throttle_RNIFL0A6Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.aileron_RNIA24U4Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.aileron_RNIE64U4Z0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.elevator_RNI0L5L6Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.elevator_RNI5Q5L6Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.throttle_RNI1T1M6Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.throttle_RNI622M6Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.throttle_RNIB72M6Z0Z_8 ;
    wire bfn_17_9_0_;
    wire \ppm_encoder_1.throttle_RNIGC2M6Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.elevator_RNIOVAA6Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.elevator_RNIT4BA6Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.elevator_RNI2ABA6Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.elevator_RNI7FBA6Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.aileron_esr_RNIG1J17Z0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire bfn_17_10_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \pid_side.state_RNIIIOOZ0Z_0 ;
    wire \pid_side.N_61_0 ;
    wire \pid_side.un11lto30_i_a2_2_and ;
    wire \pid_side.un11lto30_i_a2_3_and ;
    wire \pid_side.pid_preregZ0Z_14 ;
    wire \pid_side.pid_prereg_esr_RNIE1A2Z0Z_17_cascade_ ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ;
    wire bfn_17_13_0_;
    wire \pid_side.pid_preregZ0Z_0 ;
    wire \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_side.un1_pid_prereg_0_cry_0 ;
    wire \pid_side.un1_pid_prereg_0_cry_1 ;
    wire \pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ;
    wire \pid_side.un1_pid_prereg_0_cry_2 ;
    wire \pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ;
    wire \pid_side.pid_preregZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_0_cry_3 ;
    wire \pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ;
    wire \pid_side.pid_preregZ0Z_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_4 ;
    wire \pid_side.pid_preregZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_0_cry_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_6 ;
    wire \pid_side.pid_preregZ0Z_7 ;
    wire bfn_17_14_0_;
    wire \pid_side.pid_preregZ0Z_8 ;
    wire \pid_side.un1_pid_prereg_0_cry_7 ;
    wire \pid_side.un1_pid_prereg_0_cry_8 ;
    wire \pid_side.pid_preregZ0Z_10 ;
    wire \pid_side.un1_pid_prereg_0_cry_9 ;
    wire \pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ;
    wire \pid_side.pid_preregZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_0_cry_10 ;
    wire \pid_side.pid_preregZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_11 ;
    wire \pid_side.un1_pid_prereg_0_cry_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_side.un1_pid_prereg_0_cry_13 ;
    wire \pid_side.un1_pid_prereg_0_cry_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNINPDOKZ0Z_12 ;
    wire \pid_side.pid_preregZ0Z_15 ;
    wire bfn_17_15_0_;
    wire \pid_side.error_d_reg_prev_esr_RNITHHEAZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIJ1F8FZ0Z_12 ;
    wire \pid_side.pid_preregZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_cry_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ;
    wire \pid_side.pid_preregZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_cry_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ;
    wire \pid_side.pid_preregZ0Z_18 ;
    wire \pid_side.un1_pid_prereg_0_cry_17 ;
    wire \pid_side.pid_preregZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_0_cry_18 ;
    wire \pid_side.pid_preregZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_cry_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ;
    wire \pid_side.pid_preregZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ;
    wire \pid_side.pid_preregZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_0_cry_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ;
    wire \pid_side.pid_preregZ0Z_23 ;
    wire bfn_17_16_0_;
    wire \pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_cry_23 ;
    wire \pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_cry_24 ;
    wire \pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_26 ;
    wire \pid_side.un1_pid_prereg_0_cry_25 ;
    wire \pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_27 ;
    wire \pid_side.un1_pid_prereg_0_cry_26 ;
    wire \pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_28 ;
    wire \pid_side.un1_pid_prereg_0_cry_27 ;
    wire \pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_29 ;
    wire \pid_side.un1_pid_prereg_0_cry_28 ;
    wire \pid_side.un1_pid_prereg_0_axb_30 ;
    wire \pid_side.un1_pid_prereg_0_cry_29 ;
    wire \pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ;
    wire \pid_side.un1_pid_prereg_0_21_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ;
    wire \pid_side.error_i_reg_esr_RNISESSZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_20 ;
    wire \pid_side.un1_pid_prereg_0_19 ;
    wire \pid_side.un1_pid_prereg_0_18 ;
    wire \pid_side.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ;
    wire \pid_side.error_d_reg_prevZ0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ;
    wire \pid_side.error_d_reg_prevZ0Z_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire uart_drone_data_3;
    wire drone_H_disp_side_11;
    wire side_command_7;
    wire uart_drone_data_4;
    wire uart_drone_data_7;
    wire \dron_frame_decoder_1.drone_H_disp_side_7 ;
    wire \pid_side.N_12_1 ;
    wire \pid_side.N_126_cascade_ ;
    wire \pid_side.m131_0_ns_1_cascade_ ;
    wire \pid_side.m21_2_03_0 ;
    wire \pid_side.N_89_0 ;
    wire \pid_side.m93_0_ns_1 ;
    wire \pid_side.m13_2_03_4_i_0 ;
    wire pid_side_N_166;
    wire \pid_side.m13_2_03_4_i_0_cascade_ ;
    wire \pid_side.error_i_regZ0Z_9 ;
    wire \pid_side.N_88_0 ;
    wire \pid_side.N_88_0_cascade_ ;
    wire \pid_side.N_126 ;
    wire \pid_side.N_127 ;
    wire \pid_side.error_cry_4_c_RNINOG52Z0Z_1 ;
    wire \pid_side.N_36_0_0_cascade_ ;
    wire \pid_side.g0_9_1_cascade_ ;
    wire \pid_side.N_22_0_0_cascade_ ;
    wire \pid_side.N_57_0_0 ;
    wire \pid_side.g1_cascade_ ;
    wire \pid_side.error_i_regZ0Z_20 ;
    wire \pid_side.g3 ;
    wire \pid_side.m88_0_ns_1_0_cascade_ ;
    wire \pid_side.m48_ns_1 ;
    wire \pid_side.m21_1_cascade_ ;
    wire \pid_side.N_22_0 ;
    wire \pid_side.m30_1_ns_1 ;
    wire \pid_side.error_cry_4_c_RNINOGZ0Z52 ;
    wire \pid_side.N_30_1 ;
    wire \pid_side.m1_0_03 ;
    wire \pid_side.m1_0_03_cascade_ ;
    wire xy_ki_2_rep2;
    wire \pid_side.m1_2_03 ;
    wire \pid_side.N_126_0 ;
    wire \pid_side.g3_0 ;
    wire \pid_side.g1_0_cascade_ ;
    wire \pid_side.error_i_regZ0Z_21 ;
    wire \pid_side.N_89_0_0 ;
    wire \pid_side.N_116_0_0_cascade_ ;
    wire \pid_side.un4_error_i_reg_31_ns_1_0 ;
    wire \pid_side.g2_cascade_ ;
    wire \pid_side.N_117_0 ;
    wire \pid_side.g0_i_m4_0_1 ;
    wire \pid_side.N_10 ;
    wire xy_ki_2_rep1;
    wire \pid_side.N_61_0_0 ;
    wire \pid_side.N_60_0_0_cascade_ ;
    wire \pid_side.un4_error_i_reg_30_ns_1_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.N_2569_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_153_d ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \pid_side.pid_preregZ0Z_1 ;
    wire side_order_1;
    wire \pid_side.pid_preregZ0Z_2 ;
    wire side_order_2;
    wire \pid_side.N_75 ;
    wire \pid_side.pid_preregZ0Z_3 ;
    wire side_order_3;
    wire \pid_side.N_76 ;
    wire \pid_side.pid_preregZ0Z_9 ;
    wire side_order_9;
    wire \pid_side.pid_preregZ0Z_30 ;
    wire \pid_side.N_98 ;
    wire \pid_side.pid_preregZ0Z_13 ;
    wire side_order_13;
    wire \pid_side.state_0_1 ;
    wire \pid_side.un1_reset_0_i ;
    wire \pid_side.state_RNINK4UZ0Z_0_cascade_ ;
    wire debug_CH1_0A_c;
    wire \pid_side.stateZ0Z_0 ;
    wire \pid_side.state_ns_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ;
    wire \pid_side.error_i_acumm_preregZ0Z_28 ;
    wire \pid_side.stateZ0Z_1 ;
    wire \pid_side.error_i_acumm_3_sqmuxa ;
    wire \pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire \pid_side.un1_pid_prereg_0_2 ;
    wire \pid_side.un1_pid_prereg_0_3 ;
    wire \pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ;
    wire \pid_side.un1_pid_prereg_0_5_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_5 ;
    wire \pid_side.un1_pid_prereg_0_6_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ;
    wire \pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_4 ;
    wire \pid_side.error_d_reg_prev_esr_RNI83KO4Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI3AMCBZ0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_153_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIO56DBZ0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ;
    wire \pid_side.un1_pid_prereg_9_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ;
    wire \pid_side.un1_pid_prereg_0_7 ;
    wire \pid_side.un1_pid_prereg_0_6 ;
    wire \pid_side.un1_pid_prereg_0_8_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_9 ;
    wire \pid_side.un1_pid_prereg_0_9_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_8 ;
    wire \pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ;
    wire \pid_side.un1_pid_prereg_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ;
    wire \pid_side.error_i_acumm_preregZ0Z_16 ;
    wire \pid_side.error_i_acumm_preregZ0Z_17 ;
    wire \pid_side.un10lto27_10_cascade_ ;
    wire \pid_side.un10lto27_11 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ;
    wire \pid_side.error_i_acumm_preregZ0Z_21 ;
    wire \pid_side.un10lto27_9 ;
    wire \pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ;
    wire \pid_side.error_i_acumm_preregZ0Z_18 ;
    wire \pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ;
    wire \pid_side.error_i_acumm_preregZ0Z_19 ;
    wire \pid_side.error_i_acumm_preregZ0Z_14 ;
    wire \pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ;
    wire \pid_side.error_i_acumm_preregZ0Z_20 ;
    wire \pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ;
    wire \pid_side.error_i_acumm_preregZ0Z_15 ;
    wire uart_drone_data_5;
    wire \dron_frame_decoder_1.drone_H_disp_side_5 ;
    wire drone_H_disp_side_2;
    wire uart_drone_data_6;
    wire \dron_frame_decoder_1.drone_H_disp_side_6 ;
    wire \pid_side.error_axb_0 ;
    wire bfn_18_19_0_;
    wire \pid_side.error_axbZ0Z_1 ;
    wire \pid_side.error_cry_0 ;
    wire \pid_side.error_axbZ0Z_2 ;
    wire \pid_side.error_cry_1 ;
    wire \pid_side.error_axbZ0Z_3 ;
    wire \pid_side.error_cry_2 ;
    wire side_command_0;
    wire drone_H_disp_side_i_4;
    wire \pid_side.error_cry_3 ;
    wire side_command_1;
    wire drone_H_disp_side_i_5;
    wire \pid_side.error_cry_0_0 ;
    wire drone_H_disp_side_i_6;
    wire side_command_2;
    wire \pid_side.error_cry_1_0 ;
    wire drone_H_disp_side_i_7;
    wire side_command_3;
    wire \pid_side.error_cry_2_0 ;
    wire \pid_side.error_cry_3_0 ;
    wire side_command_4;
    wire bfn_18_20_0_;
    wire drone_H_disp_side_i_9;
    wire side_command_5;
    wire \pid_side.error_9 ;
    wire \pid_side.error_cry_4 ;
    wire side_command_6;
    wire \pid_side.error_cry_5 ;
    wire \pid_side.error_axbZ0Z_7 ;
    wire \pid_side.error_cry_6 ;
    wire \pid_side.error_axb_8_l_ofxZ0 ;
    wire drone_H_disp_side_12;
    wire \pid_side.error_cry_7 ;
    wire drone_H_disp_side_i_12;
    wire drone_H_disp_side_13;
    wire \pid_side.error_cry_8 ;
    wire drone_H_disp_side_i_13;
    wire \pid_side.error_cry_9 ;
    wire drone_H_disp_side_15;
    wire drone_H_disp_side_14;
    wire \pid_side.error_cry_10 ;
    wire \pid_side.m87_0_ns_1 ;
    wire \pid_side.error_10 ;
    wire \pid_side.m87_0_ns_1_0_cascade_ ;
    wire \pid_side.N_88_0_0 ;
    wire \pid_side.error_11 ;
    wire xy_ki_0;
    wire \pid_side.error_12 ;
    wire \pid_side.error_13 ;
    wire \pid_side.m36_1_ns_1_cascade_ ;
    wire \pid_side.error_14 ;
    wire \pid_side.N_37_1 ;
    wire xy_ki_2;
    wire xy_ki_3;
    wire \pid_side.N_37_1_cascade_ ;
    wire \pid_side.error_15 ;
    wire pid_front_N_331;
    wire xy_ki_4;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_22 ;
    wire \pid_side.error_i_regZ0Z_22 ;
    wire \pid_side.state_ns_0_0 ;
    wire drone_H_disp_side_0;
    wire \dron_frame_decoder_1.drone_H_disp_side_8 ;
    wire drone_H_disp_side_i_8;
    wire uart_drone_data_0;
    wire dron_frame_decoder_1_source_H_disp_side_fast_0;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire uart_drone_data_2;
    wire \dron_frame_decoder_1.un1_sink_data_valid_1_0 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_10 ;
    wire drone_H_disp_side_i_10;
    wire \pid_side.error_1 ;
    wire \pid_side.N_12_1_0 ;
    wire xy_ki_0_rep2;
    wire xy_ki_fast_0;
    wire uart_pc_data_1;
    wire xy_ki_1;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ;
    wire \pid_side.g0_3_1_cascade_ ;
    wire \pid_side.N_28_1_0 ;
    wire xy_ki_fast_1;
    wire \pid_side.error_2 ;
    wire \pid_side.m11_0_ns_1_0 ;
    wire \pid_side.error_3 ;
    wire xy_ki_1_rep1;
    wire \pid_side.m30_1_ns_1_0 ;
    wire \pid_side.error_4 ;
    wire \pid_side.N_15_0_0 ;
    wire xy_ki_0_rep1;
    wire \pid_side.error_5 ;
    wire \pid_side.error_6 ;
    wire \pid_side.error_8 ;
    wire \pid_side.error_7 ;
    wire \pid_side.g0_i_m4_1_cascade_ ;
    wire xy_ki_1_rep2;
    wire \pid_side.N_9_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_1_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \pid_side.O_2_6 ;
    wire \pid_side.error_p_regZ0Z_3 ;
    wire \pid_side.O_2_5 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ;
    wire \pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ;
    wire \pid_side.un1_pid_prereg_66_0_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ;
    wire \pid_side.N_1869_i ;
    wire \pid_side.N_1869_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ;
    wire \pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ;
    wire \pid_side.error_d_reg_prevZ0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ;
    wire \pid_side.error_p_reg_esr_RNIT9E37Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ;
    wire \pid_side.error_d_reg_prevZ0Z_10 ;
    wire \pid_side.error_d_reg_prevZ0Z_9 ;
    wire \pid_side.N_1893_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ;
    wire \pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ;
    wire \pid_side.error_p_regZ0Z_2 ;
    wire \pid_side.error_d_reg_prevZ0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ;
    wire \pid_side.error_d_reg_prevZ0Z_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ;
    wire \pid_side.N_1881_i ;
    wire \pid_side.N_1881_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ;
    wire \pid_side.N_1887_i ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ;
    wire \pid_front.O_6 ;
    wire \pid_front.error_d_regZ0Z_4 ;
    wire \pid_front.O_4 ;
    wire \pid_front.error_d_regZ0Z_2 ;
    wire \pid_front.O_11 ;
    wire \pid_front.error_d_regZ0Z_9 ;
    wire \pid_front.O_13 ;
    wire \pid_front.error_d_regZ0Z_11 ;
    wire \pid_front.O_5 ;
    wire \pid_front.error_d_regZ0Z_3 ;
    wire reset_system_g;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.PPM_STATE_53_d ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ;
    wire \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ;
    wire bfn_21_8_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ;
    wire \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire bfn_21_9_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ;
    wire \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire bfn_21_10_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \pid_side.O_2_7 ;
    wire \pid_side.O_1_7 ;
    wire \pid_side.O_1_8 ;
    wire \pid_side.error_d_regZ0Z_6 ;
    wire \pid_side.N_1875_i ;
    wire \pid_side.error_d_reg_prevZ0Z_7 ;
    wire \pid_side.N_478_g ;
    wire \pid_side.error_d_regZ0Z_5 ;
    wire \pid_side.error_d_reg_prevZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_6 ;
    wire \ppm_encoder_1.N_221 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \pid_side.O_1_4 ;
    wire \pid_side.error_d_regZ0Z_2 ;
    wire \pid_side.O_1_9 ;
    wire \pid_side.error_d_regZ0Z_7 ;
    wire \pid_side.O_1_11 ;
    wire \pid_side.error_d_regZ0Z_9 ;
    wire \pid_side.O_2_4 ;
    wire \pid_side.error_p_regZ0Z_1 ;
    wire \pid_side.O_1_12 ;
    wire \pid_side.error_d_regZ0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12 ;
    wire \pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_axb_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12 ;
    wire \pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ;
    wire \pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQ7S9AZ0Z_12 ;
    wire \pid_side.O_1_10 ;
    wire \pid_side.error_d_regZ0Z_8 ;
    wire \pid_side.error_d_reg_prevZ0Z_8 ;
    wire \pid_front.O_12 ;
    wire \pid_front.error_d_regZ0Z_10 ;
    wire \pid_front.O_14 ;
    wire \pid_front.error_d_regZ0Z_12 ;
    wire \pid_front.O_15 ;
    wire \pid_front.error_d_regZ0Z_13 ;
    wire uart_pc_data_4;
    wire xy_kd_4;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ;
    wire \pid_side.error_d_reg_prevZ0Z_4 ;
    wire \pid_side.error_p_regZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ;
    wire \pid_side.error_d_reg_prevZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ;
    wire \pid_side.error_d_reg_prevZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ;
    wire \pid_side.un1_pid_prereg_167_0_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_167_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIOZ0Z_13 ;
    wire \pid_side.error_d_reg_prevZ0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNIMERG_0Z0Z_12 ;
    wire \pid_side.error_p_reg_esr_RNIR3TQ1Z0Z_12 ;
    wire uart_pc_data_0;
    wire xy_kd_0;
    wire uart_pc_data_2;
    wire xy_kd_2;
    wire uart_pc_data_5;
    wire xy_kd_5;
    wire uart_pc_data_7;
    wire xy_kd_7;
    wire uart_pc_data_3;
    wire xy_kd_3;
    wire \pid_side.O_1_5 ;
    wire \pid_side.error_d_regZ0Z_3 ;
    wire \pid_side.O_1_6 ;
    wire \pid_side.error_d_regZ0Z_4 ;
    wire \pid_side.error_d_reg_prevZ0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ;
    wire \pid_side.error_d_reg_prevZ0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ;
    wire \pid_side.O_1_13 ;
    wire \pid_side.N_1905_i ;
    wire \pid_side.N_1905_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIR3TQ1_0Z0Z_12 ;
    wire \pid_side.un1_pid_prereg_79 ;
    wire \pid_side.un1_pid_prereg_79_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIVHA21Z0Z_12 ;
    wire \pid_side.error_p_reg_esr_RNIVKIOZ0Z_12 ;
    wire \pid_side.error_d_reg_prevZ0Z_12 ;
    wire \pid_side.N_478_0 ;
    wire \pid_side.N_1352_g ;
    wire uart_pc_data_6;
    wire xy_kd_6;
    wire \Commands_frame_decoder.state_RNITUI31Z0Z_13 ;
    wire \pid_side.O_2_24 ;
    wire \pid_side.error_p_regZ0Z_21 ;
    wire \pid_side.O_2_16 ;
    wire \pid_side.error_p_regZ0Z_13 ;
    wire \pid_side.O_2_17 ;
    wire \pid_side.error_p_regZ0Z_14 ;
    wire \pid_side.O_2_11 ;
    wire \pid_side.error_p_regZ0Z_8 ;
    wire \pid_side.O_2_19 ;
    wire \pid_side.error_p_regZ0Z_16 ;
    wire \pid_side.O_2_18 ;
    wire \pid_side.error_p_regZ0Z_15 ;
    wire \pid_side.O_2_23 ;
    wire \pid_side.O_2_12 ;
    wire \pid_side.error_p_regZ0Z_9 ;
    wire \pid_side.O_2_22 ;
    wire \pid_side.O_2_20 ;
    wire \pid_side.error_p_regZ0Z_17 ;
    wire \pid_side.O_2_21 ;
    wire \pid_side.error_p_regZ0Z_18 ;
    wire \pid_side.O_2_8 ;
    wire \pid_side.error_p_regZ0Z_5 ;
    wire \pid_side.O_2_10 ;
    wire \pid_side.error_p_regZ0Z_7 ;
    wire \pid_side.O_2_13 ;
    wire \pid_side.error_p_regZ0Z_10 ;
    wire \pid_side.O_2_9 ;
    wire \pid_side.error_p_regZ0Z_6 ;
    wire \pid_side.O_2_3 ;
    wire \pid_side.error_p_regZ0Z_0 ;
    wire \pid_side.O_1_19 ;
    wire \pid_side.error_d_regZ0Z_17 ;
    wire \pid_side.O_1_20 ;
    wire \pid_side.error_d_regZ0Z_18 ;
    wire \pid_side.O_1_18 ;
    wire \pid_side.error_d_regZ0Z_16 ;
    wire \pid_side.O_1_17 ;
    wire \pid_side.error_d_regZ0Z_15 ;
    wire \pid_side.O_1_24 ;
    wire \pid_side.error_d_regZ0Z_22 ;
    wire \pid_side.error_p_regZ0Z_19 ;
    wire \pid_side.error_d_reg_prevZ0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ;
    wire \pid_side.O_1_21 ;
    wire \pid_side.error_d_regZ0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ;
    wire \pid_side.error_d_regZ0Z_11 ;
    wire \pid_side.error_d_reg_prevZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_135_0 ;
    wire \pid_side.O_2_14 ;
    wire \pid_side.error_p_regZ0Z_11 ;
    wire \pid_side.error_p_regZ0Z_20 ;
    wire \pid_side.error_d_reg_prevZ0Z_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ;
    wire \pid_side.O_0_2 ;
    wire \pid_side.error_d_regZ0Z_0 ;
    wire \pid_side.O_1_3 ;
    wire \pid_side.error_d_regZ0Z_1 ;
    wire \pid_side.O_2_15 ;
    wire \pid_side.error_p_regZ0Z_12 ;
    wire \pid_side.O_1_14 ;
    wire \pid_side.error_d_regZ0Z_12 ;
    wire \pid_side.O_1_15 ;
    wire \pid_side.error_d_regZ0Z_13 ;
    wire \pid_side.O_1_16 ;
    wire \pid_side.error_d_regZ0Z_14 ;
    wire \pid_side.O_1_23 ;
    wire \pid_side.error_d_regZ0Z_21 ;
    wire \pid_side.O_1_22 ;
    wire \pid_side.error_d_regZ0Z_20 ;
    wire \pid_side.N_513_0 ;
    wire \pid_front.O_10 ;
    wire \pid_front.error_d_regZ0Z_8 ;
    wire \pid_front.O_19 ;
    wire \pid_front.error_d_regZ0Z_17 ;
    wire \pid_front.O_20 ;
    wire \pid_front.error_d_regZ0Z_18 ;
    wire \pid_front.O_21 ;
    wire \pid_front.error_d_regZ0Z_19 ;
    wire \pid_front.O_22 ;
    wire \pid_front.error_d_regZ0Z_20 ;
    wire \pid_front.O_23 ;
    wire \pid_front.error_d_regZ0Z_21 ;
    wire \pid_front.O_24 ;
    wire \pid_front.error_d_regZ0Z_22 ;
    wire \pid_front.O_18 ;
    wire \pid_front.error_d_regZ0Z_16 ;
    wire \pid_front.O_17 ;
    wire \pid_front.error_d_regZ0Z_15 ;
    wire \pid_front.O_16 ;
    wire \pid_front.error_d_regZ0Z_14 ;
    wire _gnd_net_;
    wire clk_system_pll_g;
    wire \pid_front.N_429_0 ;
    wire N_580_g;

    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .TEST_MODE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVR=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVQ=3'b110;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVF=7'b0111111;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \Pc2drone_pll_inst.Pc2drone_pll_inst_pll  (
            .PLLOUTGLOBAL(),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__60571),
            .PLLOUTCORE(\Pc2drone_pll_inst.clk_system_pll ),
            .LOCK(),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__84558));
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60669),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60668),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__31846,N__31492,N__31531,N__31574,N__31606,N__31645,N__31687,N__31729,N__31769,N__31237,N__31276,N__31327,N__31363,N__31409,N__31441,N__34232}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__32808,N__32832,N__38790,N__37827,N__32907,N__32820,N__32796,N__38685}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_5_24 ,\pid_alt.O_5_23 ,\pid_alt.O_5_22 ,\pid_alt.O_5_21 ,\pid_alt.O_5_20 ,\pid_alt.O_5_19 ,\pid_alt.O_5_18 ,\pid_alt.O_5_17 ,\pid_alt.O_5_16 ,\pid_alt.O_5_15 ,\pid_alt.O_5_14 ,\pid_alt.O_5_13 ,\pid_alt.O_5_12 ,\pid_alt.O_5_11 ,\pid_alt.O_5_10 ,\pid_alt.O_5_9 ,\pid_alt.O_5_8 ,\pid_alt.O_5_7 ,\pid_alt.O_5_6 ,\pid_alt.O_5_5 ,\pid_alt.O_5_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60642),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60570),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__31854,N__31500,N__31536,N__31575,N__31614,N__31653,N__31691,N__31734,N__31773,N__31242,N__31284,N__31329,N__31368,N__31408,N__31449,N__34233}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__31974,N__32085,N__31986,N__32094,N__32076,N__32010,N__32022,N__31998}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_3_24 ,\pid_alt.O_3_23 ,\pid_alt.O_3_22 ,\pid_alt.O_3_21 ,\pid_alt.O_3_20 ,\pid_alt.O_3_19 ,\pid_alt.O_3_18 ,\pid_alt.O_3_17 ,\pid_alt.O_3_16 ,\pid_alt.O_3_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.O_3_5 ,\pid_alt.O_3_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60521),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60455),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .ADDSUBBOT(),
            .A({N__70100,N__70832,N__70919,N__70992,N__71240,N__71330,N__69042,N__72431,N__72347,N__72512,N__72588,N__72797,N__73070,N__73165,N__71675,N__69162}),
            .C({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133}),
            .B({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,N__79754,N__80939,N__79961,N__79146,N__79599,N__80129,N__62270,N__80330}),
            .OHOLDTOP(),
            .O({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,\pid_side.O_1_24 ,\pid_side.O_1_23 ,\pid_side.O_1_22 ,\pid_side.O_1_21 ,\pid_side.O_1_20 ,\pid_side.O_1_19 ,\pid_side.O_1_18 ,\pid_side.O_1_17 ,\pid_side.O_1_16 ,\pid_side.O_1_15 ,\pid_side.O_1_14 ,\pid_side.O_1_13 ,\pid_side.O_1_12 ,\pid_side.O_1_11 ,\pid_side.O_1_10 ,\pid_side.O_1_9 ,\pid_side.O_1_8 ,\pid_side.O_1_7 ,\pid_side.O_1_6 ,\pid_side.O_1_5 ,\pid_side.O_1_4 ,\pid_side.O_1_3 ,\pid_side.O_0_2 ,dangling_wire_149,dangling_wire_150}));
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60454),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60453),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166}),
            .ADDSUBBOT(),
            .A({N__70107,N__70839,N__70920,N__70988,N__71241,N__71331,N__69041,N__72435,N__72351,N__72516,N__72584,N__72801,N__73074,N__73170,N__71676,N__69163}),
            .C({dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182}),
            .B({dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,N__51470,N__51507,N__51530,N__38370,N__51203,N__51236,N__51272,N__51312}),
            .OHOLDTOP(),
            .O({dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,\pid_side.O_2_24 ,\pid_side.O_2_23 ,\pid_side.O_2_22 ,\pid_side.O_2_21 ,\pid_side.O_2_20 ,\pid_side.O_2_19 ,\pid_side.O_2_18 ,\pid_side.O_2_17 ,\pid_side.O_2_16 ,\pid_side.O_2_15 ,\pid_side.O_2_14 ,\pid_side.O_2_13 ,\pid_side.O_2_12 ,\pid_side.O_2_11 ,\pid_side.O_2_10 ,\pid_side.O_2_9 ,\pid_side.O_2_8 ,\pid_side.O_2_7 ,\pid_side.O_2_6 ,\pid_side.O_2_5 ,\pid_side.O_2_4 ,\pid_side.O_2_3 ,dangling_wire_198,dangling_wire_199,dangling_wire_200}));
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60572),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60522),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216}),
            .ADDSUBBOT(),
            .A({N__56534,N__56102,N__56163,N__55745,N__55833,N__53835,N__53885,N__53597,N__53519,N__50310,N__50369,N__50151,N__50222,N__49997,N__49646,N__61838}),
            .C({dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232}),
            .B({dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,N__79758,N__80943,N__79962,N__79142,N__79595,N__80133,N__62274,N__80334}),
            .OHOLDTOP(),
            .O({dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,\pid_front.O_24 ,\pid_front.O_23 ,\pid_front.O_22 ,\pid_front.O_21 ,\pid_front.O_20 ,\pid_front.O_19 ,\pid_front.O_18 ,\pid_front.O_17 ,\pid_front.O_16 ,\pid_front.O_15 ,\pid_front.O_14 ,\pid_front.O_13 ,\pid_front.O_12 ,\pid_front.O_11 ,\pid_front.O_10 ,\pid_front.O_9 ,\pid_front.O_8 ,\pid_front.O_7 ,\pid_front.O_6 ,\pid_front.O_5 ,\pid_front.O_4 ,\pid_front.O_3 ,\pid_front.O_2 ,dangling_wire_248,dangling_wire_249}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60621),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60602),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265}),
            .ADDSUBBOT(),
            .A({N__31847,N__31493,N__31532,N__31570,N__31607,N__31646,N__31692,N__31730,N__31765,N__31238,N__31277,N__31328,N__31364,N__31410,N__31442,N__34219}),
            .C({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .B({dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__30831,N__30843,N__30852,N__30864,N__30873,N__30885,N__30735,N__30747}),
            .OHOLDTOP(),
            .O({dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,\pid_alt.O_4_24 ,\pid_alt.O_4_23 ,\pid_alt.O_4_22 ,\pid_alt.O_4_21 ,\pid_alt.O_4_20 ,\pid_alt.O_4_19 ,\pid_alt.O_4_18 ,\pid_alt.O_4_17 ,\pid_alt.O_4_16 ,\pid_alt.O_4_15 ,\pid_alt.O_4_14 ,\pid_alt.O_4_13 ,\pid_alt.O_4_12 ,\pid_alt.O_4_11 ,\pid_alt.O_4_10 ,\pid_alt.O_4_9 ,\pid_alt.O_4_8 ,\pid_alt.O_4_7 ,\pid_alt.O_4_6 ,\pid_alt.O_4_5 ,\pid_alt.O_4_4 ,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300}));
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__60656),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__60655),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316}),
            .ADDSUBBOT(),
            .A({N__56535,N__56103,N__56162,N__55749,N__55829,N__53831,N__53889,N__53598,N__53523,N__50306,N__50370,N__50150,N__50223,N__49998,N__49647,N__61839}),
            .C({dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332}),
            .B({dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,N__51471,N__51506,N__51534,N__38369,N__51204,N__51240,N__51276,N__51311}),
            .OHOLDTOP(),
            .O({dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,\pid_front.O_0_24 ,\pid_front.O_0_23 ,\pid_front.O_0_22 ,\pid_front.O_0_21 ,\pid_front.O_0_20 ,\pid_front.O_0_19 ,\pid_front.O_0_18 ,\pid_front.O_0_17 ,\pid_front.O_0_16 ,\pid_front.O_0_15 ,\pid_front.O_0_14 ,\pid_front.O_0_13 ,\pid_front.O_0_12 ,\pid_front.O_0_11 ,\pid_front.O_0_10 ,\pid_front.O_0_9 ,\pid_front.O_0_8 ,\pid_front.O_0_7 ,\pid_front.O_0_6 ,\pid_front.O_0_5 ,\pid_front.O_0_4 ,\pid_front.O_0_3 ,dangling_wire_348,dangling_wire_349,dangling_wire_350}));
    IO_PAD \Pc2drone_pll_inst.Pc2drone_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__84558),
            .PACKAGEPIN(clk_system));
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__84544),
            .DIN(N__84543),
            .DOUT(N__84542),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__84544),
            .PADOUT(N__84543),
            .PADIN(N__84542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__84535),
            .DIN(N__84534),
            .DOUT(N__84533),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__84535),
            .PADOUT(N__84534),
            .PADIN(N__84533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39420),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__84526),
            .DIN(N__84525),
            .DOUT(N__84524),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__84526),
            .PADOUT(N__84525),
            .PADIN(N__84524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__84517),
            .DIN(N__84516),
            .DOUT(N__84515),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__84517),
            .PADOUT(N__84516),
            .PADIN(N__84515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__84508),
            .DIN(N__84507),
            .DOUT(N__84506),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__84508),
            .PADOUT(N__84507),
            .PADIN(N__84506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46992),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__84499),
            .DIN(N__84498),
            .DOUT(N__84497),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__84499),
            .PADOUT(N__84498),
            .PADIN(N__84497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__84490),
            .DIN(N__84489),
            .DOUT(N__84488),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__84490),
            .PADOUT(N__84489),
            .PADIN(N__84488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__84481),
            .DIN(N__84480),
            .DOUT(N__84479),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__84481),
            .PADOUT(N__84480),
            .PADIN(N__84479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__84472),
            .DIN(N__84471),
            .DOUT(N__84470),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__84472),
            .PADOUT(N__84471),
            .PADIN(N__84470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43188),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__84463),
            .DIN(N__84462),
            .DOUT(N__84461),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__84463),
            .PADOUT(N__84462),
            .PADIN(N__84461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__67389),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__20429 (
            .O(N__84444),
            .I(N__84441));
    LocalMux I__20428 (
            .O(N__84441),
            .I(N__84438));
    Odrv4 I__20427 (
            .O(N__84438),
            .I(\pid_front.O_21 ));
    InMux I__20426 (
            .O(N__84435),
            .I(N__84426));
    InMux I__20425 (
            .O(N__84434),
            .I(N__84426));
    InMux I__20424 (
            .O(N__84433),
            .I(N__84426));
    LocalMux I__20423 (
            .O(N__84426),
            .I(N__84423));
    Span4Mux_h I__20422 (
            .O(N__84423),
            .I(N__84420));
    Span4Mux_h I__20421 (
            .O(N__84420),
            .I(N__84417));
    Span4Mux_h I__20420 (
            .O(N__84417),
            .I(N__84414));
    Odrv4 I__20419 (
            .O(N__84414),
            .I(\pid_front.error_d_regZ0Z_19 ));
    InMux I__20418 (
            .O(N__84411),
            .I(N__84408));
    LocalMux I__20417 (
            .O(N__84408),
            .I(N__84405));
    Span4Mux_h I__20416 (
            .O(N__84405),
            .I(N__84402));
    Odrv4 I__20415 (
            .O(N__84402),
            .I(\pid_front.O_22 ));
    InMux I__20414 (
            .O(N__84399),
            .I(N__84396));
    LocalMux I__20413 (
            .O(N__84396),
            .I(N__84391));
    InMux I__20412 (
            .O(N__84395),
            .I(N__84386));
    InMux I__20411 (
            .O(N__84394),
            .I(N__84386));
    Span4Mux_v I__20410 (
            .O(N__84391),
            .I(N__84383));
    LocalMux I__20409 (
            .O(N__84386),
            .I(N__84380));
    Sp12to4 I__20408 (
            .O(N__84383),
            .I(N__84377));
    Span12Mux_h I__20407 (
            .O(N__84380),
            .I(N__84374));
    Span12Mux_h I__20406 (
            .O(N__84377),
            .I(N__84371));
    Span12Mux_h I__20405 (
            .O(N__84374),
            .I(N__84368));
    Odrv12 I__20404 (
            .O(N__84371),
            .I(\pid_front.error_d_regZ0Z_20 ));
    Odrv12 I__20403 (
            .O(N__84368),
            .I(\pid_front.error_d_regZ0Z_20 ));
    InMux I__20402 (
            .O(N__84363),
            .I(N__84360));
    LocalMux I__20401 (
            .O(N__84360),
            .I(N__84357));
    Span4Mux_h I__20400 (
            .O(N__84357),
            .I(N__84354));
    Odrv4 I__20399 (
            .O(N__84354),
            .I(\pid_front.O_23 ));
    InMux I__20398 (
            .O(N__84351),
            .I(N__84346));
    InMux I__20397 (
            .O(N__84350),
            .I(N__84341));
    InMux I__20396 (
            .O(N__84349),
            .I(N__84341));
    LocalMux I__20395 (
            .O(N__84346),
            .I(N__84338));
    LocalMux I__20394 (
            .O(N__84341),
            .I(N__84335));
    Span4Mux_h I__20393 (
            .O(N__84338),
            .I(N__84332));
    Span4Mux_v I__20392 (
            .O(N__84335),
            .I(N__84329));
    Sp12to4 I__20391 (
            .O(N__84332),
            .I(N__84326));
    Span4Mux_h I__20390 (
            .O(N__84329),
            .I(N__84323));
    Span12Mux_v I__20389 (
            .O(N__84326),
            .I(N__84318));
    Sp12to4 I__20388 (
            .O(N__84323),
            .I(N__84318));
    Odrv12 I__20387 (
            .O(N__84318),
            .I(\pid_front.error_d_regZ0Z_21 ));
    InMux I__20386 (
            .O(N__84315),
            .I(N__84312));
    LocalMux I__20385 (
            .O(N__84312),
            .I(N__84309));
    Span4Mux_v I__20384 (
            .O(N__84309),
            .I(N__84306));
    Odrv4 I__20383 (
            .O(N__84306),
            .I(\pid_front.O_24 ));
    CascadeMux I__20382 (
            .O(N__84303),
            .I(N__84297));
    InMux I__20381 (
            .O(N__84302),
            .I(N__84284));
    InMux I__20380 (
            .O(N__84301),
            .I(N__84281));
    InMux I__20379 (
            .O(N__84300),
            .I(N__84272));
    InMux I__20378 (
            .O(N__84297),
            .I(N__84272));
    InMux I__20377 (
            .O(N__84296),
            .I(N__84272));
    InMux I__20376 (
            .O(N__84295),
            .I(N__84272));
    InMux I__20375 (
            .O(N__84294),
            .I(N__84263));
    InMux I__20374 (
            .O(N__84293),
            .I(N__84263));
    InMux I__20373 (
            .O(N__84292),
            .I(N__84263));
    InMux I__20372 (
            .O(N__84291),
            .I(N__84263));
    InMux I__20371 (
            .O(N__84290),
            .I(N__84260));
    InMux I__20370 (
            .O(N__84289),
            .I(N__84253));
    InMux I__20369 (
            .O(N__84288),
            .I(N__84253));
    InMux I__20368 (
            .O(N__84287),
            .I(N__84253));
    LocalMux I__20367 (
            .O(N__84284),
            .I(N__84250));
    LocalMux I__20366 (
            .O(N__84281),
            .I(N__84245));
    LocalMux I__20365 (
            .O(N__84272),
            .I(N__84245));
    LocalMux I__20364 (
            .O(N__84263),
            .I(N__84240));
    LocalMux I__20363 (
            .O(N__84260),
            .I(N__84240));
    LocalMux I__20362 (
            .O(N__84253),
            .I(N__84237));
    Span4Mux_v I__20361 (
            .O(N__84250),
            .I(N__84234));
    Span4Mux_v I__20360 (
            .O(N__84245),
            .I(N__84229));
    Span4Mux_h I__20359 (
            .O(N__84240),
            .I(N__84229));
    Span4Mux_v I__20358 (
            .O(N__84237),
            .I(N__84226));
    Span4Mux_h I__20357 (
            .O(N__84234),
            .I(N__84221));
    Span4Mux_h I__20356 (
            .O(N__84229),
            .I(N__84221));
    Sp12to4 I__20355 (
            .O(N__84226),
            .I(N__84218));
    Span4Mux_h I__20354 (
            .O(N__84221),
            .I(N__84215));
    Span12Mux_h I__20353 (
            .O(N__84218),
            .I(N__84212));
    Span4Mux_h I__20352 (
            .O(N__84215),
            .I(N__84209));
    Odrv12 I__20351 (
            .O(N__84212),
            .I(\pid_front.error_d_regZ0Z_22 ));
    Odrv4 I__20350 (
            .O(N__84209),
            .I(\pid_front.error_d_regZ0Z_22 ));
    InMux I__20349 (
            .O(N__84204),
            .I(N__84201));
    LocalMux I__20348 (
            .O(N__84201),
            .I(N__84198));
    Odrv4 I__20347 (
            .O(N__84198),
            .I(\pid_front.O_18 ));
    InMux I__20346 (
            .O(N__84195),
            .I(N__84186));
    InMux I__20345 (
            .O(N__84194),
            .I(N__84186));
    InMux I__20344 (
            .O(N__84193),
            .I(N__84186));
    LocalMux I__20343 (
            .O(N__84186),
            .I(N__84183));
    Span4Mux_h I__20342 (
            .O(N__84183),
            .I(N__84180));
    Span4Mux_h I__20341 (
            .O(N__84180),
            .I(N__84177));
    Span4Mux_h I__20340 (
            .O(N__84177),
            .I(N__84174));
    Odrv4 I__20339 (
            .O(N__84174),
            .I(\pid_front.error_d_regZ0Z_16 ));
    InMux I__20338 (
            .O(N__84171),
            .I(N__84168));
    LocalMux I__20337 (
            .O(N__84168),
            .I(N__84165));
    Odrv4 I__20336 (
            .O(N__84165),
            .I(\pid_front.O_17 ));
    InMux I__20335 (
            .O(N__84162),
            .I(N__84153));
    InMux I__20334 (
            .O(N__84161),
            .I(N__84153));
    InMux I__20333 (
            .O(N__84160),
            .I(N__84153));
    LocalMux I__20332 (
            .O(N__84153),
            .I(N__84150));
    Sp12to4 I__20331 (
            .O(N__84150),
            .I(N__84147));
    Span12Mux_v I__20330 (
            .O(N__84147),
            .I(N__84144));
    Odrv12 I__20329 (
            .O(N__84144),
            .I(\pid_front.error_d_regZ0Z_15 ));
    InMux I__20328 (
            .O(N__84141),
            .I(N__84138));
    LocalMux I__20327 (
            .O(N__84138),
            .I(\pid_front.O_16 ));
    InMux I__20326 (
            .O(N__84135),
            .I(N__84126));
    InMux I__20325 (
            .O(N__84134),
            .I(N__84126));
    InMux I__20324 (
            .O(N__84133),
            .I(N__84126));
    LocalMux I__20323 (
            .O(N__84126),
            .I(N__84123));
    Span12Mux_h I__20322 (
            .O(N__84123),
            .I(N__84120));
    Span12Mux_h I__20321 (
            .O(N__84120),
            .I(N__84117));
    Odrv12 I__20320 (
            .O(N__84117),
            .I(\pid_front.error_d_regZ0Z_14 ));
    ClkMux I__20319 (
            .O(N__84114),
            .I(N__83214));
    ClkMux I__20318 (
            .O(N__84113),
            .I(N__83214));
    ClkMux I__20317 (
            .O(N__84112),
            .I(N__83214));
    ClkMux I__20316 (
            .O(N__84111),
            .I(N__83214));
    ClkMux I__20315 (
            .O(N__84110),
            .I(N__83214));
    ClkMux I__20314 (
            .O(N__84109),
            .I(N__83214));
    ClkMux I__20313 (
            .O(N__84108),
            .I(N__83214));
    ClkMux I__20312 (
            .O(N__84107),
            .I(N__83214));
    ClkMux I__20311 (
            .O(N__84106),
            .I(N__83214));
    ClkMux I__20310 (
            .O(N__84105),
            .I(N__83214));
    ClkMux I__20309 (
            .O(N__84104),
            .I(N__83214));
    ClkMux I__20308 (
            .O(N__84103),
            .I(N__83214));
    ClkMux I__20307 (
            .O(N__84102),
            .I(N__83214));
    ClkMux I__20306 (
            .O(N__84101),
            .I(N__83214));
    ClkMux I__20305 (
            .O(N__84100),
            .I(N__83214));
    ClkMux I__20304 (
            .O(N__84099),
            .I(N__83214));
    ClkMux I__20303 (
            .O(N__84098),
            .I(N__83214));
    ClkMux I__20302 (
            .O(N__84097),
            .I(N__83214));
    ClkMux I__20301 (
            .O(N__84096),
            .I(N__83214));
    ClkMux I__20300 (
            .O(N__84095),
            .I(N__83214));
    ClkMux I__20299 (
            .O(N__84094),
            .I(N__83214));
    ClkMux I__20298 (
            .O(N__84093),
            .I(N__83214));
    ClkMux I__20297 (
            .O(N__84092),
            .I(N__83214));
    ClkMux I__20296 (
            .O(N__84091),
            .I(N__83214));
    ClkMux I__20295 (
            .O(N__84090),
            .I(N__83214));
    ClkMux I__20294 (
            .O(N__84089),
            .I(N__83214));
    ClkMux I__20293 (
            .O(N__84088),
            .I(N__83214));
    ClkMux I__20292 (
            .O(N__84087),
            .I(N__83214));
    ClkMux I__20291 (
            .O(N__84086),
            .I(N__83214));
    ClkMux I__20290 (
            .O(N__84085),
            .I(N__83214));
    ClkMux I__20289 (
            .O(N__84084),
            .I(N__83214));
    ClkMux I__20288 (
            .O(N__84083),
            .I(N__83214));
    ClkMux I__20287 (
            .O(N__84082),
            .I(N__83214));
    ClkMux I__20286 (
            .O(N__84081),
            .I(N__83214));
    ClkMux I__20285 (
            .O(N__84080),
            .I(N__83214));
    ClkMux I__20284 (
            .O(N__84079),
            .I(N__83214));
    ClkMux I__20283 (
            .O(N__84078),
            .I(N__83214));
    ClkMux I__20282 (
            .O(N__84077),
            .I(N__83214));
    ClkMux I__20281 (
            .O(N__84076),
            .I(N__83214));
    ClkMux I__20280 (
            .O(N__84075),
            .I(N__83214));
    ClkMux I__20279 (
            .O(N__84074),
            .I(N__83214));
    ClkMux I__20278 (
            .O(N__84073),
            .I(N__83214));
    ClkMux I__20277 (
            .O(N__84072),
            .I(N__83214));
    ClkMux I__20276 (
            .O(N__84071),
            .I(N__83214));
    ClkMux I__20275 (
            .O(N__84070),
            .I(N__83214));
    ClkMux I__20274 (
            .O(N__84069),
            .I(N__83214));
    ClkMux I__20273 (
            .O(N__84068),
            .I(N__83214));
    ClkMux I__20272 (
            .O(N__84067),
            .I(N__83214));
    ClkMux I__20271 (
            .O(N__84066),
            .I(N__83214));
    ClkMux I__20270 (
            .O(N__84065),
            .I(N__83214));
    ClkMux I__20269 (
            .O(N__84064),
            .I(N__83214));
    ClkMux I__20268 (
            .O(N__84063),
            .I(N__83214));
    ClkMux I__20267 (
            .O(N__84062),
            .I(N__83214));
    ClkMux I__20266 (
            .O(N__84061),
            .I(N__83214));
    ClkMux I__20265 (
            .O(N__84060),
            .I(N__83214));
    ClkMux I__20264 (
            .O(N__84059),
            .I(N__83214));
    ClkMux I__20263 (
            .O(N__84058),
            .I(N__83214));
    ClkMux I__20262 (
            .O(N__84057),
            .I(N__83214));
    ClkMux I__20261 (
            .O(N__84056),
            .I(N__83214));
    ClkMux I__20260 (
            .O(N__84055),
            .I(N__83214));
    ClkMux I__20259 (
            .O(N__84054),
            .I(N__83214));
    ClkMux I__20258 (
            .O(N__84053),
            .I(N__83214));
    ClkMux I__20257 (
            .O(N__84052),
            .I(N__83214));
    ClkMux I__20256 (
            .O(N__84051),
            .I(N__83214));
    ClkMux I__20255 (
            .O(N__84050),
            .I(N__83214));
    ClkMux I__20254 (
            .O(N__84049),
            .I(N__83214));
    ClkMux I__20253 (
            .O(N__84048),
            .I(N__83214));
    ClkMux I__20252 (
            .O(N__84047),
            .I(N__83214));
    ClkMux I__20251 (
            .O(N__84046),
            .I(N__83214));
    ClkMux I__20250 (
            .O(N__84045),
            .I(N__83214));
    ClkMux I__20249 (
            .O(N__84044),
            .I(N__83214));
    ClkMux I__20248 (
            .O(N__84043),
            .I(N__83214));
    ClkMux I__20247 (
            .O(N__84042),
            .I(N__83214));
    ClkMux I__20246 (
            .O(N__84041),
            .I(N__83214));
    ClkMux I__20245 (
            .O(N__84040),
            .I(N__83214));
    ClkMux I__20244 (
            .O(N__84039),
            .I(N__83214));
    ClkMux I__20243 (
            .O(N__84038),
            .I(N__83214));
    ClkMux I__20242 (
            .O(N__84037),
            .I(N__83214));
    ClkMux I__20241 (
            .O(N__84036),
            .I(N__83214));
    ClkMux I__20240 (
            .O(N__84035),
            .I(N__83214));
    ClkMux I__20239 (
            .O(N__84034),
            .I(N__83214));
    ClkMux I__20238 (
            .O(N__84033),
            .I(N__83214));
    ClkMux I__20237 (
            .O(N__84032),
            .I(N__83214));
    ClkMux I__20236 (
            .O(N__84031),
            .I(N__83214));
    ClkMux I__20235 (
            .O(N__84030),
            .I(N__83214));
    ClkMux I__20234 (
            .O(N__84029),
            .I(N__83214));
    ClkMux I__20233 (
            .O(N__84028),
            .I(N__83214));
    ClkMux I__20232 (
            .O(N__84027),
            .I(N__83214));
    ClkMux I__20231 (
            .O(N__84026),
            .I(N__83214));
    ClkMux I__20230 (
            .O(N__84025),
            .I(N__83214));
    ClkMux I__20229 (
            .O(N__84024),
            .I(N__83214));
    ClkMux I__20228 (
            .O(N__84023),
            .I(N__83214));
    ClkMux I__20227 (
            .O(N__84022),
            .I(N__83214));
    ClkMux I__20226 (
            .O(N__84021),
            .I(N__83214));
    ClkMux I__20225 (
            .O(N__84020),
            .I(N__83214));
    ClkMux I__20224 (
            .O(N__84019),
            .I(N__83214));
    ClkMux I__20223 (
            .O(N__84018),
            .I(N__83214));
    ClkMux I__20222 (
            .O(N__84017),
            .I(N__83214));
    ClkMux I__20221 (
            .O(N__84016),
            .I(N__83214));
    ClkMux I__20220 (
            .O(N__84015),
            .I(N__83214));
    ClkMux I__20219 (
            .O(N__84014),
            .I(N__83214));
    ClkMux I__20218 (
            .O(N__84013),
            .I(N__83214));
    ClkMux I__20217 (
            .O(N__84012),
            .I(N__83214));
    ClkMux I__20216 (
            .O(N__84011),
            .I(N__83214));
    ClkMux I__20215 (
            .O(N__84010),
            .I(N__83214));
    ClkMux I__20214 (
            .O(N__84009),
            .I(N__83214));
    ClkMux I__20213 (
            .O(N__84008),
            .I(N__83214));
    ClkMux I__20212 (
            .O(N__84007),
            .I(N__83214));
    ClkMux I__20211 (
            .O(N__84006),
            .I(N__83214));
    ClkMux I__20210 (
            .O(N__84005),
            .I(N__83214));
    ClkMux I__20209 (
            .O(N__84004),
            .I(N__83214));
    ClkMux I__20208 (
            .O(N__84003),
            .I(N__83214));
    ClkMux I__20207 (
            .O(N__84002),
            .I(N__83214));
    ClkMux I__20206 (
            .O(N__84001),
            .I(N__83214));
    ClkMux I__20205 (
            .O(N__84000),
            .I(N__83214));
    ClkMux I__20204 (
            .O(N__83999),
            .I(N__83214));
    ClkMux I__20203 (
            .O(N__83998),
            .I(N__83214));
    ClkMux I__20202 (
            .O(N__83997),
            .I(N__83214));
    ClkMux I__20201 (
            .O(N__83996),
            .I(N__83214));
    ClkMux I__20200 (
            .O(N__83995),
            .I(N__83214));
    ClkMux I__20199 (
            .O(N__83994),
            .I(N__83214));
    ClkMux I__20198 (
            .O(N__83993),
            .I(N__83214));
    ClkMux I__20197 (
            .O(N__83992),
            .I(N__83214));
    ClkMux I__20196 (
            .O(N__83991),
            .I(N__83214));
    ClkMux I__20195 (
            .O(N__83990),
            .I(N__83214));
    ClkMux I__20194 (
            .O(N__83989),
            .I(N__83214));
    ClkMux I__20193 (
            .O(N__83988),
            .I(N__83214));
    ClkMux I__20192 (
            .O(N__83987),
            .I(N__83214));
    ClkMux I__20191 (
            .O(N__83986),
            .I(N__83214));
    ClkMux I__20190 (
            .O(N__83985),
            .I(N__83214));
    ClkMux I__20189 (
            .O(N__83984),
            .I(N__83214));
    ClkMux I__20188 (
            .O(N__83983),
            .I(N__83214));
    ClkMux I__20187 (
            .O(N__83982),
            .I(N__83214));
    ClkMux I__20186 (
            .O(N__83981),
            .I(N__83214));
    ClkMux I__20185 (
            .O(N__83980),
            .I(N__83214));
    ClkMux I__20184 (
            .O(N__83979),
            .I(N__83214));
    ClkMux I__20183 (
            .O(N__83978),
            .I(N__83214));
    ClkMux I__20182 (
            .O(N__83977),
            .I(N__83214));
    ClkMux I__20181 (
            .O(N__83976),
            .I(N__83214));
    ClkMux I__20180 (
            .O(N__83975),
            .I(N__83214));
    ClkMux I__20179 (
            .O(N__83974),
            .I(N__83214));
    ClkMux I__20178 (
            .O(N__83973),
            .I(N__83214));
    ClkMux I__20177 (
            .O(N__83972),
            .I(N__83214));
    ClkMux I__20176 (
            .O(N__83971),
            .I(N__83214));
    ClkMux I__20175 (
            .O(N__83970),
            .I(N__83214));
    ClkMux I__20174 (
            .O(N__83969),
            .I(N__83214));
    ClkMux I__20173 (
            .O(N__83968),
            .I(N__83214));
    ClkMux I__20172 (
            .O(N__83967),
            .I(N__83214));
    ClkMux I__20171 (
            .O(N__83966),
            .I(N__83214));
    ClkMux I__20170 (
            .O(N__83965),
            .I(N__83214));
    ClkMux I__20169 (
            .O(N__83964),
            .I(N__83214));
    ClkMux I__20168 (
            .O(N__83963),
            .I(N__83214));
    ClkMux I__20167 (
            .O(N__83962),
            .I(N__83214));
    ClkMux I__20166 (
            .O(N__83961),
            .I(N__83214));
    ClkMux I__20165 (
            .O(N__83960),
            .I(N__83214));
    ClkMux I__20164 (
            .O(N__83959),
            .I(N__83214));
    ClkMux I__20163 (
            .O(N__83958),
            .I(N__83214));
    ClkMux I__20162 (
            .O(N__83957),
            .I(N__83214));
    ClkMux I__20161 (
            .O(N__83956),
            .I(N__83214));
    ClkMux I__20160 (
            .O(N__83955),
            .I(N__83214));
    ClkMux I__20159 (
            .O(N__83954),
            .I(N__83214));
    ClkMux I__20158 (
            .O(N__83953),
            .I(N__83214));
    ClkMux I__20157 (
            .O(N__83952),
            .I(N__83214));
    ClkMux I__20156 (
            .O(N__83951),
            .I(N__83214));
    ClkMux I__20155 (
            .O(N__83950),
            .I(N__83214));
    ClkMux I__20154 (
            .O(N__83949),
            .I(N__83214));
    ClkMux I__20153 (
            .O(N__83948),
            .I(N__83214));
    ClkMux I__20152 (
            .O(N__83947),
            .I(N__83214));
    ClkMux I__20151 (
            .O(N__83946),
            .I(N__83214));
    ClkMux I__20150 (
            .O(N__83945),
            .I(N__83214));
    ClkMux I__20149 (
            .O(N__83944),
            .I(N__83214));
    ClkMux I__20148 (
            .O(N__83943),
            .I(N__83214));
    ClkMux I__20147 (
            .O(N__83942),
            .I(N__83214));
    ClkMux I__20146 (
            .O(N__83941),
            .I(N__83214));
    ClkMux I__20145 (
            .O(N__83940),
            .I(N__83214));
    ClkMux I__20144 (
            .O(N__83939),
            .I(N__83214));
    ClkMux I__20143 (
            .O(N__83938),
            .I(N__83214));
    ClkMux I__20142 (
            .O(N__83937),
            .I(N__83214));
    ClkMux I__20141 (
            .O(N__83936),
            .I(N__83214));
    ClkMux I__20140 (
            .O(N__83935),
            .I(N__83214));
    ClkMux I__20139 (
            .O(N__83934),
            .I(N__83214));
    ClkMux I__20138 (
            .O(N__83933),
            .I(N__83214));
    ClkMux I__20137 (
            .O(N__83932),
            .I(N__83214));
    ClkMux I__20136 (
            .O(N__83931),
            .I(N__83214));
    ClkMux I__20135 (
            .O(N__83930),
            .I(N__83214));
    ClkMux I__20134 (
            .O(N__83929),
            .I(N__83214));
    ClkMux I__20133 (
            .O(N__83928),
            .I(N__83214));
    ClkMux I__20132 (
            .O(N__83927),
            .I(N__83214));
    ClkMux I__20131 (
            .O(N__83926),
            .I(N__83214));
    ClkMux I__20130 (
            .O(N__83925),
            .I(N__83214));
    ClkMux I__20129 (
            .O(N__83924),
            .I(N__83214));
    ClkMux I__20128 (
            .O(N__83923),
            .I(N__83214));
    ClkMux I__20127 (
            .O(N__83922),
            .I(N__83214));
    ClkMux I__20126 (
            .O(N__83921),
            .I(N__83214));
    ClkMux I__20125 (
            .O(N__83920),
            .I(N__83214));
    ClkMux I__20124 (
            .O(N__83919),
            .I(N__83214));
    ClkMux I__20123 (
            .O(N__83918),
            .I(N__83214));
    ClkMux I__20122 (
            .O(N__83917),
            .I(N__83214));
    ClkMux I__20121 (
            .O(N__83916),
            .I(N__83214));
    ClkMux I__20120 (
            .O(N__83915),
            .I(N__83214));
    ClkMux I__20119 (
            .O(N__83914),
            .I(N__83214));
    ClkMux I__20118 (
            .O(N__83913),
            .I(N__83214));
    ClkMux I__20117 (
            .O(N__83912),
            .I(N__83214));
    ClkMux I__20116 (
            .O(N__83911),
            .I(N__83214));
    ClkMux I__20115 (
            .O(N__83910),
            .I(N__83214));
    ClkMux I__20114 (
            .O(N__83909),
            .I(N__83214));
    ClkMux I__20113 (
            .O(N__83908),
            .I(N__83214));
    ClkMux I__20112 (
            .O(N__83907),
            .I(N__83214));
    ClkMux I__20111 (
            .O(N__83906),
            .I(N__83214));
    ClkMux I__20110 (
            .O(N__83905),
            .I(N__83214));
    ClkMux I__20109 (
            .O(N__83904),
            .I(N__83214));
    ClkMux I__20108 (
            .O(N__83903),
            .I(N__83214));
    ClkMux I__20107 (
            .O(N__83902),
            .I(N__83214));
    ClkMux I__20106 (
            .O(N__83901),
            .I(N__83214));
    ClkMux I__20105 (
            .O(N__83900),
            .I(N__83214));
    ClkMux I__20104 (
            .O(N__83899),
            .I(N__83214));
    ClkMux I__20103 (
            .O(N__83898),
            .I(N__83214));
    ClkMux I__20102 (
            .O(N__83897),
            .I(N__83214));
    ClkMux I__20101 (
            .O(N__83896),
            .I(N__83214));
    ClkMux I__20100 (
            .O(N__83895),
            .I(N__83214));
    ClkMux I__20099 (
            .O(N__83894),
            .I(N__83214));
    ClkMux I__20098 (
            .O(N__83893),
            .I(N__83214));
    ClkMux I__20097 (
            .O(N__83892),
            .I(N__83214));
    ClkMux I__20096 (
            .O(N__83891),
            .I(N__83214));
    ClkMux I__20095 (
            .O(N__83890),
            .I(N__83214));
    ClkMux I__20094 (
            .O(N__83889),
            .I(N__83214));
    ClkMux I__20093 (
            .O(N__83888),
            .I(N__83214));
    ClkMux I__20092 (
            .O(N__83887),
            .I(N__83214));
    ClkMux I__20091 (
            .O(N__83886),
            .I(N__83214));
    ClkMux I__20090 (
            .O(N__83885),
            .I(N__83214));
    ClkMux I__20089 (
            .O(N__83884),
            .I(N__83214));
    ClkMux I__20088 (
            .O(N__83883),
            .I(N__83214));
    ClkMux I__20087 (
            .O(N__83882),
            .I(N__83214));
    ClkMux I__20086 (
            .O(N__83881),
            .I(N__83214));
    ClkMux I__20085 (
            .O(N__83880),
            .I(N__83214));
    ClkMux I__20084 (
            .O(N__83879),
            .I(N__83214));
    ClkMux I__20083 (
            .O(N__83878),
            .I(N__83214));
    ClkMux I__20082 (
            .O(N__83877),
            .I(N__83214));
    ClkMux I__20081 (
            .O(N__83876),
            .I(N__83214));
    ClkMux I__20080 (
            .O(N__83875),
            .I(N__83214));
    ClkMux I__20079 (
            .O(N__83874),
            .I(N__83214));
    ClkMux I__20078 (
            .O(N__83873),
            .I(N__83214));
    ClkMux I__20077 (
            .O(N__83872),
            .I(N__83214));
    ClkMux I__20076 (
            .O(N__83871),
            .I(N__83214));
    ClkMux I__20075 (
            .O(N__83870),
            .I(N__83214));
    ClkMux I__20074 (
            .O(N__83869),
            .I(N__83214));
    ClkMux I__20073 (
            .O(N__83868),
            .I(N__83214));
    ClkMux I__20072 (
            .O(N__83867),
            .I(N__83214));
    ClkMux I__20071 (
            .O(N__83866),
            .I(N__83214));
    ClkMux I__20070 (
            .O(N__83865),
            .I(N__83214));
    ClkMux I__20069 (
            .O(N__83864),
            .I(N__83214));
    ClkMux I__20068 (
            .O(N__83863),
            .I(N__83214));
    ClkMux I__20067 (
            .O(N__83862),
            .I(N__83214));
    ClkMux I__20066 (
            .O(N__83861),
            .I(N__83214));
    ClkMux I__20065 (
            .O(N__83860),
            .I(N__83214));
    ClkMux I__20064 (
            .O(N__83859),
            .I(N__83214));
    ClkMux I__20063 (
            .O(N__83858),
            .I(N__83214));
    ClkMux I__20062 (
            .O(N__83857),
            .I(N__83214));
    ClkMux I__20061 (
            .O(N__83856),
            .I(N__83214));
    ClkMux I__20060 (
            .O(N__83855),
            .I(N__83214));
    ClkMux I__20059 (
            .O(N__83854),
            .I(N__83214));
    ClkMux I__20058 (
            .O(N__83853),
            .I(N__83214));
    ClkMux I__20057 (
            .O(N__83852),
            .I(N__83214));
    ClkMux I__20056 (
            .O(N__83851),
            .I(N__83214));
    ClkMux I__20055 (
            .O(N__83850),
            .I(N__83214));
    ClkMux I__20054 (
            .O(N__83849),
            .I(N__83214));
    ClkMux I__20053 (
            .O(N__83848),
            .I(N__83214));
    ClkMux I__20052 (
            .O(N__83847),
            .I(N__83214));
    ClkMux I__20051 (
            .O(N__83846),
            .I(N__83214));
    ClkMux I__20050 (
            .O(N__83845),
            .I(N__83214));
    ClkMux I__20049 (
            .O(N__83844),
            .I(N__83214));
    ClkMux I__20048 (
            .O(N__83843),
            .I(N__83214));
    ClkMux I__20047 (
            .O(N__83842),
            .I(N__83214));
    ClkMux I__20046 (
            .O(N__83841),
            .I(N__83214));
    ClkMux I__20045 (
            .O(N__83840),
            .I(N__83214));
    ClkMux I__20044 (
            .O(N__83839),
            .I(N__83214));
    ClkMux I__20043 (
            .O(N__83838),
            .I(N__83214));
    ClkMux I__20042 (
            .O(N__83837),
            .I(N__83214));
    ClkMux I__20041 (
            .O(N__83836),
            .I(N__83214));
    ClkMux I__20040 (
            .O(N__83835),
            .I(N__83214));
    ClkMux I__20039 (
            .O(N__83834),
            .I(N__83214));
    ClkMux I__20038 (
            .O(N__83833),
            .I(N__83214));
    ClkMux I__20037 (
            .O(N__83832),
            .I(N__83214));
    ClkMux I__20036 (
            .O(N__83831),
            .I(N__83214));
    ClkMux I__20035 (
            .O(N__83830),
            .I(N__83214));
    ClkMux I__20034 (
            .O(N__83829),
            .I(N__83214));
    ClkMux I__20033 (
            .O(N__83828),
            .I(N__83214));
    ClkMux I__20032 (
            .O(N__83827),
            .I(N__83214));
    ClkMux I__20031 (
            .O(N__83826),
            .I(N__83214));
    ClkMux I__20030 (
            .O(N__83825),
            .I(N__83214));
    ClkMux I__20029 (
            .O(N__83824),
            .I(N__83214));
    ClkMux I__20028 (
            .O(N__83823),
            .I(N__83214));
    ClkMux I__20027 (
            .O(N__83822),
            .I(N__83214));
    ClkMux I__20026 (
            .O(N__83821),
            .I(N__83214));
    ClkMux I__20025 (
            .O(N__83820),
            .I(N__83214));
    ClkMux I__20024 (
            .O(N__83819),
            .I(N__83214));
    ClkMux I__20023 (
            .O(N__83818),
            .I(N__83214));
    ClkMux I__20022 (
            .O(N__83817),
            .I(N__83214));
    ClkMux I__20021 (
            .O(N__83816),
            .I(N__83214));
    ClkMux I__20020 (
            .O(N__83815),
            .I(N__83214));
    GlobalMux I__20019 (
            .O(N__83214),
            .I(N__83211));
    gio2CtrlBuf I__20018 (
            .O(N__83211),
            .I(clk_system_pll_g));
    CEMux I__20017 (
            .O(N__83208),
            .I(N__83205));
    LocalMux I__20016 (
            .O(N__83205),
            .I(N__83198));
    CEMux I__20015 (
            .O(N__83204),
            .I(N__83195));
    CEMux I__20014 (
            .O(N__83203),
            .I(N__83192));
    CEMux I__20013 (
            .O(N__83202),
            .I(N__83189));
    CEMux I__20012 (
            .O(N__83201),
            .I(N__83185));
    Span4Mux_v I__20011 (
            .O(N__83198),
            .I(N__83175));
    LocalMux I__20010 (
            .O(N__83195),
            .I(N__83175));
    LocalMux I__20009 (
            .O(N__83192),
            .I(N__83175));
    LocalMux I__20008 (
            .O(N__83189),
            .I(N__83172));
    CEMux I__20007 (
            .O(N__83188),
            .I(N__83169));
    LocalMux I__20006 (
            .O(N__83185),
            .I(N__83166));
    CEMux I__20005 (
            .O(N__83184),
            .I(N__83163));
    CEMux I__20004 (
            .O(N__83183),
            .I(N__83160));
    CEMux I__20003 (
            .O(N__83182),
            .I(N__83157));
    Span4Mux_v I__20002 (
            .O(N__83175),
            .I(N__83149));
    Span4Mux_v I__20001 (
            .O(N__83172),
            .I(N__83149));
    LocalMux I__20000 (
            .O(N__83169),
            .I(N__83149));
    Span4Mux_v I__19999 (
            .O(N__83166),
            .I(N__83146));
    LocalMux I__19998 (
            .O(N__83163),
            .I(N__83141));
    LocalMux I__19997 (
            .O(N__83160),
            .I(N__83141));
    LocalMux I__19996 (
            .O(N__83157),
            .I(N__83138));
    CEMux I__19995 (
            .O(N__83156),
            .I(N__83135));
    Span4Mux_h I__19994 (
            .O(N__83149),
            .I(N__83128));
    Span4Mux_h I__19993 (
            .O(N__83146),
            .I(N__83119));
    Span4Mux_v I__19992 (
            .O(N__83141),
            .I(N__83119));
    Span4Mux_v I__19991 (
            .O(N__83138),
            .I(N__83119));
    LocalMux I__19990 (
            .O(N__83135),
            .I(N__83119));
    CEMux I__19989 (
            .O(N__83134),
            .I(N__83116));
    CEMux I__19988 (
            .O(N__83133),
            .I(N__83113));
    CEMux I__19987 (
            .O(N__83132),
            .I(N__83110));
    CEMux I__19986 (
            .O(N__83131),
            .I(N__83107));
    Span4Mux_h I__19985 (
            .O(N__83128),
            .I(N__83103));
    Span4Mux_h I__19984 (
            .O(N__83119),
            .I(N__83100));
    LocalMux I__19983 (
            .O(N__83116),
            .I(N__83097));
    LocalMux I__19982 (
            .O(N__83113),
            .I(N__83094));
    LocalMux I__19981 (
            .O(N__83110),
            .I(N__83091));
    LocalMux I__19980 (
            .O(N__83107),
            .I(N__83087));
    CEMux I__19979 (
            .O(N__83106),
            .I(N__83084));
    Span4Mux_h I__19978 (
            .O(N__83103),
            .I(N__83077));
    Span4Mux_h I__19977 (
            .O(N__83100),
            .I(N__83077));
    Span4Mux_v I__19976 (
            .O(N__83097),
            .I(N__83077));
    Span4Mux_h I__19975 (
            .O(N__83094),
            .I(N__83072));
    Span4Mux_h I__19974 (
            .O(N__83091),
            .I(N__83072));
    CEMux I__19973 (
            .O(N__83090),
            .I(N__83069));
    Span4Mux_h I__19972 (
            .O(N__83087),
            .I(N__83066));
    LocalMux I__19971 (
            .O(N__83084),
            .I(N__83063));
    Span4Mux_h I__19970 (
            .O(N__83077),
            .I(N__83056));
    Span4Mux_h I__19969 (
            .O(N__83072),
            .I(N__83056));
    LocalMux I__19968 (
            .O(N__83069),
            .I(N__83056));
    Span4Mux_h I__19967 (
            .O(N__83066),
            .I(N__83051));
    Span4Mux_v I__19966 (
            .O(N__83063),
            .I(N__83051));
    Span4Mux_v I__19965 (
            .O(N__83056),
            .I(N__83048));
    Odrv4 I__19964 (
            .O(N__83051),
            .I(\pid_front.N_429_0 ));
    Odrv4 I__19963 (
            .O(N__83048),
            .I(\pid_front.N_429_0 ));
    InMux I__19962 (
            .O(N__83043),
            .I(N__82990));
    InMux I__19961 (
            .O(N__83042),
            .I(N__82990));
    InMux I__19960 (
            .O(N__83041),
            .I(N__82990));
    InMux I__19959 (
            .O(N__83040),
            .I(N__82990));
    InMux I__19958 (
            .O(N__83039),
            .I(N__82990));
    InMux I__19957 (
            .O(N__83038),
            .I(N__82985));
    InMux I__19956 (
            .O(N__83037),
            .I(N__82985));
    InMux I__19955 (
            .O(N__83036),
            .I(N__82968));
    InMux I__19954 (
            .O(N__83035),
            .I(N__82968));
    InMux I__19953 (
            .O(N__83034),
            .I(N__82968));
    InMux I__19952 (
            .O(N__83033),
            .I(N__82968));
    InMux I__19951 (
            .O(N__83032),
            .I(N__82968));
    InMux I__19950 (
            .O(N__83031),
            .I(N__82968));
    InMux I__19949 (
            .O(N__83030),
            .I(N__82968));
    InMux I__19948 (
            .O(N__83029),
            .I(N__82968));
    InMux I__19947 (
            .O(N__83028),
            .I(N__82965));
    InMux I__19946 (
            .O(N__83027),
            .I(N__82962));
    InMux I__19945 (
            .O(N__83026),
            .I(N__82959));
    InMux I__19944 (
            .O(N__83025),
            .I(N__82956));
    InMux I__19943 (
            .O(N__83024),
            .I(N__82951));
    InMux I__19942 (
            .O(N__83023),
            .I(N__82951));
    InMux I__19941 (
            .O(N__83022),
            .I(N__82936));
    InMux I__19940 (
            .O(N__83021),
            .I(N__82936));
    InMux I__19939 (
            .O(N__83020),
            .I(N__82936));
    InMux I__19938 (
            .O(N__83019),
            .I(N__82936));
    InMux I__19937 (
            .O(N__83018),
            .I(N__82936));
    InMux I__19936 (
            .O(N__83017),
            .I(N__82936));
    InMux I__19935 (
            .O(N__83016),
            .I(N__82936));
    InMux I__19934 (
            .O(N__83015),
            .I(N__82933));
    InMux I__19933 (
            .O(N__83014),
            .I(N__82928));
    InMux I__19932 (
            .O(N__83013),
            .I(N__82928));
    InMux I__19931 (
            .O(N__83012),
            .I(N__82925));
    InMux I__19930 (
            .O(N__83011),
            .I(N__82916));
    InMux I__19929 (
            .O(N__83010),
            .I(N__82916));
    InMux I__19928 (
            .O(N__83009),
            .I(N__82916));
    InMux I__19927 (
            .O(N__83008),
            .I(N__82916));
    InMux I__19926 (
            .O(N__83007),
            .I(N__82913));
    InMux I__19925 (
            .O(N__83006),
            .I(N__82910));
    InMux I__19924 (
            .O(N__83005),
            .I(N__82907));
    InMux I__19923 (
            .O(N__83004),
            .I(N__82904));
    InMux I__19922 (
            .O(N__83003),
            .I(N__82901));
    InMux I__19921 (
            .O(N__83002),
            .I(N__82898));
    InMux I__19920 (
            .O(N__83001),
            .I(N__82895));
    LocalMux I__19919 (
            .O(N__82990),
            .I(N__82846));
    LocalMux I__19918 (
            .O(N__82985),
            .I(N__82843));
    LocalMux I__19917 (
            .O(N__82968),
            .I(N__82840));
    LocalMux I__19916 (
            .O(N__82965),
            .I(N__82837));
    LocalMux I__19915 (
            .O(N__82962),
            .I(N__82834));
    LocalMux I__19914 (
            .O(N__82959),
            .I(N__82831));
    LocalMux I__19913 (
            .O(N__82956),
            .I(N__82828));
    LocalMux I__19912 (
            .O(N__82951),
            .I(N__82825));
    LocalMux I__19911 (
            .O(N__82936),
            .I(N__82822));
    LocalMux I__19910 (
            .O(N__82933),
            .I(N__82819));
    LocalMux I__19909 (
            .O(N__82928),
            .I(N__82816));
    LocalMux I__19908 (
            .O(N__82925),
            .I(N__82813));
    LocalMux I__19907 (
            .O(N__82916),
            .I(N__82810));
    LocalMux I__19906 (
            .O(N__82913),
            .I(N__82807));
    LocalMux I__19905 (
            .O(N__82910),
            .I(N__82804));
    LocalMux I__19904 (
            .O(N__82907),
            .I(N__82801));
    LocalMux I__19903 (
            .O(N__82904),
            .I(N__82798));
    LocalMux I__19902 (
            .O(N__82901),
            .I(N__82795));
    LocalMux I__19901 (
            .O(N__82898),
            .I(N__82792));
    LocalMux I__19900 (
            .O(N__82895),
            .I(N__82789));
    SRMux I__19899 (
            .O(N__82894),
            .I(N__82656));
    SRMux I__19898 (
            .O(N__82893),
            .I(N__82656));
    SRMux I__19897 (
            .O(N__82892),
            .I(N__82656));
    SRMux I__19896 (
            .O(N__82891),
            .I(N__82656));
    SRMux I__19895 (
            .O(N__82890),
            .I(N__82656));
    SRMux I__19894 (
            .O(N__82889),
            .I(N__82656));
    SRMux I__19893 (
            .O(N__82888),
            .I(N__82656));
    SRMux I__19892 (
            .O(N__82887),
            .I(N__82656));
    SRMux I__19891 (
            .O(N__82886),
            .I(N__82656));
    SRMux I__19890 (
            .O(N__82885),
            .I(N__82656));
    SRMux I__19889 (
            .O(N__82884),
            .I(N__82656));
    SRMux I__19888 (
            .O(N__82883),
            .I(N__82656));
    SRMux I__19887 (
            .O(N__82882),
            .I(N__82656));
    SRMux I__19886 (
            .O(N__82881),
            .I(N__82656));
    SRMux I__19885 (
            .O(N__82880),
            .I(N__82656));
    SRMux I__19884 (
            .O(N__82879),
            .I(N__82656));
    SRMux I__19883 (
            .O(N__82878),
            .I(N__82656));
    SRMux I__19882 (
            .O(N__82877),
            .I(N__82656));
    SRMux I__19881 (
            .O(N__82876),
            .I(N__82656));
    SRMux I__19880 (
            .O(N__82875),
            .I(N__82656));
    SRMux I__19879 (
            .O(N__82874),
            .I(N__82656));
    SRMux I__19878 (
            .O(N__82873),
            .I(N__82656));
    SRMux I__19877 (
            .O(N__82872),
            .I(N__82656));
    SRMux I__19876 (
            .O(N__82871),
            .I(N__82656));
    SRMux I__19875 (
            .O(N__82870),
            .I(N__82656));
    SRMux I__19874 (
            .O(N__82869),
            .I(N__82656));
    SRMux I__19873 (
            .O(N__82868),
            .I(N__82656));
    SRMux I__19872 (
            .O(N__82867),
            .I(N__82656));
    SRMux I__19871 (
            .O(N__82866),
            .I(N__82656));
    SRMux I__19870 (
            .O(N__82865),
            .I(N__82656));
    SRMux I__19869 (
            .O(N__82864),
            .I(N__82656));
    SRMux I__19868 (
            .O(N__82863),
            .I(N__82656));
    SRMux I__19867 (
            .O(N__82862),
            .I(N__82656));
    SRMux I__19866 (
            .O(N__82861),
            .I(N__82656));
    SRMux I__19865 (
            .O(N__82860),
            .I(N__82656));
    SRMux I__19864 (
            .O(N__82859),
            .I(N__82656));
    SRMux I__19863 (
            .O(N__82858),
            .I(N__82656));
    SRMux I__19862 (
            .O(N__82857),
            .I(N__82656));
    SRMux I__19861 (
            .O(N__82856),
            .I(N__82656));
    SRMux I__19860 (
            .O(N__82855),
            .I(N__82656));
    SRMux I__19859 (
            .O(N__82854),
            .I(N__82656));
    SRMux I__19858 (
            .O(N__82853),
            .I(N__82656));
    SRMux I__19857 (
            .O(N__82852),
            .I(N__82656));
    SRMux I__19856 (
            .O(N__82851),
            .I(N__82656));
    SRMux I__19855 (
            .O(N__82850),
            .I(N__82656));
    SRMux I__19854 (
            .O(N__82849),
            .I(N__82656));
    Glb2LocalMux I__19853 (
            .O(N__82846),
            .I(N__82656));
    Glb2LocalMux I__19852 (
            .O(N__82843),
            .I(N__82656));
    Glb2LocalMux I__19851 (
            .O(N__82840),
            .I(N__82656));
    Glb2LocalMux I__19850 (
            .O(N__82837),
            .I(N__82656));
    Glb2LocalMux I__19849 (
            .O(N__82834),
            .I(N__82656));
    Glb2LocalMux I__19848 (
            .O(N__82831),
            .I(N__82656));
    Glb2LocalMux I__19847 (
            .O(N__82828),
            .I(N__82656));
    Glb2LocalMux I__19846 (
            .O(N__82825),
            .I(N__82656));
    Glb2LocalMux I__19845 (
            .O(N__82822),
            .I(N__82656));
    Glb2LocalMux I__19844 (
            .O(N__82819),
            .I(N__82656));
    Glb2LocalMux I__19843 (
            .O(N__82816),
            .I(N__82656));
    Glb2LocalMux I__19842 (
            .O(N__82813),
            .I(N__82656));
    Glb2LocalMux I__19841 (
            .O(N__82810),
            .I(N__82656));
    Glb2LocalMux I__19840 (
            .O(N__82807),
            .I(N__82656));
    Glb2LocalMux I__19839 (
            .O(N__82804),
            .I(N__82656));
    Glb2LocalMux I__19838 (
            .O(N__82801),
            .I(N__82656));
    Glb2LocalMux I__19837 (
            .O(N__82798),
            .I(N__82656));
    Glb2LocalMux I__19836 (
            .O(N__82795),
            .I(N__82656));
    Glb2LocalMux I__19835 (
            .O(N__82792),
            .I(N__82656));
    Glb2LocalMux I__19834 (
            .O(N__82789),
            .I(N__82656));
    GlobalMux I__19833 (
            .O(N__82656),
            .I(N__82653));
    gio2CtrlBuf I__19832 (
            .O(N__82653),
            .I(N_580_g));
    InMux I__19831 (
            .O(N__82650),
            .I(N__82647));
    LocalMux I__19830 (
            .O(N__82647),
            .I(\pid_side.O_1_14 ));
    InMux I__19829 (
            .O(N__82644),
            .I(N__82641));
    LocalMux I__19828 (
            .O(N__82641),
            .I(N__82637));
    InMux I__19827 (
            .O(N__82640),
            .I(N__82634));
    Span4Mux_h I__19826 (
            .O(N__82637),
            .I(N__82627));
    LocalMux I__19825 (
            .O(N__82634),
            .I(N__82627));
    InMux I__19824 (
            .O(N__82633),
            .I(N__82624));
    InMux I__19823 (
            .O(N__82632),
            .I(N__82621));
    Span4Mux_h I__19822 (
            .O(N__82627),
            .I(N__82614));
    LocalMux I__19821 (
            .O(N__82624),
            .I(N__82609));
    LocalMux I__19820 (
            .O(N__82621),
            .I(N__82609));
    InMux I__19819 (
            .O(N__82620),
            .I(N__82604));
    InMux I__19818 (
            .O(N__82619),
            .I(N__82604));
    InMux I__19817 (
            .O(N__82618),
            .I(N__82599));
    InMux I__19816 (
            .O(N__82617),
            .I(N__82599));
    Odrv4 I__19815 (
            .O(N__82614),
            .I(\pid_side.error_d_regZ0Z_12 ));
    Odrv4 I__19814 (
            .O(N__82609),
            .I(\pid_side.error_d_regZ0Z_12 ));
    LocalMux I__19813 (
            .O(N__82604),
            .I(\pid_side.error_d_regZ0Z_12 ));
    LocalMux I__19812 (
            .O(N__82599),
            .I(\pid_side.error_d_regZ0Z_12 ));
    InMux I__19811 (
            .O(N__82590),
            .I(N__82587));
    LocalMux I__19810 (
            .O(N__82587),
            .I(\pid_side.O_1_15 ));
    InMux I__19809 (
            .O(N__82584),
            .I(N__82579));
    InMux I__19808 (
            .O(N__82583),
            .I(N__82576));
    CascadeMux I__19807 (
            .O(N__82582),
            .I(N__82573));
    LocalMux I__19806 (
            .O(N__82579),
            .I(N__82569));
    LocalMux I__19805 (
            .O(N__82576),
            .I(N__82566));
    InMux I__19804 (
            .O(N__82573),
            .I(N__82561));
    InMux I__19803 (
            .O(N__82572),
            .I(N__82561));
    Span4Mux_h I__19802 (
            .O(N__82569),
            .I(N__82558));
    Span4Mux_v I__19801 (
            .O(N__82566),
            .I(N__82553));
    LocalMux I__19800 (
            .O(N__82561),
            .I(N__82553));
    Odrv4 I__19799 (
            .O(N__82558),
            .I(\pid_side.error_d_regZ0Z_13 ));
    Odrv4 I__19798 (
            .O(N__82553),
            .I(\pid_side.error_d_regZ0Z_13 ));
    InMux I__19797 (
            .O(N__82548),
            .I(N__82545));
    LocalMux I__19796 (
            .O(N__82545),
            .I(\pid_side.O_1_16 ));
    InMux I__19795 (
            .O(N__82542),
            .I(N__82536));
    InMux I__19794 (
            .O(N__82541),
            .I(N__82536));
    LocalMux I__19793 (
            .O(N__82536),
            .I(N__82532));
    InMux I__19792 (
            .O(N__82535),
            .I(N__82529));
    Span4Mux_v I__19791 (
            .O(N__82532),
            .I(N__82524));
    LocalMux I__19790 (
            .O(N__82529),
            .I(N__82524));
    Odrv4 I__19789 (
            .O(N__82524),
            .I(\pid_side.error_d_regZ0Z_14 ));
    InMux I__19788 (
            .O(N__82521),
            .I(N__82518));
    LocalMux I__19787 (
            .O(N__82518),
            .I(\pid_side.O_1_23 ));
    InMux I__19786 (
            .O(N__82515),
            .I(N__82506));
    InMux I__19785 (
            .O(N__82514),
            .I(N__82506));
    InMux I__19784 (
            .O(N__82513),
            .I(N__82506));
    LocalMux I__19783 (
            .O(N__82506),
            .I(N__82503));
    Span4Mux_h I__19782 (
            .O(N__82503),
            .I(N__82500));
    Span4Mux_h I__19781 (
            .O(N__82500),
            .I(N__82497));
    Odrv4 I__19780 (
            .O(N__82497),
            .I(\pid_side.error_d_regZ0Z_21 ));
    InMux I__19779 (
            .O(N__82494),
            .I(N__82491));
    LocalMux I__19778 (
            .O(N__82491),
            .I(\pid_side.O_1_22 ));
    InMux I__19777 (
            .O(N__82488),
            .I(N__82482));
    InMux I__19776 (
            .O(N__82487),
            .I(N__82482));
    LocalMux I__19775 (
            .O(N__82482),
            .I(N__82479));
    Span4Mux_h I__19774 (
            .O(N__82479),
            .I(N__82476));
    Span4Mux_h I__19773 (
            .O(N__82476),
            .I(N__82472));
    InMux I__19772 (
            .O(N__82475),
            .I(N__82469));
    Odrv4 I__19771 (
            .O(N__82472),
            .I(\pid_side.error_d_regZ0Z_20 ));
    LocalMux I__19770 (
            .O(N__82469),
            .I(\pid_side.error_d_regZ0Z_20 ));
    CEMux I__19769 (
            .O(N__82464),
            .I(N__82461));
    LocalMux I__19768 (
            .O(N__82461),
            .I(N__82448));
    CEMux I__19767 (
            .O(N__82460),
            .I(N__82445));
    CEMux I__19766 (
            .O(N__82459),
            .I(N__82442));
    CEMux I__19765 (
            .O(N__82458),
            .I(N__82439));
    CEMux I__19764 (
            .O(N__82457),
            .I(N__82436));
    CEMux I__19763 (
            .O(N__82456),
            .I(N__82433));
    CEMux I__19762 (
            .O(N__82455),
            .I(N__82428));
    CEMux I__19761 (
            .O(N__82454),
            .I(N__82425));
    CEMux I__19760 (
            .O(N__82453),
            .I(N__82422));
    CEMux I__19759 (
            .O(N__82452),
            .I(N__82419));
    CEMux I__19758 (
            .O(N__82451),
            .I(N__82416));
    Span4Mux_v I__19757 (
            .O(N__82448),
            .I(N__82409));
    LocalMux I__19756 (
            .O(N__82445),
            .I(N__82409));
    LocalMux I__19755 (
            .O(N__82442),
            .I(N__82406));
    LocalMux I__19754 (
            .O(N__82439),
            .I(N__82403));
    LocalMux I__19753 (
            .O(N__82436),
            .I(N__82400));
    LocalMux I__19752 (
            .O(N__82433),
            .I(N__82397));
    CEMux I__19751 (
            .O(N__82432),
            .I(N__82394));
    CEMux I__19750 (
            .O(N__82431),
            .I(N__82391));
    LocalMux I__19749 (
            .O(N__82428),
            .I(N__82386));
    LocalMux I__19748 (
            .O(N__82425),
            .I(N__82386));
    LocalMux I__19747 (
            .O(N__82422),
            .I(N__82383));
    LocalMux I__19746 (
            .O(N__82419),
            .I(N__82380));
    LocalMux I__19745 (
            .O(N__82416),
            .I(N__82377));
    CEMux I__19744 (
            .O(N__82415),
            .I(N__82374));
    CEMux I__19743 (
            .O(N__82414),
            .I(N__82371));
    Span4Mux_s2_h I__19742 (
            .O(N__82409),
            .I(N__82368));
    Span4Mux_v I__19741 (
            .O(N__82406),
            .I(N__82363));
    Span4Mux_v I__19740 (
            .O(N__82403),
            .I(N__82363));
    Span4Mux_h I__19739 (
            .O(N__82400),
            .I(N__82354));
    Span4Mux_v I__19738 (
            .O(N__82397),
            .I(N__82354));
    LocalMux I__19737 (
            .O(N__82394),
            .I(N__82354));
    LocalMux I__19736 (
            .O(N__82391),
            .I(N__82354));
    Span4Mux_v I__19735 (
            .O(N__82386),
            .I(N__82343));
    Span4Mux_v I__19734 (
            .O(N__82383),
            .I(N__82343));
    Span4Mux_s1_h I__19733 (
            .O(N__82380),
            .I(N__82343));
    Span4Mux_v I__19732 (
            .O(N__82377),
            .I(N__82343));
    LocalMux I__19731 (
            .O(N__82374),
            .I(N__82343));
    LocalMux I__19730 (
            .O(N__82371),
            .I(N__82340));
    Span4Mux_h I__19729 (
            .O(N__82368),
            .I(N__82337));
    Span4Mux_h I__19728 (
            .O(N__82363),
            .I(N__82332));
    Span4Mux_v I__19727 (
            .O(N__82354),
            .I(N__82332));
    Span4Mux_h I__19726 (
            .O(N__82343),
            .I(N__82327));
    Span4Mux_v I__19725 (
            .O(N__82340),
            .I(N__82327));
    Odrv4 I__19724 (
            .O(N__82337),
            .I(\pid_side.N_513_0 ));
    Odrv4 I__19723 (
            .O(N__82332),
            .I(\pid_side.N_513_0 ));
    Odrv4 I__19722 (
            .O(N__82327),
            .I(\pid_side.N_513_0 ));
    InMux I__19721 (
            .O(N__82320),
            .I(N__82317));
    LocalMux I__19720 (
            .O(N__82317),
            .I(N__82314));
    Span4Mux_v I__19719 (
            .O(N__82314),
            .I(N__82311));
    Odrv4 I__19718 (
            .O(N__82311),
            .I(\pid_front.O_10 ));
    InMux I__19717 (
            .O(N__82308),
            .I(N__82302));
    InMux I__19716 (
            .O(N__82307),
            .I(N__82302));
    LocalMux I__19715 (
            .O(N__82302),
            .I(N__82299));
    Span4Mux_h I__19714 (
            .O(N__82299),
            .I(N__82294));
    InMux I__19713 (
            .O(N__82298),
            .I(N__82289));
    InMux I__19712 (
            .O(N__82297),
            .I(N__82289));
    Span4Mux_h I__19711 (
            .O(N__82294),
            .I(N__82286));
    LocalMux I__19710 (
            .O(N__82289),
            .I(N__82283));
    Span4Mux_h I__19709 (
            .O(N__82286),
            .I(N__82280));
    Span12Mux_h I__19708 (
            .O(N__82283),
            .I(N__82277));
    Odrv4 I__19707 (
            .O(N__82280),
            .I(\pid_front.error_d_regZ0Z_8 ));
    Odrv12 I__19706 (
            .O(N__82277),
            .I(\pid_front.error_d_regZ0Z_8 ));
    InMux I__19705 (
            .O(N__82272),
            .I(N__82269));
    LocalMux I__19704 (
            .O(N__82269),
            .I(N__82266));
    Span4Mux_h I__19703 (
            .O(N__82266),
            .I(N__82263));
    Odrv4 I__19702 (
            .O(N__82263),
            .I(\pid_front.O_19 ));
    InMux I__19701 (
            .O(N__82260),
            .I(N__82251));
    InMux I__19700 (
            .O(N__82259),
            .I(N__82251));
    InMux I__19699 (
            .O(N__82258),
            .I(N__82251));
    LocalMux I__19698 (
            .O(N__82251),
            .I(N__82248));
    Span12Mux_v I__19697 (
            .O(N__82248),
            .I(N__82245));
    Span12Mux_h I__19696 (
            .O(N__82245),
            .I(N__82242));
    Odrv12 I__19695 (
            .O(N__82242),
            .I(\pid_front.error_d_regZ0Z_17 ));
    InMux I__19694 (
            .O(N__82239),
            .I(N__82236));
    LocalMux I__19693 (
            .O(N__82236),
            .I(N__82233));
    Odrv4 I__19692 (
            .O(N__82233),
            .I(\pid_front.O_20 ));
    InMux I__19691 (
            .O(N__82230),
            .I(N__82223));
    InMux I__19690 (
            .O(N__82229),
            .I(N__82223));
    InMux I__19689 (
            .O(N__82228),
            .I(N__82220));
    LocalMux I__19688 (
            .O(N__82223),
            .I(N__82217));
    LocalMux I__19687 (
            .O(N__82220),
            .I(N__82214));
    Span4Mux_h I__19686 (
            .O(N__82217),
            .I(N__82211));
    Span4Mux_h I__19685 (
            .O(N__82214),
            .I(N__82208));
    Span4Mux_h I__19684 (
            .O(N__82211),
            .I(N__82205));
    Span4Mux_h I__19683 (
            .O(N__82208),
            .I(N__82202));
    Span4Mux_h I__19682 (
            .O(N__82205),
            .I(N__82199));
    Span4Mux_h I__19681 (
            .O(N__82202),
            .I(N__82196));
    Odrv4 I__19680 (
            .O(N__82199),
            .I(\pid_front.error_d_regZ0Z_18 ));
    Odrv4 I__19679 (
            .O(N__82196),
            .I(\pid_front.error_d_regZ0Z_18 ));
    InMux I__19678 (
            .O(N__82191),
            .I(N__82187));
    InMux I__19677 (
            .O(N__82190),
            .I(N__82184));
    LocalMux I__19676 (
            .O(N__82187),
            .I(N__82179));
    LocalMux I__19675 (
            .O(N__82184),
            .I(N__82179));
    Span4Mux_v I__19674 (
            .O(N__82179),
            .I(N__82176));
    Odrv4 I__19673 (
            .O(N__82176),
            .I(\pid_side.error_p_regZ0Z_19 ));
    InMux I__19672 (
            .O(N__82173),
            .I(N__82169));
    InMux I__19671 (
            .O(N__82172),
            .I(N__82166));
    LocalMux I__19670 (
            .O(N__82169),
            .I(\pid_side.error_d_reg_prevZ0Z_19 ));
    LocalMux I__19669 (
            .O(N__82166),
            .I(\pid_side.error_d_reg_prevZ0Z_19 ));
    InMux I__19668 (
            .O(N__82161),
            .I(N__82158));
    LocalMux I__19667 (
            .O(N__82158),
            .I(N__82154));
    InMux I__19666 (
            .O(N__82157),
            .I(N__82151));
    Span4Mux_v I__19665 (
            .O(N__82154),
            .I(N__82146));
    LocalMux I__19664 (
            .O(N__82151),
            .I(N__82146));
    Span4Mux_h I__19663 (
            .O(N__82146),
            .I(N__82143));
    Span4Mux_h I__19662 (
            .O(N__82143),
            .I(N__82140));
    Odrv4 I__19661 (
            .O(N__82140),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ));
    InMux I__19660 (
            .O(N__82137),
            .I(N__82134));
    LocalMux I__19659 (
            .O(N__82134),
            .I(N__82131));
    Odrv4 I__19658 (
            .O(N__82131),
            .I(\pid_side.O_1_21 ));
    InMux I__19657 (
            .O(N__82128),
            .I(N__82123));
    InMux I__19656 (
            .O(N__82127),
            .I(N__82118));
    InMux I__19655 (
            .O(N__82126),
            .I(N__82118));
    LocalMux I__19654 (
            .O(N__82123),
            .I(\pid_side.error_d_regZ0Z_19 ));
    LocalMux I__19653 (
            .O(N__82118),
            .I(\pid_side.error_d_regZ0Z_19 ));
    InMux I__19652 (
            .O(N__82113),
            .I(N__82107));
    InMux I__19651 (
            .O(N__82112),
            .I(N__82107));
    LocalMux I__19650 (
            .O(N__82107),
            .I(N__82104));
    Odrv12 I__19649 (
            .O(N__82104),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ));
    InMux I__19648 (
            .O(N__82101),
            .I(N__82096));
    InMux I__19647 (
            .O(N__82100),
            .I(N__82091));
    InMux I__19646 (
            .O(N__82099),
            .I(N__82091));
    LocalMux I__19645 (
            .O(N__82096),
            .I(\pid_side.error_d_regZ0Z_11 ));
    LocalMux I__19644 (
            .O(N__82091),
            .I(\pid_side.error_d_regZ0Z_11 ));
    InMux I__19643 (
            .O(N__82086),
            .I(N__82079));
    InMux I__19642 (
            .O(N__82085),
            .I(N__82079));
    InMux I__19641 (
            .O(N__82084),
            .I(N__82076));
    LocalMux I__19640 (
            .O(N__82079),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    LocalMux I__19639 (
            .O(N__82076),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    CascadeMux I__19638 (
            .O(N__82071),
            .I(N__82066));
    InMux I__19637 (
            .O(N__82070),
            .I(N__82063));
    InMux I__19636 (
            .O(N__82069),
            .I(N__82060));
    InMux I__19635 (
            .O(N__82066),
            .I(N__82056));
    LocalMux I__19634 (
            .O(N__82063),
            .I(N__82051));
    LocalMux I__19633 (
            .O(N__82060),
            .I(N__82051));
    InMux I__19632 (
            .O(N__82059),
            .I(N__82048));
    LocalMux I__19631 (
            .O(N__82056),
            .I(N__82043));
    Span4Mux_v I__19630 (
            .O(N__82051),
            .I(N__82043));
    LocalMux I__19629 (
            .O(N__82048),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    Odrv4 I__19628 (
            .O(N__82043),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    InMux I__19627 (
            .O(N__82038),
            .I(N__82035));
    LocalMux I__19626 (
            .O(N__82035),
            .I(N__82032));
    Span4Mux_v I__19625 (
            .O(N__82032),
            .I(N__82029));
    Odrv4 I__19624 (
            .O(N__82029),
            .I(\pid_side.O_2_14 ));
    InMux I__19623 (
            .O(N__82026),
            .I(N__82019));
    InMux I__19622 (
            .O(N__82025),
            .I(N__82019));
    InMux I__19621 (
            .O(N__82024),
            .I(N__82016));
    LocalMux I__19620 (
            .O(N__82019),
            .I(\pid_side.error_p_regZ0Z_11 ));
    LocalMux I__19619 (
            .O(N__82016),
            .I(\pid_side.error_p_regZ0Z_11 ));
    InMux I__19618 (
            .O(N__82011),
            .I(N__82008));
    LocalMux I__19617 (
            .O(N__82008),
            .I(N__82005));
    Span4Mux_h I__19616 (
            .O(N__82005),
            .I(N__82001));
    InMux I__19615 (
            .O(N__82004),
            .I(N__81998));
    Span4Mux_h I__19614 (
            .O(N__82001),
            .I(N__81995));
    LocalMux I__19613 (
            .O(N__81998),
            .I(N__81992));
    Odrv4 I__19612 (
            .O(N__81995),
            .I(\pid_side.error_p_regZ0Z_20 ));
    Odrv12 I__19611 (
            .O(N__81992),
            .I(\pid_side.error_p_regZ0Z_20 ));
    InMux I__19610 (
            .O(N__81987),
            .I(N__81984));
    LocalMux I__19609 (
            .O(N__81984),
            .I(N__81981));
    Span4Mux_s2_h I__19608 (
            .O(N__81981),
            .I(N__81977));
    InMux I__19607 (
            .O(N__81980),
            .I(N__81974));
    Span4Mux_h I__19606 (
            .O(N__81977),
            .I(N__81971));
    LocalMux I__19605 (
            .O(N__81974),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    Odrv4 I__19604 (
            .O(N__81971),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    InMux I__19603 (
            .O(N__81966),
            .I(N__81963));
    LocalMux I__19602 (
            .O(N__81963),
            .I(N__81959));
    InMux I__19601 (
            .O(N__81962),
            .I(N__81956));
    Span4Mux_v I__19600 (
            .O(N__81959),
            .I(N__81951));
    LocalMux I__19599 (
            .O(N__81956),
            .I(N__81951));
    Span4Mux_h I__19598 (
            .O(N__81951),
            .I(N__81948));
    Span4Mux_h I__19597 (
            .O(N__81948),
            .I(N__81945));
    Odrv4 I__19596 (
            .O(N__81945),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ));
    InMux I__19595 (
            .O(N__81942),
            .I(N__81939));
    LocalMux I__19594 (
            .O(N__81939),
            .I(\pid_side.O_0_2 ));
    InMux I__19593 (
            .O(N__81936),
            .I(N__81930));
    InMux I__19592 (
            .O(N__81935),
            .I(N__81930));
    LocalMux I__19591 (
            .O(N__81930),
            .I(N__81924));
    InMux I__19590 (
            .O(N__81929),
            .I(N__81917));
    InMux I__19589 (
            .O(N__81928),
            .I(N__81917));
    InMux I__19588 (
            .O(N__81927),
            .I(N__81917));
    Span4Mux_h I__19587 (
            .O(N__81924),
            .I(N__81914));
    LocalMux I__19586 (
            .O(N__81917),
            .I(N__81911));
    Odrv4 I__19585 (
            .O(N__81914),
            .I(\pid_side.error_d_regZ0Z_0 ));
    Odrv12 I__19584 (
            .O(N__81911),
            .I(\pid_side.error_d_regZ0Z_0 ));
    InMux I__19583 (
            .O(N__81906),
            .I(N__81903));
    LocalMux I__19582 (
            .O(N__81903),
            .I(\pid_side.O_1_3 ));
    InMux I__19581 (
            .O(N__81900),
            .I(N__81895));
    InMux I__19580 (
            .O(N__81899),
            .I(N__81890));
    InMux I__19579 (
            .O(N__81898),
            .I(N__81890));
    LocalMux I__19578 (
            .O(N__81895),
            .I(N__81882));
    LocalMux I__19577 (
            .O(N__81890),
            .I(N__81882));
    InMux I__19576 (
            .O(N__81889),
            .I(N__81875));
    InMux I__19575 (
            .O(N__81888),
            .I(N__81875));
    InMux I__19574 (
            .O(N__81887),
            .I(N__81875));
    Span4Mux_h I__19573 (
            .O(N__81882),
            .I(N__81872));
    LocalMux I__19572 (
            .O(N__81875),
            .I(N__81869));
    Odrv4 I__19571 (
            .O(N__81872),
            .I(\pid_side.error_d_regZ0Z_1 ));
    Odrv12 I__19570 (
            .O(N__81869),
            .I(\pid_side.error_d_regZ0Z_1 ));
    InMux I__19569 (
            .O(N__81864),
            .I(N__81861));
    LocalMux I__19568 (
            .O(N__81861),
            .I(N__81858));
    Span4Mux_v I__19567 (
            .O(N__81858),
            .I(N__81855));
    Odrv4 I__19566 (
            .O(N__81855),
            .I(\pid_side.O_2_15 ));
    InMux I__19565 (
            .O(N__81852),
            .I(N__81848));
    InMux I__19564 (
            .O(N__81851),
            .I(N__81845));
    LocalMux I__19563 (
            .O(N__81848),
            .I(N__81842));
    LocalMux I__19562 (
            .O(N__81845),
            .I(N__81839));
    Span4Mux_h I__19561 (
            .O(N__81842),
            .I(N__81833));
    Span4Mux_h I__19560 (
            .O(N__81839),
            .I(N__81830));
    InMux I__19559 (
            .O(N__81838),
            .I(N__81823));
    InMux I__19558 (
            .O(N__81837),
            .I(N__81823));
    InMux I__19557 (
            .O(N__81836),
            .I(N__81823));
    Odrv4 I__19556 (
            .O(N__81833),
            .I(\pid_side.error_p_regZ0Z_12 ));
    Odrv4 I__19555 (
            .O(N__81830),
            .I(\pid_side.error_p_regZ0Z_12 ));
    LocalMux I__19554 (
            .O(N__81823),
            .I(\pid_side.error_p_regZ0Z_12 ));
    InMux I__19553 (
            .O(N__81816),
            .I(N__81813));
    LocalMux I__19552 (
            .O(N__81813),
            .I(\pid_side.O_2_13 ));
    CascadeMux I__19551 (
            .O(N__81810),
            .I(N__81805));
    CascadeMux I__19550 (
            .O(N__81809),
            .I(N__81802));
    InMux I__19549 (
            .O(N__81808),
            .I(N__81799));
    InMux I__19548 (
            .O(N__81805),
            .I(N__81794));
    InMux I__19547 (
            .O(N__81802),
            .I(N__81794));
    LocalMux I__19546 (
            .O(N__81799),
            .I(N__81791));
    LocalMux I__19545 (
            .O(N__81794),
            .I(N__81788));
    Span4Mux_v I__19544 (
            .O(N__81791),
            .I(N__81783));
    Span4Mux_v I__19543 (
            .O(N__81788),
            .I(N__81783));
    Odrv4 I__19542 (
            .O(N__81783),
            .I(\pid_side.error_p_regZ0Z_10 ));
    InMux I__19541 (
            .O(N__81780),
            .I(N__81777));
    LocalMux I__19540 (
            .O(N__81777),
            .I(\pid_side.O_2_9 ));
    CascadeMux I__19539 (
            .O(N__81774),
            .I(N__81770));
    InMux I__19538 (
            .O(N__81773),
            .I(N__81767));
    InMux I__19537 (
            .O(N__81770),
            .I(N__81764));
    LocalMux I__19536 (
            .O(N__81767),
            .I(N__81759));
    LocalMux I__19535 (
            .O(N__81764),
            .I(N__81759));
    Span4Mux_v I__19534 (
            .O(N__81759),
            .I(N__81756));
    Odrv4 I__19533 (
            .O(N__81756),
            .I(\pid_side.error_p_regZ0Z_6 ));
    InMux I__19532 (
            .O(N__81753),
            .I(N__81750));
    LocalMux I__19531 (
            .O(N__81750),
            .I(N__81747));
    Span4Mux_v I__19530 (
            .O(N__81747),
            .I(N__81744));
    Odrv4 I__19529 (
            .O(N__81744),
            .I(\pid_side.O_2_3 ));
    CascadeMux I__19528 (
            .O(N__81741),
            .I(N__81738));
    InMux I__19527 (
            .O(N__81738),
            .I(N__81735));
    LocalMux I__19526 (
            .O(N__81735),
            .I(N__81731));
    InMux I__19525 (
            .O(N__81734),
            .I(N__81728));
    Span4Mux_v I__19524 (
            .O(N__81731),
            .I(N__81723));
    LocalMux I__19523 (
            .O(N__81728),
            .I(N__81723));
    Span4Mux_h I__19522 (
            .O(N__81723),
            .I(N__81720));
    Odrv4 I__19521 (
            .O(N__81720),
            .I(\pid_side.error_p_regZ0Z_0 ));
    InMux I__19520 (
            .O(N__81717),
            .I(N__81714));
    LocalMux I__19519 (
            .O(N__81714),
            .I(N__81711));
    Span4Mux_h I__19518 (
            .O(N__81711),
            .I(N__81708));
    Odrv4 I__19517 (
            .O(N__81708),
            .I(\pid_side.O_1_19 ));
    InMux I__19516 (
            .O(N__81705),
            .I(N__81700));
    InMux I__19515 (
            .O(N__81704),
            .I(N__81697));
    InMux I__19514 (
            .O(N__81703),
            .I(N__81694));
    LocalMux I__19513 (
            .O(N__81700),
            .I(N__81691));
    LocalMux I__19512 (
            .O(N__81697),
            .I(N__81688));
    LocalMux I__19511 (
            .O(N__81694),
            .I(N__81683));
    Span4Mux_v I__19510 (
            .O(N__81691),
            .I(N__81683));
    Span4Mux_h I__19509 (
            .O(N__81688),
            .I(N__81680));
    Odrv4 I__19508 (
            .O(N__81683),
            .I(\pid_side.error_d_regZ0Z_17 ));
    Odrv4 I__19507 (
            .O(N__81680),
            .I(\pid_side.error_d_regZ0Z_17 ));
    InMux I__19506 (
            .O(N__81675),
            .I(N__81672));
    LocalMux I__19505 (
            .O(N__81672),
            .I(N__81669));
    Odrv4 I__19504 (
            .O(N__81669),
            .I(\pid_side.O_1_20 ));
    InMux I__19503 (
            .O(N__81666),
            .I(N__81657));
    InMux I__19502 (
            .O(N__81665),
            .I(N__81657));
    InMux I__19501 (
            .O(N__81664),
            .I(N__81657));
    LocalMux I__19500 (
            .O(N__81657),
            .I(\pid_side.error_d_regZ0Z_18 ));
    InMux I__19499 (
            .O(N__81654),
            .I(N__81651));
    LocalMux I__19498 (
            .O(N__81651),
            .I(N__81648));
    Odrv4 I__19497 (
            .O(N__81648),
            .I(\pid_side.O_1_18 ));
    InMux I__19496 (
            .O(N__81645),
            .I(N__81636));
    InMux I__19495 (
            .O(N__81644),
            .I(N__81636));
    InMux I__19494 (
            .O(N__81643),
            .I(N__81636));
    LocalMux I__19493 (
            .O(N__81636),
            .I(N__81633));
    Odrv4 I__19492 (
            .O(N__81633),
            .I(\pid_side.error_d_regZ0Z_16 ));
    InMux I__19491 (
            .O(N__81630),
            .I(N__81627));
    LocalMux I__19490 (
            .O(N__81627),
            .I(N__81624));
    Odrv4 I__19489 (
            .O(N__81624),
            .I(\pid_side.O_1_17 ));
    InMux I__19488 (
            .O(N__81621),
            .I(N__81612));
    InMux I__19487 (
            .O(N__81620),
            .I(N__81612));
    InMux I__19486 (
            .O(N__81619),
            .I(N__81612));
    LocalMux I__19485 (
            .O(N__81612),
            .I(N__81609));
    Odrv4 I__19484 (
            .O(N__81609),
            .I(\pid_side.error_d_regZ0Z_15 ));
    InMux I__19483 (
            .O(N__81606),
            .I(N__81603));
    LocalMux I__19482 (
            .O(N__81603),
            .I(N__81600));
    Span4Mux_h I__19481 (
            .O(N__81600),
            .I(N__81597));
    Odrv4 I__19480 (
            .O(N__81597),
            .I(\pid_side.O_1_24 ));
    CascadeMux I__19479 (
            .O(N__81594),
            .I(N__81588));
    InMux I__19478 (
            .O(N__81593),
            .I(N__81578));
    InMux I__19477 (
            .O(N__81592),
            .I(N__81578));
    InMux I__19476 (
            .O(N__81591),
            .I(N__81578));
    InMux I__19475 (
            .O(N__81588),
            .I(N__81575));
    InMux I__19474 (
            .O(N__81587),
            .I(N__81563));
    InMux I__19473 (
            .O(N__81586),
            .I(N__81563));
    InMux I__19472 (
            .O(N__81585),
            .I(N__81563));
    LocalMux I__19471 (
            .O(N__81578),
            .I(N__81558));
    LocalMux I__19470 (
            .O(N__81575),
            .I(N__81558));
    InMux I__19469 (
            .O(N__81574),
            .I(N__81553));
    InMux I__19468 (
            .O(N__81573),
            .I(N__81553));
    CascadeMux I__19467 (
            .O(N__81572),
            .I(N__81550));
    CascadeMux I__19466 (
            .O(N__81571),
            .I(N__81547));
    CascadeMux I__19465 (
            .O(N__81570),
            .I(N__81544));
    LocalMux I__19464 (
            .O(N__81563),
            .I(N__81539));
    Span4Mux_v I__19463 (
            .O(N__81558),
            .I(N__81534));
    LocalMux I__19462 (
            .O(N__81553),
            .I(N__81534));
    InMux I__19461 (
            .O(N__81550),
            .I(N__81523));
    InMux I__19460 (
            .O(N__81547),
            .I(N__81523));
    InMux I__19459 (
            .O(N__81544),
            .I(N__81523));
    InMux I__19458 (
            .O(N__81543),
            .I(N__81523));
    InMux I__19457 (
            .O(N__81542),
            .I(N__81523));
    Span4Mux_h I__19456 (
            .O(N__81539),
            .I(N__81520));
    Span4Mux_h I__19455 (
            .O(N__81534),
            .I(N__81517));
    LocalMux I__19454 (
            .O(N__81523),
            .I(N__81514));
    Span4Mux_h I__19453 (
            .O(N__81520),
            .I(N__81511));
    Span4Mux_h I__19452 (
            .O(N__81517),
            .I(N__81508));
    Span12Mux_h I__19451 (
            .O(N__81514),
            .I(N__81505));
    Odrv4 I__19450 (
            .O(N__81511),
            .I(\pid_side.error_d_regZ0Z_22 ));
    Odrv4 I__19449 (
            .O(N__81508),
            .I(\pid_side.error_d_regZ0Z_22 ));
    Odrv12 I__19448 (
            .O(N__81505),
            .I(\pid_side.error_d_regZ0Z_22 ));
    InMux I__19447 (
            .O(N__81498),
            .I(N__81495));
    LocalMux I__19446 (
            .O(N__81495),
            .I(N__81492));
    Odrv4 I__19445 (
            .O(N__81492),
            .I(\pid_side.O_2_19 ));
    InMux I__19444 (
            .O(N__81489),
            .I(N__81483));
    InMux I__19443 (
            .O(N__81488),
            .I(N__81483));
    LocalMux I__19442 (
            .O(N__81483),
            .I(N__81480));
    Span4Mux_v I__19441 (
            .O(N__81480),
            .I(N__81477));
    Odrv4 I__19440 (
            .O(N__81477),
            .I(\pid_side.error_p_regZ0Z_16 ));
    InMux I__19439 (
            .O(N__81474),
            .I(N__81471));
    LocalMux I__19438 (
            .O(N__81471),
            .I(N__81468));
    Odrv4 I__19437 (
            .O(N__81468),
            .I(\pid_side.O_2_18 ));
    InMux I__19436 (
            .O(N__81465),
            .I(N__81459));
    InMux I__19435 (
            .O(N__81464),
            .I(N__81459));
    LocalMux I__19434 (
            .O(N__81459),
            .I(N__81456));
    Span4Mux_v I__19433 (
            .O(N__81456),
            .I(N__81453));
    Odrv4 I__19432 (
            .O(N__81453),
            .I(\pid_side.error_p_regZ0Z_15 ));
    InMux I__19431 (
            .O(N__81450),
            .I(N__81447));
    LocalMux I__19430 (
            .O(N__81447),
            .I(N__81444));
    Odrv4 I__19429 (
            .O(N__81444),
            .I(\pid_side.O_2_23 ));
    InMux I__19428 (
            .O(N__81441),
            .I(N__81438));
    LocalMux I__19427 (
            .O(N__81438),
            .I(\pid_side.O_2_12 ));
    InMux I__19426 (
            .O(N__81435),
            .I(N__81429));
    InMux I__19425 (
            .O(N__81434),
            .I(N__81429));
    LocalMux I__19424 (
            .O(N__81429),
            .I(N__81426));
    Span12Mux_h I__19423 (
            .O(N__81426),
            .I(N__81423));
    Odrv12 I__19422 (
            .O(N__81423),
            .I(\pid_side.error_p_regZ0Z_9 ));
    InMux I__19421 (
            .O(N__81420),
            .I(N__81417));
    LocalMux I__19420 (
            .O(N__81417),
            .I(\pid_side.O_2_22 ));
    InMux I__19419 (
            .O(N__81414),
            .I(N__81411));
    LocalMux I__19418 (
            .O(N__81411),
            .I(\pid_side.O_2_20 ));
    InMux I__19417 (
            .O(N__81408),
            .I(N__81404));
    InMux I__19416 (
            .O(N__81407),
            .I(N__81401));
    LocalMux I__19415 (
            .O(N__81404),
            .I(N__81396));
    LocalMux I__19414 (
            .O(N__81401),
            .I(N__81396));
    Span4Mux_v I__19413 (
            .O(N__81396),
            .I(N__81393));
    Odrv4 I__19412 (
            .O(N__81393),
            .I(\pid_side.error_p_regZ0Z_17 ));
    InMux I__19411 (
            .O(N__81390),
            .I(N__81387));
    LocalMux I__19410 (
            .O(N__81387),
            .I(\pid_side.O_2_21 ));
    InMux I__19409 (
            .O(N__81384),
            .I(N__81378));
    InMux I__19408 (
            .O(N__81383),
            .I(N__81378));
    LocalMux I__19407 (
            .O(N__81378),
            .I(N__81375));
    Span4Mux_h I__19406 (
            .O(N__81375),
            .I(N__81372));
    Odrv4 I__19405 (
            .O(N__81372),
            .I(\pid_side.error_p_regZ0Z_18 ));
    InMux I__19404 (
            .O(N__81369),
            .I(N__81366));
    LocalMux I__19403 (
            .O(N__81366),
            .I(\pid_side.O_2_8 ));
    CascadeMux I__19402 (
            .O(N__81363),
            .I(N__81359));
    InMux I__19401 (
            .O(N__81362),
            .I(N__81354));
    InMux I__19400 (
            .O(N__81359),
            .I(N__81354));
    LocalMux I__19399 (
            .O(N__81354),
            .I(N__81351));
    Span4Mux_h I__19398 (
            .O(N__81351),
            .I(N__81348));
    Odrv4 I__19397 (
            .O(N__81348),
            .I(\pid_side.error_p_regZ0Z_5 ));
    InMux I__19396 (
            .O(N__81345),
            .I(N__81342));
    LocalMux I__19395 (
            .O(N__81342),
            .I(\pid_side.O_2_10 ));
    CascadeMux I__19394 (
            .O(N__81339),
            .I(N__81336));
    InMux I__19393 (
            .O(N__81336),
            .I(N__81330));
    InMux I__19392 (
            .O(N__81335),
            .I(N__81330));
    LocalMux I__19391 (
            .O(N__81330),
            .I(N__81327));
    Span4Mux_v I__19390 (
            .O(N__81327),
            .I(N__81324));
    Odrv4 I__19389 (
            .O(N__81324),
            .I(\pid_side.error_p_regZ0Z_7 ));
    InMux I__19388 (
            .O(N__81321),
            .I(N__81318));
    LocalMux I__19387 (
            .O(N__81318),
            .I(N__81315));
    Odrv4 I__19386 (
            .O(N__81315),
            .I(\pid_side.error_p_reg_esr_RNIVKIOZ0Z_12 ));
    InMux I__19385 (
            .O(N__81312),
            .I(N__81309));
    LocalMux I__19384 (
            .O(N__81309),
            .I(N__81305));
    InMux I__19383 (
            .O(N__81308),
            .I(N__81300));
    Span4Mux_h I__19382 (
            .O(N__81305),
            .I(N__81297));
    CascadeMux I__19381 (
            .O(N__81304),
            .I(N__81292));
    CascadeMux I__19380 (
            .O(N__81303),
            .I(N__81289));
    LocalMux I__19379 (
            .O(N__81300),
            .I(N__81285));
    Span4Mux_h I__19378 (
            .O(N__81297),
            .I(N__81282));
    InMux I__19377 (
            .O(N__81296),
            .I(N__81279));
    InMux I__19376 (
            .O(N__81295),
            .I(N__81276));
    InMux I__19375 (
            .O(N__81292),
            .I(N__81269));
    InMux I__19374 (
            .O(N__81289),
            .I(N__81269));
    InMux I__19373 (
            .O(N__81288),
            .I(N__81269));
    Odrv4 I__19372 (
            .O(N__81285),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__19371 (
            .O(N__81282),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19370 (
            .O(N__81279),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19369 (
            .O(N__81276),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19368 (
            .O(N__81269),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    CEMux I__19367 (
            .O(N__81258),
            .I(N__81253));
    CEMux I__19366 (
            .O(N__81257),
            .I(N__81250));
    CEMux I__19365 (
            .O(N__81256),
            .I(N__81244));
    LocalMux I__19364 (
            .O(N__81253),
            .I(N__81240));
    LocalMux I__19363 (
            .O(N__81250),
            .I(N__81237));
    CEMux I__19362 (
            .O(N__81249),
            .I(N__81234));
    CEMux I__19361 (
            .O(N__81248),
            .I(N__81231));
    CEMux I__19360 (
            .O(N__81247),
            .I(N__81227));
    LocalMux I__19359 (
            .O(N__81244),
            .I(N__81224));
    CEMux I__19358 (
            .O(N__81243),
            .I(N__81221));
    Span4Mux_v I__19357 (
            .O(N__81240),
            .I(N__81216));
    Span4Mux_v I__19356 (
            .O(N__81237),
            .I(N__81216));
    LocalMux I__19355 (
            .O(N__81234),
            .I(N__81211));
    LocalMux I__19354 (
            .O(N__81231),
            .I(N__81211));
    CEMux I__19353 (
            .O(N__81230),
            .I(N__81208));
    LocalMux I__19352 (
            .O(N__81227),
            .I(N__81205));
    Span4Mux_v I__19351 (
            .O(N__81224),
            .I(N__81200));
    LocalMux I__19350 (
            .O(N__81221),
            .I(N__81200));
    Span4Mux_h I__19349 (
            .O(N__81216),
            .I(N__81192));
    Span4Mux_v I__19348 (
            .O(N__81211),
            .I(N__81192));
    LocalMux I__19347 (
            .O(N__81208),
            .I(N__81192));
    Span4Mux_v I__19346 (
            .O(N__81205),
            .I(N__81186));
    Span4Mux_v I__19345 (
            .O(N__81200),
            .I(N__81183));
    CEMux I__19344 (
            .O(N__81199),
            .I(N__81180));
    Span4Mux_h I__19343 (
            .O(N__81192),
            .I(N__81177));
    CEMux I__19342 (
            .O(N__81191),
            .I(N__81174));
    CEMux I__19341 (
            .O(N__81190),
            .I(N__81171));
    CEMux I__19340 (
            .O(N__81189),
            .I(N__81168));
    Odrv4 I__19339 (
            .O(N__81186),
            .I(\pid_side.N_478_0 ));
    Odrv4 I__19338 (
            .O(N__81183),
            .I(\pid_side.N_478_0 ));
    LocalMux I__19337 (
            .O(N__81180),
            .I(\pid_side.N_478_0 ));
    Odrv4 I__19336 (
            .O(N__81177),
            .I(\pid_side.N_478_0 ));
    LocalMux I__19335 (
            .O(N__81174),
            .I(\pid_side.N_478_0 ));
    LocalMux I__19334 (
            .O(N__81171),
            .I(\pid_side.N_478_0 ));
    LocalMux I__19333 (
            .O(N__81168),
            .I(\pid_side.N_478_0 ));
    InMux I__19332 (
            .O(N__81153),
            .I(N__81150));
    LocalMux I__19331 (
            .O(N__81150),
            .I(N__81135));
    SRMux I__19330 (
            .O(N__81149),
            .I(N__81108));
    SRMux I__19329 (
            .O(N__81148),
            .I(N__81108));
    SRMux I__19328 (
            .O(N__81147),
            .I(N__81108));
    SRMux I__19327 (
            .O(N__81146),
            .I(N__81108));
    SRMux I__19326 (
            .O(N__81145),
            .I(N__81108));
    SRMux I__19325 (
            .O(N__81144),
            .I(N__81108));
    SRMux I__19324 (
            .O(N__81143),
            .I(N__81108));
    SRMux I__19323 (
            .O(N__81142),
            .I(N__81108));
    SRMux I__19322 (
            .O(N__81141),
            .I(N__81108));
    SRMux I__19321 (
            .O(N__81140),
            .I(N__81108));
    SRMux I__19320 (
            .O(N__81139),
            .I(N__81108));
    SRMux I__19319 (
            .O(N__81138),
            .I(N__81108));
    Glb2LocalMux I__19318 (
            .O(N__81135),
            .I(N__81108));
    GlobalMux I__19317 (
            .O(N__81108),
            .I(N__81105));
    gio2CtrlBuf I__19316 (
            .O(N__81105),
            .I(\pid_side.N_1352_g ));
    InMux I__19315 (
            .O(N__81102),
            .I(N__81097));
    InMux I__19314 (
            .O(N__81101),
            .I(N__81094));
    InMux I__19313 (
            .O(N__81100),
            .I(N__81090));
    LocalMux I__19312 (
            .O(N__81097),
            .I(N__81087));
    LocalMux I__19311 (
            .O(N__81094),
            .I(N__81082));
    InMux I__19310 (
            .O(N__81093),
            .I(N__81077));
    LocalMux I__19309 (
            .O(N__81090),
            .I(N__81072));
    Span4Mux_v I__19308 (
            .O(N__81087),
            .I(N__81069));
    InMux I__19307 (
            .O(N__81086),
            .I(N__81066));
    InMux I__19306 (
            .O(N__81085),
            .I(N__81063));
    Span4Mux_v I__19305 (
            .O(N__81082),
            .I(N__81060));
    InMux I__19304 (
            .O(N__81081),
            .I(N__81056));
    InMux I__19303 (
            .O(N__81080),
            .I(N__81053));
    LocalMux I__19302 (
            .O(N__81077),
            .I(N__81050));
    InMux I__19301 (
            .O(N__81076),
            .I(N__81047));
    InMux I__19300 (
            .O(N__81075),
            .I(N__81044));
    Span4Mux_h I__19299 (
            .O(N__81072),
            .I(N__81041));
    Sp12to4 I__19298 (
            .O(N__81069),
            .I(N__81038));
    LocalMux I__19297 (
            .O(N__81066),
            .I(N__81035));
    LocalMux I__19296 (
            .O(N__81063),
            .I(N__81032));
    Span4Mux_h I__19295 (
            .O(N__81060),
            .I(N__81029));
    InMux I__19294 (
            .O(N__81059),
            .I(N__81026));
    LocalMux I__19293 (
            .O(N__81056),
            .I(N__81023));
    LocalMux I__19292 (
            .O(N__81053),
            .I(N__81020));
    Span4Mux_v I__19291 (
            .O(N__81050),
            .I(N__81017));
    LocalMux I__19290 (
            .O(N__81047),
            .I(N__81014));
    LocalMux I__19289 (
            .O(N__81044),
            .I(N__81011));
    Sp12to4 I__19288 (
            .O(N__81041),
            .I(N__81007));
    Span12Mux_h I__19287 (
            .O(N__81038),
            .I(N__81000));
    Sp12to4 I__19286 (
            .O(N__81035),
            .I(N__81000));
    Span12Mux_s8_h I__19285 (
            .O(N__81032),
            .I(N__81000));
    Span4Mux_v I__19284 (
            .O(N__81029),
            .I(N__80997));
    LocalMux I__19283 (
            .O(N__81026),
            .I(N__80992));
    Span4Mux_h I__19282 (
            .O(N__81023),
            .I(N__80992));
    Span4Mux_v I__19281 (
            .O(N__81020),
            .I(N__80989));
    Span4Mux_h I__19280 (
            .O(N__81017),
            .I(N__80986));
    Span4Mux_h I__19279 (
            .O(N__81014),
            .I(N__80983));
    Span4Mux_h I__19278 (
            .O(N__81011),
            .I(N__80979));
    InMux I__19277 (
            .O(N__81010),
            .I(N__80976));
    Span12Mux_v I__19276 (
            .O(N__81007),
            .I(N__80971));
    Span12Mux_v I__19275 (
            .O(N__81000),
            .I(N__80971));
    Span4Mux_v I__19274 (
            .O(N__80997),
            .I(N__80964));
    Span4Mux_v I__19273 (
            .O(N__80992),
            .I(N__80964));
    Span4Mux_h I__19272 (
            .O(N__80989),
            .I(N__80964));
    Span4Mux_h I__19271 (
            .O(N__80986),
            .I(N__80959));
    Span4Mux_h I__19270 (
            .O(N__80983),
            .I(N__80959));
    InMux I__19269 (
            .O(N__80982),
            .I(N__80956));
    Odrv4 I__19268 (
            .O(N__80979),
            .I(uart_pc_data_6));
    LocalMux I__19267 (
            .O(N__80976),
            .I(uart_pc_data_6));
    Odrv12 I__19266 (
            .O(N__80971),
            .I(uart_pc_data_6));
    Odrv4 I__19265 (
            .O(N__80964),
            .I(uart_pc_data_6));
    Odrv4 I__19264 (
            .O(N__80959),
            .I(uart_pc_data_6));
    LocalMux I__19263 (
            .O(N__80956),
            .I(uart_pc_data_6));
    InMux I__19262 (
            .O(N__80943),
            .I(N__80940));
    LocalMux I__19261 (
            .O(N__80940),
            .I(N__80936));
    InMux I__19260 (
            .O(N__80939),
            .I(N__80933));
    Span4Mux_s1_h I__19259 (
            .O(N__80936),
            .I(N__80930));
    LocalMux I__19258 (
            .O(N__80933),
            .I(N__80927));
    Span4Mux_v I__19257 (
            .O(N__80930),
            .I(N__80922));
    Span4Mux_s1_h I__19256 (
            .O(N__80927),
            .I(N__80922));
    Odrv4 I__19255 (
            .O(N__80922),
            .I(xy_kd_6));
    CEMux I__19254 (
            .O(N__80919),
            .I(N__80915));
    CEMux I__19253 (
            .O(N__80918),
            .I(N__80909));
    LocalMux I__19252 (
            .O(N__80915),
            .I(N__80906));
    CEMux I__19251 (
            .O(N__80914),
            .I(N__80903));
    CEMux I__19250 (
            .O(N__80913),
            .I(N__80900));
    CEMux I__19249 (
            .O(N__80912),
            .I(N__80897));
    LocalMux I__19248 (
            .O(N__80909),
            .I(N__80894));
    Span4Mux_v I__19247 (
            .O(N__80906),
            .I(N__80891));
    LocalMux I__19246 (
            .O(N__80903),
            .I(N__80886));
    LocalMux I__19245 (
            .O(N__80900),
            .I(N__80886));
    LocalMux I__19244 (
            .O(N__80897),
            .I(N__80883));
    Span4Mux_h I__19243 (
            .O(N__80894),
            .I(N__80878));
    Span4Mux_h I__19242 (
            .O(N__80891),
            .I(N__80878));
    Span4Mux_v I__19241 (
            .O(N__80886),
            .I(N__80875));
    Span4Mux_h I__19240 (
            .O(N__80883),
            .I(N__80872));
    Sp12to4 I__19239 (
            .O(N__80878),
            .I(N__80869));
    Sp12to4 I__19238 (
            .O(N__80875),
            .I(N__80866));
    Span4Mux_h I__19237 (
            .O(N__80872),
            .I(N__80863));
    Span12Mux_v I__19236 (
            .O(N__80869),
            .I(N__80858));
    Span12Mux_s6_h I__19235 (
            .O(N__80866),
            .I(N__80858));
    Span4Mux_v I__19234 (
            .O(N__80863),
            .I(N__80855));
    Span12Mux_h I__19233 (
            .O(N__80858),
            .I(N__80852));
    Span4Mux_h I__19232 (
            .O(N__80855),
            .I(N__80849));
    Odrv12 I__19231 (
            .O(N__80852),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    Odrv4 I__19230 (
            .O(N__80849),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    InMux I__19229 (
            .O(N__80844),
            .I(N__80841));
    LocalMux I__19228 (
            .O(N__80841),
            .I(N__80838));
    Odrv4 I__19227 (
            .O(N__80838),
            .I(\pid_side.O_2_24 ));
    InMux I__19226 (
            .O(N__80835),
            .I(N__80827));
    InMux I__19225 (
            .O(N__80834),
            .I(N__80822));
    InMux I__19224 (
            .O(N__80833),
            .I(N__80822));
    InMux I__19223 (
            .O(N__80832),
            .I(N__80815));
    InMux I__19222 (
            .O(N__80831),
            .I(N__80815));
    InMux I__19221 (
            .O(N__80830),
            .I(N__80815));
    LocalMux I__19220 (
            .O(N__80827),
            .I(N__80799));
    LocalMux I__19219 (
            .O(N__80822),
            .I(N__80799));
    LocalMux I__19218 (
            .O(N__80815),
            .I(N__80799));
    InMux I__19217 (
            .O(N__80814),
            .I(N__80788));
    InMux I__19216 (
            .O(N__80813),
            .I(N__80788));
    InMux I__19215 (
            .O(N__80812),
            .I(N__80788));
    InMux I__19214 (
            .O(N__80811),
            .I(N__80788));
    InMux I__19213 (
            .O(N__80810),
            .I(N__80788));
    InMux I__19212 (
            .O(N__80809),
            .I(N__80779));
    InMux I__19211 (
            .O(N__80808),
            .I(N__80779));
    InMux I__19210 (
            .O(N__80807),
            .I(N__80779));
    InMux I__19209 (
            .O(N__80806),
            .I(N__80779));
    Span4Mux_v I__19208 (
            .O(N__80799),
            .I(N__80774));
    LocalMux I__19207 (
            .O(N__80788),
            .I(N__80774));
    LocalMux I__19206 (
            .O(N__80779),
            .I(N__80771));
    Span4Mux_v I__19205 (
            .O(N__80774),
            .I(N__80768));
    Span4Mux_v I__19204 (
            .O(N__80771),
            .I(N__80765));
    Sp12to4 I__19203 (
            .O(N__80768),
            .I(N__80762));
    Span4Mux_v I__19202 (
            .O(N__80765),
            .I(N__80759));
    Span12Mux_h I__19201 (
            .O(N__80762),
            .I(N__80756));
    Span4Mux_h I__19200 (
            .O(N__80759),
            .I(N__80753));
    Odrv12 I__19199 (
            .O(N__80756),
            .I(\pid_side.error_p_regZ0Z_21 ));
    Odrv4 I__19198 (
            .O(N__80753),
            .I(\pid_side.error_p_regZ0Z_21 ));
    InMux I__19197 (
            .O(N__80748),
            .I(N__80745));
    LocalMux I__19196 (
            .O(N__80745),
            .I(N__80742));
    Odrv4 I__19195 (
            .O(N__80742),
            .I(\pid_side.O_2_16 ));
    InMux I__19194 (
            .O(N__80739),
            .I(N__80734));
    InMux I__19193 (
            .O(N__80738),
            .I(N__80729));
    InMux I__19192 (
            .O(N__80737),
            .I(N__80729));
    LocalMux I__19191 (
            .O(N__80734),
            .I(N__80726));
    LocalMux I__19190 (
            .O(N__80729),
            .I(N__80723));
    Span4Mux_h I__19189 (
            .O(N__80726),
            .I(N__80720));
    Span4Mux_h I__19188 (
            .O(N__80723),
            .I(N__80717));
    Span4Mux_v I__19187 (
            .O(N__80720),
            .I(N__80714));
    Span4Mux_v I__19186 (
            .O(N__80717),
            .I(N__80711));
    Odrv4 I__19185 (
            .O(N__80714),
            .I(\pid_side.error_p_regZ0Z_13 ));
    Odrv4 I__19184 (
            .O(N__80711),
            .I(\pid_side.error_p_regZ0Z_13 ));
    InMux I__19183 (
            .O(N__80706),
            .I(N__80703));
    LocalMux I__19182 (
            .O(N__80703),
            .I(N__80700));
    Odrv4 I__19181 (
            .O(N__80700),
            .I(\pid_side.O_2_17 ));
    InMux I__19180 (
            .O(N__80697),
            .I(N__80693));
    InMux I__19179 (
            .O(N__80696),
            .I(N__80690));
    LocalMux I__19178 (
            .O(N__80693),
            .I(N__80687));
    LocalMux I__19177 (
            .O(N__80690),
            .I(N__80682));
    Span4Mux_v I__19176 (
            .O(N__80687),
            .I(N__80682));
    Span4Mux_v I__19175 (
            .O(N__80682),
            .I(N__80679));
    Odrv4 I__19174 (
            .O(N__80679),
            .I(\pid_side.error_p_regZ0Z_14 ));
    InMux I__19173 (
            .O(N__80676),
            .I(N__80673));
    LocalMux I__19172 (
            .O(N__80673),
            .I(\pid_side.O_2_11 ));
    InMux I__19171 (
            .O(N__80670),
            .I(N__80664));
    InMux I__19170 (
            .O(N__80669),
            .I(N__80664));
    LocalMux I__19169 (
            .O(N__80664),
            .I(N__80661));
    Span4Mux_h I__19168 (
            .O(N__80661),
            .I(N__80658));
    Span4Mux_v I__19167 (
            .O(N__80658),
            .I(N__80655));
    Odrv4 I__19166 (
            .O(N__80655),
            .I(\pid_side.error_p_regZ0Z_8 ));
    InMux I__19165 (
            .O(N__80652),
            .I(N__80646));
    InMux I__19164 (
            .O(N__80651),
            .I(N__80646));
    LocalMux I__19163 (
            .O(N__80646),
            .I(\pid_side.error_d_reg_prevZ0Z_18 ));
    InMux I__19162 (
            .O(N__80643),
            .I(N__80640));
    LocalMux I__19161 (
            .O(N__80640),
            .I(N__80637));
    Span4Mux_h I__19160 (
            .O(N__80637),
            .I(N__80633));
    InMux I__19159 (
            .O(N__80636),
            .I(N__80630));
    Span4Mux_h I__19158 (
            .O(N__80633),
            .I(N__80627));
    LocalMux I__19157 (
            .O(N__80630),
            .I(N__80624));
    Odrv4 I__19156 (
            .O(N__80627),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ));
    Odrv12 I__19155 (
            .O(N__80624),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ));
    InMux I__19154 (
            .O(N__80619),
            .I(N__80616));
    LocalMux I__19153 (
            .O(N__80616),
            .I(N__80612));
    InMux I__19152 (
            .O(N__80615),
            .I(N__80609));
    Span4Mux_v I__19151 (
            .O(N__80612),
            .I(N__80604));
    LocalMux I__19150 (
            .O(N__80609),
            .I(N__80604));
    Span4Mux_h I__19149 (
            .O(N__80604),
            .I(N__80601));
    Odrv4 I__19148 (
            .O(N__80601),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ));
    InMux I__19147 (
            .O(N__80598),
            .I(N__80595));
    LocalMux I__19146 (
            .O(N__80595),
            .I(N__80592));
    Span4Mux_v I__19145 (
            .O(N__80592),
            .I(N__80589));
    Odrv4 I__19144 (
            .O(N__80589),
            .I(\pid_side.O_1_13 ));
    InMux I__19143 (
            .O(N__80586),
            .I(N__80582));
    InMux I__19142 (
            .O(N__80585),
            .I(N__80579));
    LocalMux I__19141 (
            .O(N__80582),
            .I(\pid_side.N_1905_i ));
    LocalMux I__19140 (
            .O(N__80579),
            .I(\pid_side.N_1905_i ));
    CascadeMux I__19139 (
            .O(N__80574),
            .I(\pid_side.N_1905_i_cascade_ ));
    CascadeMux I__19138 (
            .O(N__80571),
            .I(N__80568));
    InMux I__19137 (
            .O(N__80568),
            .I(N__80562));
    InMux I__19136 (
            .O(N__80567),
            .I(N__80562));
    LocalMux I__19135 (
            .O(N__80562),
            .I(N__80559));
    Span4Mux_h I__19134 (
            .O(N__80559),
            .I(N__80556));
    Span4Mux_h I__19133 (
            .O(N__80556),
            .I(N__80553));
    Odrv4 I__19132 (
            .O(N__80553),
            .I(\pid_side.error_p_reg_esr_RNIR3TQ1_0Z0Z_12 ));
    CascadeMux I__19131 (
            .O(N__80550),
            .I(N__80547));
    InMux I__19130 (
            .O(N__80547),
            .I(N__80542));
    InMux I__19129 (
            .O(N__80546),
            .I(N__80539));
    InMux I__19128 (
            .O(N__80545),
            .I(N__80536));
    LocalMux I__19127 (
            .O(N__80542),
            .I(\pid_side.un1_pid_prereg_79 ));
    LocalMux I__19126 (
            .O(N__80539),
            .I(\pid_side.un1_pid_prereg_79 ));
    LocalMux I__19125 (
            .O(N__80536),
            .I(\pid_side.un1_pid_prereg_79 ));
    CascadeMux I__19124 (
            .O(N__80529),
            .I(\pid_side.un1_pid_prereg_79_cascade_ ));
    InMux I__19123 (
            .O(N__80526),
            .I(N__80523));
    LocalMux I__19122 (
            .O(N__80523),
            .I(N__80520));
    Odrv4 I__19121 (
            .O(N__80520),
            .I(\pid_side.error_p_reg_esr_RNIVHA21Z0Z_12 ));
    InMux I__19120 (
            .O(N__80517),
            .I(N__80511));
    InMux I__19119 (
            .O(N__80516),
            .I(N__80506));
    InMux I__19118 (
            .O(N__80515),
            .I(N__80501));
    InMux I__19117 (
            .O(N__80514),
            .I(N__80497));
    LocalMux I__19116 (
            .O(N__80511),
            .I(N__80494));
    InMux I__19115 (
            .O(N__80510),
            .I(N__80488));
    InMux I__19114 (
            .O(N__80509),
            .I(N__80488));
    LocalMux I__19113 (
            .O(N__80506),
            .I(N__80485));
    InMux I__19112 (
            .O(N__80505),
            .I(N__80482));
    InMux I__19111 (
            .O(N__80504),
            .I(N__80478));
    LocalMux I__19110 (
            .O(N__80501),
            .I(N__80475));
    InMux I__19109 (
            .O(N__80500),
            .I(N__80472));
    LocalMux I__19108 (
            .O(N__80497),
            .I(N__80468));
    Span4Mux_v I__19107 (
            .O(N__80494),
            .I(N__80464));
    InMux I__19106 (
            .O(N__80493),
            .I(N__80460));
    LocalMux I__19105 (
            .O(N__80488),
            .I(N__80457));
    Span4Mux_v I__19104 (
            .O(N__80485),
            .I(N__80454));
    LocalMux I__19103 (
            .O(N__80482),
            .I(N__80451));
    InMux I__19102 (
            .O(N__80481),
            .I(N__80448));
    LocalMux I__19101 (
            .O(N__80478),
            .I(N__80445));
    Span4Mux_v I__19100 (
            .O(N__80475),
            .I(N__80440));
    LocalMux I__19099 (
            .O(N__80472),
            .I(N__80440));
    InMux I__19098 (
            .O(N__80471),
            .I(N__80437));
    Span4Mux_v I__19097 (
            .O(N__80468),
            .I(N__80434));
    InMux I__19096 (
            .O(N__80467),
            .I(N__80429));
    Span4Mux_h I__19095 (
            .O(N__80464),
            .I(N__80426));
    InMux I__19094 (
            .O(N__80463),
            .I(N__80423));
    LocalMux I__19093 (
            .O(N__80460),
            .I(N__80420));
    Sp12to4 I__19092 (
            .O(N__80457),
            .I(N__80417));
    Sp12to4 I__19091 (
            .O(N__80454),
            .I(N__80414));
    Span4Mux_h I__19090 (
            .O(N__80451),
            .I(N__80409));
    LocalMux I__19089 (
            .O(N__80448),
            .I(N__80404));
    Span4Mux_h I__19088 (
            .O(N__80445),
            .I(N__80404));
    Span4Mux_h I__19087 (
            .O(N__80440),
            .I(N__80401));
    LocalMux I__19086 (
            .O(N__80437),
            .I(N__80396));
    Sp12to4 I__19085 (
            .O(N__80434),
            .I(N__80396));
    InMux I__19084 (
            .O(N__80433),
            .I(N__80390));
    InMux I__19083 (
            .O(N__80432),
            .I(N__80390));
    LocalMux I__19082 (
            .O(N__80429),
            .I(N__80381));
    Sp12to4 I__19081 (
            .O(N__80426),
            .I(N__80381));
    LocalMux I__19080 (
            .O(N__80423),
            .I(N__80381));
    Span12Mux_h I__19079 (
            .O(N__80420),
            .I(N__80381));
    Span12Mux_v I__19078 (
            .O(N__80417),
            .I(N__80376));
    Span12Mux_s6_h I__19077 (
            .O(N__80414),
            .I(N__80376));
    InMux I__19076 (
            .O(N__80413),
            .I(N__80373));
    InMux I__19075 (
            .O(N__80412),
            .I(N__80370));
    Span4Mux_h I__19074 (
            .O(N__80409),
            .I(N__80367));
    Span4Mux_v I__19073 (
            .O(N__80404),
            .I(N__80362));
    Span4Mux_v I__19072 (
            .O(N__80401),
            .I(N__80362));
    Span12Mux_v I__19071 (
            .O(N__80396),
            .I(N__80359));
    InMux I__19070 (
            .O(N__80395),
            .I(N__80356));
    LocalMux I__19069 (
            .O(N__80390),
            .I(N__80347));
    Span12Mux_v I__19068 (
            .O(N__80381),
            .I(N__80347));
    Span12Mux_h I__19067 (
            .O(N__80376),
            .I(N__80347));
    LocalMux I__19066 (
            .O(N__80373),
            .I(N__80347));
    LocalMux I__19065 (
            .O(N__80370),
            .I(uart_pc_data_0));
    Odrv4 I__19064 (
            .O(N__80367),
            .I(uart_pc_data_0));
    Odrv4 I__19063 (
            .O(N__80362),
            .I(uart_pc_data_0));
    Odrv12 I__19062 (
            .O(N__80359),
            .I(uart_pc_data_0));
    LocalMux I__19061 (
            .O(N__80356),
            .I(uart_pc_data_0));
    Odrv12 I__19060 (
            .O(N__80347),
            .I(uart_pc_data_0));
    InMux I__19059 (
            .O(N__80334),
            .I(N__80331));
    LocalMux I__19058 (
            .O(N__80331),
            .I(N__80327));
    InMux I__19057 (
            .O(N__80330),
            .I(N__80324));
    Span4Mux_s2_h I__19056 (
            .O(N__80327),
            .I(N__80321));
    LocalMux I__19055 (
            .O(N__80324),
            .I(N__80318));
    Span4Mux_v I__19054 (
            .O(N__80321),
            .I(N__80313));
    Span4Mux_s2_h I__19053 (
            .O(N__80318),
            .I(N__80313));
    Odrv4 I__19052 (
            .O(N__80313),
            .I(xy_kd_0));
    InMux I__19051 (
            .O(N__80310),
            .I(N__80298));
    InMux I__19050 (
            .O(N__80309),
            .I(N__80298));
    InMux I__19049 (
            .O(N__80308),
            .I(N__80298));
    InMux I__19048 (
            .O(N__80307),
            .I(N__80298));
    LocalMux I__19047 (
            .O(N__80298),
            .I(N__80292));
    InMux I__19046 (
            .O(N__80297),
            .I(N__80288));
    InMux I__19045 (
            .O(N__80296),
            .I(N__80285));
    InMux I__19044 (
            .O(N__80295),
            .I(N__80282));
    Span4Mux_v I__19043 (
            .O(N__80292),
            .I(N__80279));
    InMux I__19042 (
            .O(N__80291),
            .I(N__80276));
    LocalMux I__19041 (
            .O(N__80288),
            .I(N__80272));
    LocalMux I__19040 (
            .O(N__80285),
            .I(N__80269));
    LocalMux I__19039 (
            .O(N__80282),
            .I(N__80266));
    Span4Mux_h I__19038 (
            .O(N__80279),
            .I(N__80263));
    LocalMux I__19037 (
            .O(N__80276),
            .I(N__80259));
    InMux I__19036 (
            .O(N__80275),
            .I(N__80255));
    Span4Mux_v I__19035 (
            .O(N__80272),
            .I(N__80250));
    Span4Mux_v I__19034 (
            .O(N__80269),
            .I(N__80250));
    Span4Mux_v I__19033 (
            .O(N__80266),
            .I(N__80245));
    Span4Mux_h I__19032 (
            .O(N__80263),
            .I(N__80242));
    InMux I__19031 (
            .O(N__80262),
            .I(N__80239));
    Span4Mux_h I__19030 (
            .O(N__80259),
            .I(N__80235));
    InMux I__19029 (
            .O(N__80258),
            .I(N__80232));
    LocalMux I__19028 (
            .O(N__80255),
            .I(N__80229));
    Sp12to4 I__19027 (
            .O(N__80250),
            .I(N__80226));
    InMux I__19026 (
            .O(N__80249),
            .I(N__80223));
    InMux I__19025 (
            .O(N__80248),
            .I(N__80220));
    Span4Mux_v I__19024 (
            .O(N__80245),
            .I(N__80217));
    Sp12to4 I__19023 (
            .O(N__80242),
            .I(N__80212));
    LocalMux I__19022 (
            .O(N__80239),
            .I(N__80212));
    InMux I__19021 (
            .O(N__80238),
            .I(N__80209));
    Sp12to4 I__19020 (
            .O(N__80235),
            .I(N__80206));
    LocalMux I__19019 (
            .O(N__80232),
            .I(N__80200));
    Span4Mux_s3_h I__19018 (
            .O(N__80229),
            .I(N__80196));
    Span12Mux_h I__19017 (
            .O(N__80226),
            .I(N__80191));
    LocalMux I__19016 (
            .O(N__80223),
            .I(N__80191));
    LocalMux I__19015 (
            .O(N__80220),
            .I(N__80188));
    Sp12to4 I__19014 (
            .O(N__80217),
            .I(N__80178));
    Span12Mux_v I__19013 (
            .O(N__80212),
            .I(N__80178));
    LocalMux I__19012 (
            .O(N__80209),
            .I(N__80178));
    Span12Mux_v I__19011 (
            .O(N__80206),
            .I(N__80178));
    InMux I__19010 (
            .O(N__80205),
            .I(N__80173));
    InMux I__19009 (
            .O(N__80204),
            .I(N__80173));
    InMux I__19008 (
            .O(N__80203),
            .I(N__80170));
    Span4Mux_h I__19007 (
            .O(N__80200),
            .I(N__80167));
    InMux I__19006 (
            .O(N__80199),
            .I(N__80164));
    Span4Mux_h I__19005 (
            .O(N__80196),
            .I(N__80161));
    Span12Mux_v I__19004 (
            .O(N__80191),
            .I(N__80156));
    Span12Mux_s8_v I__19003 (
            .O(N__80188),
            .I(N__80156));
    InMux I__19002 (
            .O(N__80187),
            .I(N__80153));
    Span12Mux_h I__19001 (
            .O(N__80178),
            .I(N__80146));
    LocalMux I__19000 (
            .O(N__80173),
            .I(N__80146));
    LocalMux I__18999 (
            .O(N__80170),
            .I(N__80146));
    Odrv4 I__18998 (
            .O(N__80167),
            .I(uart_pc_data_2));
    LocalMux I__18997 (
            .O(N__80164),
            .I(uart_pc_data_2));
    Odrv4 I__18996 (
            .O(N__80161),
            .I(uart_pc_data_2));
    Odrv12 I__18995 (
            .O(N__80156),
            .I(uart_pc_data_2));
    LocalMux I__18994 (
            .O(N__80153),
            .I(uart_pc_data_2));
    Odrv12 I__18993 (
            .O(N__80146),
            .I(uart_pc_data_2));
    InMux I__18992 (
            .O(N__80133),
            .I(N__80130));
    LocalMux I__18991 (
            .O(N__80130),
            .I(N__80126));
    InMux I__18990 (
            .O(N__80129),
            .I(N__80123));
    Span4Mux_s2_h I__18989 (
            .O(N__80126),
            .I(N__80120));
    LocalMux I__18988 (
            .O(N__80123),
            .I(N__80117));
    Span4Mux_v I__18987 (
            .O(N__80120),
            .I(N__80112));
    Span4Mux_s2_h I__18986 (
            .O(N__80117),
            .I(N__80112));
    Odrv4 I__18985 (
            .O(N__80112),
            .I(xy_kd_2));
    InMux I__18984 (
            .O(N__80109),
            .I(N__80101));
    InMux I__18983 (
            .O(N__80108),
            .I(N__80096));
    InMux I__18982 (
            .O(N__80107),
            .I(N__80093));
    InMux I__18981 (
            .O(N__80106),
            .I(N__80090));
    InMux I__18980 (
            .O(N__80105),
            .I(N__80085));
    InMux I__18979 (
            .O(N__80104),
            .I(N__80082));
    LocalMux I__18978 (
            .O(N__80101),
            .I(N__80078));
    InMux I__18977 (
            .O(N__80100),
            .I(N__80075));
    InMux I__18976 (
            .O(N__80099),
            .I(N__80071));
    LocalMux I__18975 (
            .O(N__80096),
            .I(N__80068));
    LocalMux I__18974 (
            .O(N__80093),
            .I(N__80063));
    LocalMux I__18973 (
            .O(N__80090),
            .I(N__80063));
    InMux I__18972 (
            .O(N__80089),
            .I(N__80060));
    InMux I__18971 (
            .O(N__80088),
            .I(N__80057));
    LocalMux I__18970 (
            .O(N__80085),
            .I(N__80052));
    LocalMux I__18969 (
            .O(N__80082),
            .I(N__80052));
    InMux I__18968 (
            .O(N__80081),
            .I(N__80049));
    Span4Mux_v I__18967 (
            .O(N__80078),
            .I(N__80046));
    LocalMux I__18966 (
            .O(N__80075),
            .I(N__80041));
    InMux I__18965 (
            .O(N__80074),
            .I(N__80038));
    LocalMux I__18964 (
            .O(N__80071),
            .I(N__80034));
    Span4Mux_v I__18963 (
            .O(N__80068),
            .I(N__80031));
    Span4Mux_v I__18962 (
            .O(N__80063),
            .I(N__80028));
    LocalMux I__18961 (
            .O(N__80060),
            .I(N__80025));
    LocalMux I__18960 (
            .O(N__80057),
            .I(N__80022));
    Span4Mux_v I__18959 (
            .O(N__80052),
            .I(N__80019));
    LocalMux I__18958 (
            .O(N__80049),
            .I(N__80014));
    Sp12to4 I__18957 (
            .O(N__80046),
            .I(N__80014));
    InMux I__18956 (
            .O(N__80045),
            .I(N__80009));
    InMux I__18955 (
            .O(N__80044),
            .I(N__80009));
    Span4Mux_h I__18954 (
            .O(N__80041),
            .I(N__80004));
    LocalMux I__18953 (
            .O(N__80038),
            .I(N__80004));
    InMux I__18952 (
            .O(N__80037),
            .I(N__80000));
    Span4Mux_v I__18951 (
            .O(N__80034),
            .I(N__79995));
    Span4Mux_h I__18950 (
            .O(N__80031),
            .I(N__79995));
    Sp12to4 I__18949 (
            .O(N__80028),
            .I(N__79990));
    Span12Mux_v I__18948 (
            .O(N__80025),
            .I(N__79990));
    Span12Mux_s8_h I__18947 (
            .O(N__80022),
            .I(N__79983));
    Sp12to4 I__18946 (
            .O(N__80019),
            .I(N__79983));
    Span12Mux_h I__18945 (
            .O(N__80014),
            .I(N__79983));
    LocalMux I__18944 (
            .O(N__80009),
            .I(N__79978));
    Span4Mux_h I__18943 (
            .O(N__80004),
            .I(N__79978));
    InMux I__18942 (
            .O(N__80003),
            .I(N__79975));
    LocalMux I__18941 (
            .O(N__80000),
            .I(uart_pc_data_5));
    Odrv4 I__18940 (
            .O(N__79995),
            .I(uart_pc_data_5));
    Odrv12 I__18939 (
            .O(N__79990),
            .I(uart_pc_data_5));
    Odrv12 I__18938 (
            .O(N__79983),
            .I(uart_pc_data_5));
    Odrv4 I__18937 (
            .O(N__79978),
            .I(uart_pc_data_5));
    LocalMux I__18936 (
            .O(N__79975),
            .I(uart_pc_data_5));
    InMux I__18935 (
            .O(N__79962),
            .I(N__79958));
    InMux I__18934 (
            .O(N__79961),
            .I(N__79955));
    LocalMux I__18933 (
            .O(N__79958),
            .I(N__79952));
    LocalMux I__18932 (
            .O(N__79955),
            .I(N__79949));
    Span4Mux_v I__18931 (
            .O(N__79952),
            .I(N__79946));
    Span4Mux_v I__18930 (
            .O(N__79949),
            .I(N__79943));
    Span4Mux_v I__18929 (
            .O(N__79946),
            .I(N__79938));
    Span4Mux_s0_h I__18928 (
            .O(N__79943),
            .I(N__79938));
    Sp12to4 I__18927 (
            .O(N__79938),
            .I(N__79935));
    Odrv12 I__18926 (
            .O(N__79935),
            .I(xy_kd_5));
    InMux I__18925 (
            .O(N__79932),
            .I(N__79927));
    InMux I__18924 (
            .O(N__79931),
            .I(N__79924));
    InMux I__18923 (
            .O(N__79930),
            .I(N__79921));
    LocalMux I__18922 (
            .O(N__79927),
            .I(N__79918));
    LocalMux I__18921 (
            .O(N__79924),
            .I(N__79915));
    LocalMux I__18920 (
            .O(N__79921),
            .I(N__79910));
    Span4Mux_v I__18919 (
            .O(N__79918),
            .I(N__79910));
    Span4Mux_v I__18918 (
            .O(N__79915),
            .I(N__79905));
    Span4Mux_v I__18917 (
            .O(N__79910),
            .I(N__79902));
    InMux I__18916 (
            .O(N__79909),
            .I(N__79899));
    InMux I__18915 (
            .O(N__79908),
            .I(N__79896));
    Span4Mux_h I__18914 (
            .O(N__79905),
            .I(N__79893));
    Span4Mux_v I__18913 (
            .O(N__79902),
            .I(N__79885));
    LocalMux I__18912 (
            .O(N__79899),
            .I(N__79882));
    LocalMux I__18911 (
            .O(N__79896),
            .I(N__79877));
    Span4Mux_h I__18910 (
            .O(N__79893),
            .I(N__79877));
    InMux I__18909 (
            .O(N__79892),
            .I(N__79874));
    InMux I__18908 (
            .O(N__79891),
            .I(N__79871));
    InMux I__18907 (
            .O(N__79890),
            .I(N__79867));
    InMux I__18906 (
            .O(N__79889),
            .I(N__79861));
    InMux I__18905 (
            .O(N__79888),
            .I(N__79858));
    Span4Mux_v I__18904 (
            .O(N__79885),
            .I(N__79852));
    Span4Mux_s3_h I__18903 (
            .O(N__79882),
            .I(N__79852));
    Span4Mux_v I__18902 (
            .O(N__79877),
            .I(N__79847));
    LocalMux I__18901 (
            .O(N__79874),
            .I(N__79847));
    LocalMux I__18900 (
            .O(N__79871),
            .I(N__79844));
    InMux I__18899 (
            .O(N__79870),
            .I(N__79841));
    LocalMux I__18898 (
            .O(N__79867),
            .I(N__79838));
    InMux I__18897 (
            .O(N__79866),
            .I(N__79832));
    InMux I__18896 (
            .O(N__79865),
            .I(N__79832));
    InMux I__18895 (
            .O(N__79864),
            .I(N__79829));
    LocalMux I__18894 (
            .O(N__79861),
            .I(N__79826));
    LocalMux I__18893 (
            .O(N__79858),
            .I(N__79823));
    InMux I__18892 (
            .O(N__79857),
            .I(N__79820));
    Span4Mux_v I__18891 (
            .O(N__79852),
            .I(N__79817));
    Span4Mux_h I__18890 (
            .O(N__79847),
            .I(N__79814));
    Span4Mux_v I__18889 (
            .O(N__79844),
            .I(N__79809));
    LocalMux I__18888 (
            .O(N__79841),
            .I(N__79809));
    Span4Mux_h I__18887 (
            .O(N__79838),
            .I(N__79806));
    CascadeMux I__18886 (
            .O(N__79837),
            .I(N__79803));
    LocalMux I__18885 (
            .O(N__79832),
            .I(N__79800));
    LocalMux I__18884 (
            .O(N__79829),
            .I(N__79797));
    Span12Mux_v I__18883 (
            .O(N__79826),
            .I(N__79794));
    Span4Mux_h I__18882 (
            .O(N__79823),
            .I(N__79791));
    LocalMux I__18881 (
            .O(N__79820),
            .I(N__79784));
    Span4Mux_h I__18880 (
            .O(N__79817),
            .I(N__79784));
    Span4Mux_v I__18879 (
            .O(N__79814),
            .I(N__79784));
    Span4Mux_v I__18878 (
            .O(N__79809),
            .I(N__79779));
    Span4Mux_h I__18877 (
            .O(N__79806),
            .I(N__79779));
    InMux I__18876 (
            .O(N__79803),
            .I(N__79776));
    Span4Mux_v I__18875 (
            .O(N__79800),
            .I(N__79771));
    Span4Mux_v I__18874 (
            .O(N__79797),
            .I(N__79771));
    Odrv12 I__18873 (
            .O(N__79794),
            .I(uart_pc_data_7));
    Odrv4 I__18872 (
            .O(N__79791),
            .I(uart_pc_data_7));
    Odrv4 I__18871 (
            .O(N__79784),
            .I(uart_pc_data_7));
    Odrv4 I__18870 (
            .O(N__79779),
            .I(uart_pc_data_7));
    LocalMux I__18869 (
            .O(N__79776),
            .I(uart_pc_data_7));
    Odrv4 I__18868 (
            .O(N__79771),
            .I(uart_pc_data_7));
    InMux I__18867 (
            .O(N__79758),
            .I(N__79755));
    LocalMux I__18866 (
            .O(N__79755),
            .I(N__79751));
    InMux I__18865 (
            .O(N__79754),
            .I(N__79748));
    Span4Mux_s2_h I__18864 (
            .O(N__79751),
            .I(N__79745));
    LocalMux I__18863 (
            .O(N__79748),
            .I(N__79742));
    Span4Mux_v I__18862 (
            .O(N__79745),
            .I(N__79737));
    Span4Mux_s2_h I__18861 (
            .O(N__79742),
            .I(N__79737));
    Odrv4 I__18860 (
            .O(N__79737),
            .I(xy_kd_7));
    InMux I__18859 (
            .O(N__79734),
            .I(N__79731));
    LocalMux I__18858 (
            .O(N__79731),
            .I(N__79727));
    InMux I__18857 (
            .O(N__79730),
            .I(N__79721));
    Span4Mux_v I__18856 (
            .O(N__79727),
            .I(N__79717));
    InMux I__18855 (
            .O(N__79726),
            .I(N__79710));
    InMux I__18854 (
            .O(N__79725),
            .I(N__79707));
    InMux I__18853 (
            .O(N__79724),
            .I(N__79704));
    LocalMux I__18852 (
            .O(N__79721),
            .I(N__79701));
    InMux I__18851 (
            .O(N__79720),
            .I(N__79698));
    Span4Mux_v I__18850 (
            .O(N__79717),
            .I(N__79694));
    InMux I__18849 (
            .O(N__79716),
            .I(N__79691));
    InMux I__18848 (
            .O(N__79715),
            .I(N__79688));
    InMux I__18847 (
            .O(N__79714),
            .I(N__79685));
    InMux I__18846 (
            .O(N__79713),
            .I(N__79681));
    LocalMux I__18845 (
            .O(N__79710),
            .I(N__79678));
    LocalMux I__18844 (
            .O(N__79707),
            .I(N__79675));
    LocalMux I__18843 (
            .O(N__79704),
            .I(N__79672));
    Span12Mux_s9_v I__18842 (
            .O(N__79701),
            .I(N__79669));
    LocalMux I__18841 (
            .O(N__79698),
            .I(N__79666));
    InMux I__18840 (
            .O(N__79697),
            .I(N__79663));
    Sp12to4 I__18839 (
            .O(N__79694),
            .I(N__79658));
    LocalMux I__18838 (
            .O(N__79691),
            .I(N__79658));
    LocalMux I__18837 (
            .O(N__79688),
            .I(N__79655));
    LocalMux I__18836 (
            .O(N__79685),
            .I(N__79652));
    InMux I__18835 (
            .O(N__79684),
            .I(N__79649));
    LocalMux I__18834 (
            .O(N__79681),
            .I(N__79644));
    Span4Mux_h I__18833 (
            .O(N__79678),
            .I(N__79644));
    Span4Mux_v I__18832 (
            .O(N__79675),
            .I(N__79641));
    Span12Mux_s11_h I__18831 (
            .O(N__79672),
            .I(N__79636));
    Span12Mux_h I__18830 (
            .O(N__79669),
            .I(N__79636));
    Sp12to4 I__18829 (
            .O(N__79666),
            .I(N__79631));
    LocalMux I__18828 (
            .O(N__79663),
            .I(N__79631));
    Span12Mux_h I__18827 (
            .O(N__79658),
            .I(N__79623));
    Span12Mux_s7_h I__18826 (
            .O(N__79655),
            .I(N__79623));
    Span12Mux_v I__18825 (
            .O(N__79652),
            .I(N__79623));
    LocalMux I__18824 (
            .O(N__79649),
            .I(N__79618));
    Span4Mux_v I__18823 (
            .O(N__79644),
            .I(N__79618));
    Sp12to4 I__18822 (
            .O(N__79641),
            .I(N__79611));
    Span12Mux_v I__18821 (
            .O(N__79636),
            .I(N__79611));
    Span12Mux_s8_v I__18820 (
            .O(N__79631),
            .I(N__79611));
    InMux I__18819 (
            .O(N__79630),
            .I(N__79608));
    Odrv12 I__18818 (
            .O(N__79623),
            .I(uart_pc_data_3));
    Odrv4 I__18817 (
            .O(N__79618),
            .I(uart_pc_data_3));
    Odrv12 I__18816 (
            .O(N__79611),
            .I(uart_pc_data_3));
    LocalMux I__18815 (
            .O(N__79608),
            .I(uart_pc_data_3));
    InMux I__18814 (
            .O(N__79599),
            .I(N__79596));
    LocalMux I__18813 (
            .O(N__79596),
            .I(N__79592));
    InMux I__18812 (
            .O(N__79595),
            .I(N__79589));
    Span4Mux_s2_h I__18811 (
            .O(N__79592),
            .I(N__79586));
    LocalMux I__18810 (
            .O(N__79589),
            .I(N__79583));
    Span4Mux_v I__18809 (
            .O(N__79586),
            .I(N__79578));
    Span4Mux_s2_h I__18808 (
            .O(N__79583),
            .I(N__79578));
    Odrv4 I__18807 (
            .O(N__79578),
            .I(xy_kd_3));
    InMux I__18806 (
            .O(N__79575),
            .I(N__79572));
    LocalMux I__18805 (
            .O(N__79572),
            .I(N__79569));
    Span4Mux_v I__18804 (
            .O(N__79569),
            .I(N__79566));
    Odrv4 I__18803 (
            .O(N__79566),
            .I(\pid_side.O_1_5 ));
    InMux I__18802 (
            .O(N__79563),
            .I(N__79554));
    InMux I__18801 (
            .O(N__79562),
            .I(N__79554));
    InMux I__18800 (
            .O(N__79561),
            .I(N__79554));
    LocalMux I__18799 (
            .O(N__79554),
            .I(N__79551));
    Span4Mux_h I__18798 (
            .O(N__79551),
            .I(N__79548));
    Span4Mux_h I__18797 (
            .O(N__79548),
            .I(N__79545));
    Odrv4 I__18796 (
            .O(N__79545),
            .I(\pid_side.error_d_regZ0Z_3 ));
    InMux I__18795 (
            .O(N__79542),
            .I(N__79539));
    LocalMux I__18794 (
            .O(N__79539),
            .I(N__79536));
    Span4Mux_v I__18793 (
            .O(N__79536),
            .I(N__79533));
    Odrv4 I__18792 (
            .O(N__79533),
            .I(\pid_side.O_1_6 ));
    InMux I__18791 (
            .O(N__79530),
            .I(N__79527));
    LocalMux I__18790 (
            .O(N__79527),
            .I(N__79523));
    InMux I__18789 (
            .O(N__79526),
            .I(N__79519));
    Span4Mux_h I__18788 (
            .O(N__79523),
            .I(N__79516));
    InMux I__18787 (
            .O(N__79522),
            .I(N__79513));
    LocalMux I__18786 (
            .O(N__79519),
            .I(N__79510));
    Odrv4 I__18785 (
            .O(N__79516),
            .I(\pid_side.error_d_regZ0Z_4 ));
    LocalMux I__18784 (
            .O(N__79513),
            .I(\pid_side.error_d_regZ0Z_4 ));
    Odrv4 I__18783 (
            .O(N__79510),
            .I(\pid_side.error_d_regZ0Z_4 ));
    InMux I__18782 (
            .O(N__79503),
            .I(N__79499));
    InMux I__18781 (
            .O(N__79502),
            .I(N__79496));
    LocalMux I__18780 (
            .O(N__79499),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    LocalMux I__18779 (
            .O(N__79496),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    InMux I__18778 (
            .O(N__79491),
            .I(N__79485));
    InMux I__18777 (
            .O(N__79490),
            .I(N__79485));
    LocalMux I__18776 (
            .O(N__79485),
            .I(N__79482));
    Odrv12 I__18775 (
            .O(N__79482),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ));
    InMux I__18774 (
            .O(N__79479),
            .I(N__79473));
    InMux I__18773 (
            .O(N__79478),
            .I(N__79473));
    LocalMux I__18772 (
            .O(N__79473),
            .I(\pid_side.error_d_reg_prevZ0Z_16 ));
    InMux I__18771 (
            .O(N__79470),
            .I(N__79467));
    LocalMux I__18770 (
            .O(N__79467),
            .I(N__79463));
    InMux I__18769 (
            .O(N__79466),
            .I(N__79460));
    Span4Mux_h I__18768 (
            .O(N__79463),
            .I(N__79457));
    LocalMux I__18767 (
            .O(N__79460),
            .I(N__79454));
    Odrv4 I__18766 (
            .O(N__79457),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ));
    Odrv12 I__18765 (
            .O(N__79454),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ));
    InMux I__18764 (
            .O(N__79449),
            .I(N__79446));
    LocalMux I__18763 (
            .O(N__79446),
            .I(N__79442));
    InMux I__18762 (
            .O(N__79445),
            .I(N__79439));
    Span4Mux_v I__18761 (
            .O(N__79442),
            .I(N__79436));
    LocalMux I__18760 (
            .O(N__79439),
            .I(N__79433));
    Span4Mux_h I__18759 (
            .O(N__79436),
            .I(N__79430));
    Span12Mux_v I__18758 (
            .O(N__79433),
            .I(N__79427));
    Odrv4 I__18757 (
            .O(N__79430),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ));
    Odrv12 I__18756 (
            .O(N__79427),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ));
    InMux I__18755 (
            .O(N__79422),
            .I(N__79419));
    LocalMux I__18754 (
            .O(N__79419),
            .I(N__79416));
    Span4Mux_h I__18753 (
            .O(N__79416),
            .I(N__79412));
    InMux I__18752 (
            .O(N__79415),
            .I(N__79407));
    Span4Mux_h I__18751 (
            .O(N__79412),
            .I(N__79403));
    InMux I__18750 (
            .O(N__79411),
            .I(N__79398));
    InMux I__18749 (
            .O(N__79410),
            .I(N__79398));
    LocalMux I__18748 (
            .O(N__79407),
            .I(N__79395));
    InMux I__18747 (
            .O(N__79406),
            .I(N__79392));
    Odrv4 I__18746 (
            .O(N__79403),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    LocalMux I__18745 (
            .O(N__79398),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    Odrv12 I__18744 (
            .O(N__79395),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    LocalMux I__18743 (
            .O(N__79392),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ));
    CascadeMux I__18742 (
            .O(N__79383),
            .I(\pid_side.un1_pid_prereg_167_0_1_cascade_ ));
    InMux I__18741 (
            .O(N__79380),
            .I(N__79377));
    LocalMux I__18740 (
            .O(N__79377),
            .I(N__79374));
    Odrv12 I__18739 (
            .O(N__79374),
            .I(\pid_side.un1_pid_prereg_167_0 ));
    InMux I__18738 (
            .O(N__79371),
            .I(N__79364));
    InMux I__18737 (
            .O(N__79370),
            .I(N__79364));
    InMux I__18736 (
            .O(N__79369),
            .I(N__79361));
    LocalMux I__18735 (
            .O(N__79364),
            .I(N__79358));
    LocalMux I__18734 (
            .O(N__79361),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__18733 (
            .O(N__79358),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    CascadeMux I__18732 (
            .O(N__79353),
            .I(N__79350));
    InMux I__18731 (
            .O(N__79350),
            .I(N__79347));
    LocalMux I__18730 (
            .O(N__79347),
            .I(N__79344));
    Sp12to4 I__18729 (
            .O(N__79344),
            .I(N__79341));
    Odrv12 I__18728 (
            .O(N__79341),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIOZ0Z_13 ));
    InMux I__18727 (
            .O(N__79338),
            .I(N__79334));
    InMux I__18726 (
            .O(N__79337),
            .I(N__79331));
    LocalMux I__18725 (
            .O(N__79334),
            .I(N__79328));
    LocalMux I__18724 (
            .O(N__79331),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    Odrv4 I__18723 (
            .O(N__79328),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    InMux I__18722 (
            .O(N__79323),
            .I(N__79320));
    LocalMux I__18721 (
            .O(N__79320),
            .I(N__79317));
    Span4Mux_v I__18720 (
            .O(N__79317),
            .I(N__79313));
    InMux I__18719 (
            .O(N__79316),
            .I(N__79310));
    Span4Mux_h I__18718 (
            .O(N__79313),
            .I(N__79305));
    LocalMux I__18717 (
            .O(N__79310),
            .I(N__79305));
    Odrv4 I__18716 (
            .O(N__79305),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ));
    InMux I__18715 (
            .O(N__79302),
            .I(N__79299));
    LocalMux I__18714 (
            .O(N__79299),
            .I(\pid_side.error_d_reg_prev_esr_RNIMERG_0Z0Z_12 ));
    InMux I__18713 (
            .O(N__79296),
            .I(N__79293));
    LocalMux I__18712 (
            .O(N__79293),
            .I(\pid_side.error_p_reg_esr_RNIR3TQ1Z0Z_12 ));
    InMux I__18711 (
            .O(N__79290),
            .I(N__79285));
    InMux I__18710 (
            .O(N__79289),
            .I(N__79281));
    InMux I__18709 (
            .O(N__79288),
            .I(N__79278));
    LocalMux I__18708 (
            .O(N__79285),
            .I(N__79272));
    InMux I__18707 (
            .O(N__79284),
            .I(N__79269));
    LocalMux I__18706 (
            .O(N__79281),
            .I(N__79265));
    LocalMux I__18705 (
            .O(N__79278),
            .I(N__79262));
    InMux I__18704 (
            .O(N__79277),
            .I(N__79259));
    InMux I__18703 (
            .O(N__79276),
            .I(N__79255));
    InMux I__18702 (
            .O(N__79275),
            .I(N__79252));
    Span4Mux_v I__18701 (
            .O(N__79272),
            .I(N__79249));
    LocalMux I__18700 (
            .O(N__79269),
            .I(N__79246));
    InMux I__18699 (
            .O(N__79268),
            .I(N__79243));
    Span4Mux_v I__18698 (
            .O(N__79265),
            .I(N__79239));
    Span4Mux_h I__18697 (
            .O(N__79262),
            .I(N__79234));
    LocalMux I__18696 (
            .O(N__79259),
            .I(N__79234));
    InMux I__18695 (
            .O(N__79258),
            .I(N__79231));
    LocalMux I__18694 (
            .O(N__79255),
            .I(N__79228));
    LocalMux I__18693 (
            .O(N__79252),
            .I(N__79224));
    Sp12to4 I__18692 (
            .O(N__79249),
            .I(N__79221));
    Span4Mux_h I__18691 (
            .O(N__79246),
            .I(N__79216));
    LocalMux I__18690 (
            .O(N__79243),
            .I(N__79216));
    InMux I__18689 (
            .O(N__79242),
            .I(N__79213));
    Span4Mux_v I__18688 (
            .O(N__79239),
            .I(N__79208));
    Span4Mux_h I__18687 (
            .O(N__79234),
            .I(N__79208));
    LocalMux I__18686 (
            .O(N__79231),
            .I(N__79205));
    Span4Mux_h I__18685 (
            .O(N__79228),
            .I(N__79202));
    InMux I__18684 (
            .O(N__79227),
            .I(N__79199));
    Span12Mux_h I__18683 (
            .O(N__79224),
            .I(N__79192));
    Span12Mux_s9_h I__18682 (
            .O(N__79221),
            .I(N__79192));
    Span4Mux_v I__18681 (
            .O(N__79216),
            .I(N__79187));
    LocalMux I__18680 (
            .O(N__79213),
            .I(N__79187));
    Span4Mux_v I__18679 (
            .O(N__79208),
            .I(N__79184));
    Span4Mux_h I__18678 (
            .O(N__79205),
            .I(N__79181));
    Span4Mux_h I__18677 (
            .O(N__79202),
            .I(N__79176));
    LocalMux I__18676 (
            .O(N__79199),
            .I(N__79176));
    InMux I__18675 (
            .O(N__79198),
            .I(N__79173));
    InMux I__18674 (
            .O(N__79197),
            .I(N__79170));
    Span12Mux_v I__18673 (
            .O(N__79192),
            .I(N__79167));
    Span4Mux_h I__18672 (
            .O(N__79187),
            .I(N__79160));
    Span4Mux_v I__18671 (
            .O(N__79184),
            .I(N__79160));
    Span4Mux_h I__18670 (
            .O(N__79181),
            .I(N__79160));
    Span4Mux_v I__18669 (
            .O(N__79176),
            .I(N__79155));
    LocalMux I__18668 (
            .O(N__79173),
            .I(N__79155));
    LocalMux I__18667 (
            .O(N__79170),
            .I(uart_pc_data_4));
    Odrv12 I__18666 (
            .O(N__79167),
            .I(uart_pc_data_4));
    Odrv4 I__18665 (
            .O(N__79160),
            .I(uart_pc_data_4));
    Odrv4 I__18664 (
            .O(N__79155),
            .I(uart_pc_data_4));
    InMux I__18663 (
            .O(N__79146),
            .I(N__79143));
    LocalMux I__18662 (
            .O(N__79143),
            .I(N__79139));
    InMux I__18661 (
            .O(N__79142),
            .I(N__79136));
    Span4Mux_s3_h I__18660 (
            .O(N__79139),
            .I(N__79133));
    LocalMux I__18659 (
            .O(N__79136),
            .I(N__79130));
    Span4Mux_v I__18658 (
            .O(N__79133),
            .I(N__79125));
    Span4Mux_s3_h I__18657 (
            .O(N__79130),
            .I(N__79125));
    Odrv4 I__18656 (
            .O(N__79125),
            .I(xy_kd_4));
    InMux I__18655 (
            .O(N__79122),
            .I(N__79116));
    InMux I__18654 (
            .O(N__79121),
            .I(N__79116));
    LocalMux I__18653 (
            .O(N__79116),
            .I(N__79113));
    Span4Mux_h I__18652 (
            .O(N__79113),
            .I(N__79110));
    Odrv4 I__18651 (
            .O(N__79110),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ));
    InMux I__18650 (
            .O(N__79107),
            .I(N__79103));
    InMux I__18649 (
            .O(N__79106),
            .I(N__79100));
    LocalMux I__18648 (
            .O(N__79103),
            .I(\pid_side.error_d_reg_prevZ0Z_4 ));
    LocalMux I__18647 (
            .O(N__79100),
            .I(\pid_side.error_d_reg_prevZ0Z_4 ));
    InMux I__18646 (
            .O(N__79095),
            .I(N__79091));
    InMux I__18645 (
            .O(N__79094),
            .I(N__79088));
    LocalMux I__18644 (
            .O(N__79091),
            .I(\pid_side.error_p_regZ0Z_4 ));
    LocalMux I__18643 (
            .O(N__79088),
            .I(\pid_side.error_p_regZ0Z_4 ));
    InMux I__18642 (
            .O(N__79083),
            .I(N__79077));
    InMux I__18641 (
            .O(N__79082),
            .I(N__79077));
    LocalMux I__18640 (
            .O(N__79077),
            .I(N__79074));
    Odrv12 I__18639 (
            .O(N__79074),
            .I(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ));
    InMux I__18638 (
            .O(N__79071),
            .I(N__79068));
    LocalMux I__18637 (
            .O(N__79068),
            .I(N__79065));
    Span4Mux_v I__18636 (
            .O(N__79065),
            .I(N__79061));
    InMux I__18635 (
            .O(N__79064),
            .I(N__79058));
    Span4Mux_h I__18634 (
            .O(N__79061),
            .I(N__79053));
    LocalMux I__18633 (
            .O(N__79058),
            .I(N__79053));
    Span4Mux_h I__18632 (
            .O(N__79053),
            .I(N__79050));
    Odrv4 I__18631 (
            .O(N__79050),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ));
    InMux I__18630 (
            .O(N__79047),
            .I(N__79044));
    LocalMux I__18629 (
            .O(N__79044),
            .I(N__79040));
    InMux I__18628 (
            .O(N__79043),
            .I(N__79037));
    Span4Mux_v I__18627 (
            .O(N__79040),
            .I(N__79032));
    LocalMux I__18626 (
            .O(N__79037),
            .I(N__79032));
    Span4Mux_h I__18625 (
            .O(N__79032),
            .I(N__79029));
    Span4Mux_h I__18624 (
            .O(N__79029),
            .I(N__79026));
    Odrv4 I__18623 (
            .O(N__79026),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ));
    InMux I__18622 (
            .O(N__79023),
            .I(N__79017));
    InMux I__18621 (
            .O(N__79022),
            .I(N__79017));
    LocalMux I__18620 (
            .O(N__79017),
            .I(\pid_side.error_d_reg_prevZ0Z_15 ));
    InMux I__18619 (
            .O(N__79014),
            .I(N__79008));
    InMux I__18618 (
            .O(N__79013),
            .I(N__79008));
    LocalMux I__18617 (
            .O(N__79008),
            .I(N__79005));
    Span4Mux_h I__18616 (
            .O(N__79005),
            .I(N__79002));
    Odrv4 I__18615 (
            .O(N__79002),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ));
    InMux I__18614 (
            .O(N__78999),
            .I(N__78993));
    InMux I__18613 (
            .O(N__78998),
            .I(N__78993));
    LocalMux I__18612 (
            .O(N__78993),
            .I(N__78990));
    Odrv12 I__18611 (
            .O(N__78990),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ));
    CascadeMux I__18610 (
            .O(N__78987),
            .I(\pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13_cascade_ ));
    InMux I__18609 (
            .O(N__78984),
            .I(N__78981));
    LocalMux I__18608 (
            .O(N__78981),
            .I(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12 ));
    InMux I__18607 (
            .O(N__78978),
            .I(N__78975));
    LocalMux I__18606 (
            .O(N__78975),
            .I(N__78970));
    InMux I__18605 (
            .O(N__78974),
            .I(N__78965));
    InMux I__18604 (
            .O(N__78973),
            .I(N__78965));
    Span12Mux_v I__18603 (
            .O(N__78970),
            .I(N__78959));
    LocalMux I__18602 (
            .O(N__78965),
            .I(N__78959));
    InMux I__18601 (
            .O(N__78964),
            .I(N__78956));
    Odrv12 I__18600 (
            .O(N__78959),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    LocalMux I__18599 (
            .O(N__78956),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    InMux I__18598 (
            .O(N__78951),
            .I(N__78946));
    InMux I__18597 (
            .O(N__78950),
            .I(N__78941));
    InMux I__18596 (
            .O(N__78949),
            .I(N__78941));
    LocalMux I__18595 (
            .O(N__78946),
            .I(N__78938));
    LocalMux I__18594 (
            .O(N__78941),
            .I(N__78935));
    Span4Mux_v I__18593 (
            .O(N__78938),
            .I(N__78930));
    Span4Mux_h I__18592 (
            .O(N__78935),
            .I(N__78930));
    Odrv4 I__18591 (
            .O(N__78930),
            .I(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ));
    CascadeMux I__18590 (
            .O(N__78927),
            .I(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ));
    InMux I__18589 (
            .O(N__78924),
            .I(N__78921));
    LocalMux I__18588 (
            .O(N__78921),
            .I(\pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12 ));
    InMux I__18587 (
            .O(N__78918),
            .I(N__78914));
    CascadeMux I__18586 (
            .O(N__78917),
            .I(N__78911));
    LocalMux I__18585 (
            .O(N__78914),
            .I(N__78908));
    InMux I__18584 (
            .O(N__78911),
            .I(N__78905));
    Span4Mux_h I__18583 (
            .O(N__78908),
            .I(N__78900));
    LocalMux I__18582 (
            .O(N__78905),
            .I(N__78900));
    Span4Mux_h I__18581 (
            .O(N__78900),
            .I(N__78897));
    Odrv4 I__18580 (
            .O(N__78897),
            .I(\pid_side.error_d_reg_prev_esr_RNIQ7S9AZ0Z_12 ));
    InMux I__18579 (
            .O(N__78894),
            .I(N__78891));
    LocalMux I__18578 (
            .O(N__78891),
            .I(N__78888));
    Span4Mux_h I__18577 (
            .O(N__78888),
            .I(N__78885));
    Odrv4 I__18576 (
            .O(N__78885),
            .I(\pid_side.O_1_10 ));
    InMux I__18575 (
            .O(N__78882),
            .I(N__78876));
    InMux I__18574 (
            .O(N__78881),
            .I(N__78869));
    InMux I__18573 (
            .O(N__78880),
            .I(N__78869));
    InMux I__18572 (
            .O(N__78879),
            .I(N__78869));
    LocalMux I__18571 (
            .O(N__78876),
            .I(\pid_side.error_d_regZ0Z_8 ));
    LocalMux I__18570 (
            .O(N__78869),
            .I(\pid_side.error_d_regZ0Z_8 ));
    CascadeMux I__18569 (
            .O(N__78864),
            .I(N__78860));
    CascadeMux I__18568 (
            .O(N__78863),
            .I(N__78857));
    InMux I__18567 (
            .O(N__78860),
            .I(N__78849));
    InMux I__18566 (
            .O(N__78857),
            .I(N__78849));
    InMux I__18565 (
            .O(N__78856),
            .I(N__78849));
    LocalMux I__18564 (
            .O(N__78849),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    InMux I__18563 (
            .O(N__78846),
            .I(N__78843));
    LocalMux I__18562 (
            .O(N__78843),
            .I(N__78840));
    Span4Mux_v I__18561 (
            .O(N__78840),
            .I(N__78837));
    Span4Mux_h I__18560 (
            .O(N__78837),
            .I(N__78834));
    Odrv4 I__18559 (
            .O(N__78834),
            .I(\pid_front.O_12 ));
    InMux I__18558 (
            .O(N__78831),
            .I(N__78825));
    InMux I__18557 (
            .O(N__78830),
            .I(N__78822));
    CascadeMux I__18556 (
            .O(N__78829),
            .I(N__78818));
    InMux I__18555 (
            .O(N__78828),
            .I(N__78814));
    LocalMux I__18554 (
            .O(N__78825),
            .I(N__78809));
    LocalMux I__18553 (
            .O(N__78822),
            .I(N__78809));
    InMux I__18552 (
            .O(N__78821),
            .I(N__78802));
    InMux I__18551 (
            .O(N__78818),
            .I(N__78802));
    InMux I__18550 (
            .O(N__78817),
            .I(N__78802));
    LocalMux I__18549 (
            .O(N__78814),
            .I(N__78795));
    Span4Mux_v I__18548 (
            .O(N__78809),
            .I(N__78795));
    LocalMux I__18547 (
            .O(N__78802),
            .I(N__78795));
    Span4Mux_h I__18546 (
            .O(N__78795),
            .I(N__78792));
    Span4Mux_h I__18545 (
            .O(N__78792),
            .I(N__78789));
    Odrv4 I__18544 (
            .O(N__78789),
            .I(\pid_front.error_d_regZ0Z_10 ));
    InMux I__18543 (
            .O(N__78786),
            .I(N__78783));
    LocalMux I__18542 (
            .O(N__78783),
            .I(N__78780));
    Span4Mux_h I__18541 (
            .O(N__78780),
            .I(N__78777));
    Span4Mux_v I__18540 (
            .O(N__78777),
            .I(N__78774));
    Odrv4 I__18539 (
            .O(N__78774),
            .I(\pid_front.O_14 ));
    InMux I__18538 (
            .O(N__78771),
            .I(N__78762));
    InMux I__18537 (
            .O(N__78770),
            .I(N__78753));
    InMux I__18536 (
            .O(N__78769),
            .I(N__78753));
    InMux I__18535 (
            .O(N__78768),
            .I(N__78753));
    InMux I__18534 (
            .O(N__78767),
            .I(N__78753));
    InMux I__18533 (
            .O(N__78766),
            .I(N__78750));
    InMux I__18532 (
            .O(N__78765),
            .I(N__78746));
    LocalMux I__18531 (
            .O(N__78762),
            .I(N__78743));
    LocalMux I__18530 (
            .O(N__78753),
            .I(N__78738));
    LocalMux I__18529 (
            .O(N__78750),
            .I(N__78738));
    InMux I__18528 (
            .O(N__78749),
            .I(N__78735));
    LocalMux I__18527 (
            .O(N__78746),
            .I(N__78728));
    Span4Mux_v I__18526 (
            .O(N__78743),
            .I(N__78728));
    Span4Mux_h I__18525 (
            .O(N__78738),
            .I(N__78728));
    LocalMux I__18524 (
            .O(N__78735),
            .I(N__78725));
    Span4Mux_h I__18523 (
            .O(N__78728),
            .I(N__78722));
    Span12Mux_h I__18522 (
            .O(N__78725),
            .I(N__78719));
    Span4Mux_h I__18521 (
            .O(N__78722),
            .I(N__78716));
    Odrv12 I__18520 (
            .O(N__78719),
            .I(\pid_front.error_d_regZ0Z_12 ));
    Odrv4 I__18519 (
            .O(N__78716),
            .I(\pid_front.error_d_regZ0Z_12 ));
    InMux I__18518 (
            .O(N__78711),
            .I(N__78708));
    LocalMux I__18517 (
            .O(N__78708),
            .I(N__78705));
    Span12Mux_h I__18516 (
            .O(N__78705),
            .I(N__78702));
    Odrv12 I__18515 (
            .O(N__78702),
            .I(\pid_front.O_15 ));
    InMux I__18514 (
            .O(N__78699),
            .I(N__78691));
    InMux I__18513 (
            .O(N__78698),
            .I(N__78691));
    InMux I__18512 (
            .O(N__78697),
            .I(N__78686));
    InMux I__18511 (
            .O(N__78696),
            .I(N__78686));
    LocalMux I__18510 (
            .O(N__78691),
            .I(N__78683));
    LocalMux I__18509 (
            .O(N__78686),
            .I(N__78680));
    Span4Mux_v I__18508 (
            .O(N__78683),
            .I(N__78675));
    Span4Mux_h I__18507 (
            .O(N__78680),
            .I(N__78675));
    Span4Mux_h I__18506 (
            .O(N__78675),
            .I(N__78672));
    Span4Mux_h I__18505 (
            .O(N__78672),
            .I(N__78669));
    Odrv4 I__18504 (
            .O(N__78669),
            .I(\pid_front.error_d_regZ0Z_13 ));
    InMux I__18503 (
            .O(N__78666),
            .I(N__78663));
    LocalMux I__18502 (
            .O(N__78663),
            .I(N__78660));
    Odrv12 I__18501 (
            .O(N__78660),
            .I(\pid_side.O_1_4 ));
    InMux I__18500 (
            .O(N__78657),
            .I(N__78651));
    InMux I__18499 (
            .O(N__78656),
            .I(N__78651));
    LocalMux I__18498 (
            .O(N__78651),
            .I(N__78648));
    Span4Mux_h I__18497 (
            .O(N__78648),
            .I(N__78644));
    InMux I__18496 (
            .O(N__78647),
            .I(N__78641));
    Odrv4 I__18495 (
            .O(N__78644),
            .I(\pid_side.error_d_regZ0Z_2 ));
    LocalMux I__18494 (
            .O(N__78641),
            .I(\pid_side.error_d_regZ0Z_2 ));
    InMux I__18493 (
            .O(N__78636),
            .I(N__78633));
    LocalMux I__18492 (
            .O(N__78633),
            .I(N__78630));
    Span4Mux_v I__18491 (
            .O(N__78630),
            .I(N__78627));
    Span4Mux_h I__18490 (
            .O(N__78627),
            .I(N__78624));
    Odrv4 I__18489 (
            .O(N__78624),
            .I(\pid_side.O_1_9 ));
    InMux I__18488 (
            .O(N__78621),
            .I(N__78615));
    InMux I__18487 (
            .O(N__78620),
            .I(N__78615));
    LocalMux I__18486 (
            .O(N__78615),
            .I(N__78610));
    InMux I__18485 (
            .O(N__78614),
            .I(N__78605));
    InMux I__18484 (
            .O(N__78613),
            .I(N__78605));
    Odrv4 I__18483 (
            .O(N__78610),
            .I(\pid_side.error_d_regZ0Z_7 ));
    LocalMux I__18482 (
            .O(N__78605),
            .I(\pid_side.error_d_regZ0Z_7 ));
    InMux I__18481 (
            .O(N__78600),
            .I(N__78597));
    LocalMux I__18480 (
            .O(N__78597),
            .I(N__78594));
    Span4Mux_h I__18479 (
            .O(N__78594),
            .I(N__78591));
    Odrv4 I__18478 (
            .O(N__78591),
            .I(\pid_side.O_1_11 ));
    InMux I__18477 (
            .O(N__78588),
            .I(N__78573));
    InMux I__18476 (
            .O(N__78587),
            .I(N__78573));
    InMux I__18475 (
            .O(N__78586),
            .I(N__78573));
    InMux I__18474 (
            .O(N__78585),
            .I(N__78573));
    InMux I__18473 (
            .O(N__78584),
            .I(N__78573));
    LocalMux I__18472 (
            .O(N__78573),
            .I(\pid_side.error_d_regZ0Z_9 ));
    InMux I__18471 (
            .O(N__78570),
            .I(N__78567));
    LocalMux I__18470 (
            .O(N__78567),
            .I(N__78564));
    Span4Mux_v I__18469 (
            .O(N__78564),
            .I(N__78561));
    Span4Mux_h I__18468 (
            .O(N__78561),
            .I(N__78558));
    Odrv4 I__18467 (
            .O(N__78558),
            .I(\pid_side.O_2_4 ));
    InMux I__18466 (
            .O(N__78555),
            .I(N__78552));
    LocalMux I__18465 (
            .O(N__78552),
            .I(N__78547));
    CascadeMux I__18464 (
            .O(N__78551),
            .I(N__78544));
    CascadeMux I__18463 (
            .O(N__78550),
            .I(N__78541));
    Span4Mux_h I__18462 (
            .O(N__78547),
            .I(N__78538));
    InMux I__18461 (
            .O(N__78544),
            .I(N__78533));
    InMux I__18460 (
            .O(N__78541),
            .I(N__78533));
    Odrv4 I__18459 (
            .O(N__78538),
            .I(\pid_side.error_p_regZ0Z_1 ));
    LocalMux I__18458 (
            .O(N__78533),
            .I(\pid_side.error_p_regZ0Z_1 ));
    InMux I__18457 (
            .O(N__78528),
            .I(N__78525));
    LocalMux I__18456 (
            .O(N__78525),
            .I(N__78522));
    Span4Mux_v I__18455 (
            .O(N__78522),
            .I(N__78519));
    Odrv4 I__18454 (
            .O(N__78519),
            .I(\pid_side.O_1_12 ));
    InMux I__18453 (
            .O(N__78516),
            .I(N__78510));
    InMux I__18452 (
            .O(N__78515),
            .I(N__78510));
    LocalMux I__18451 (
            .O(N__78510),
            .I(N__78503));
    InMux I__18450 (
            .O(N__78509),
            .I(N__78494));
    InMux I__18449 (
            .O(N__78508),
            .I(N__78494));
    InMux I__18448 (
            .O(N__78507),
            .I(N__78494));
    InMux I__18447 (
            .O(N__78506),
            .I(N__78494));
    Odrv4 I__18446 (
            .O(N__78503),
            .I(\pid_side.error_d_regZ0Z_10 ));
    LocalMux I__18445 (
            .O(N__78494),
            .I(\pid_side.error_d_regZ0Z_10 ));
    InMux I__18444 (
            .O(N__78489),
            .I(N__78486));
    LocalMux I__18443 (
            .O(N__78486),
            .I(N__78482));
    InMux I__18442 (
            .O(N__78485),
            .I(N__78479));
    Span4Mux_v I__18441 (
            .O(N__78482),
            .I(N__78474));
    LocalMux I__18440 (
            .O(N__78479),
            .I(N__78474));
    Span4Mux_h I__18439 (
            .O(N__78474),
            .I(N__78471));
    Odrv4 I__18438 (
            .O(N__78471),
            .I(\pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12 ));
    CascadeMux I__18437 (
            .O(N__78468),
            .I(\pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12_cascade_ ));
    CascadeMux I__18436 (
            .O(N__78465),
            .I(\pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12_cascade_ ));
    InMux I__18435 (
            .O(N__78462),
            .I(N__78459));
    LocalMux I__18434 (
            .O(N__78459),
            .I(N__78455));
    InMux I__18433 (
            .O(N__78458),
            .I(N__78452));
    Span4Mux_h I__18432 (
            .O(N__78455),
            .I(N__78447));
    LocalMux I__18431 (
            .O(N__78452),
            .I(N__78447));
    Span4Mux_v I__18430 (
            .O(N__78447),
            .I(N__78444));
    Odrv4 I__18429 (
            .O(N__78444),
            .I(\pid_side.un1_pid_prereg_0_axb_14 ));
    InMux I__18428 (
            .O(N__78441),
            .I(N__78438));
    LocalMux I__18427 (
            .O(N__78438),
            .I(N__78435));
    Span4Mux_h I__18426 (
            .O(N__78435),
            .I(N__78432));
    Odrv4 I__18425 (
            .O(N__78432),
            .I(\pid_side.O_1_7 ));
    InMux I__18424 (
            .O(N__78429),
            .I(N__78426));
    LocalMux I__18423 (
            .O(N__78426),
            .I(N__78423));
    Span4Mux_h I__18422 (
            .O(N__78423),
            .I(N__78420));
    Odrv4 I__18421 (
            .O(N__78420),
            .I(\pid_side.O_1_8 ));
    InMux I__18420 (
            .O(N__78417),
            .I(N__78405));
    InMux I__18419 (
            .O(N__78416),
            .I(N__78405));
    InMux I__18418 (
            .O(N__78415),
            .I(N__78405));
    InMux I__18417 (
            .O(N__78414),
            .I(N__78405));
    LocalMux I__18416 (
            .O(N__78405),
            .I(\pid_side.error_d_regZ0Z_6 ));
    InMux I__18415 (
            .O(N__78402),
            .I(N__78396));
    InMux I__18414 (
            .O(N__78401),
            .I(N__78396));
    LocalMux I__18413 (
            .O(N__78396),
            .I(\pid_side.N_1875_i ));
    CascadeMux I__18412 (
            .O(N__78393),
            .I(N__78390));
    InMux I__18411 (
            .O(N__78390),
            .I(N__78384));
    InMux I__18410 (
            .O(N__78389),
            .I(N__78384));
    LocalMux I__18409 (
            .O(N__78384),
            .I(N__78381));
    Span4Mux_v I__18408 (
            .O(N__78381),
            .I(N__78377));
    InMux I__18407 (
            .O(N__78380),
            .I(N__78374));
    Odrv4 I__18406 (
            .O(N__78377),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    LocalMux I__18405 (
            .O(N__78374),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    InMux I__18404 (
            .O(N__78369),
            .I(N__78365));
    InMux I__18403 (
            .O(N__78368),
            .I(N__78362));
    LocalMux I__18402 (
            .O(N__78365),
            .I(N__78349));
    LocalMux I__18401 (
            .O(N__78362),
            .I(N__78346));
    CEMux I__18400 (
            .O(N__78361),
            .I(N__78321));
    CEMux I__18399 (
            .O(N__78360),
            .I(N__78321));
    CEMux I__18398 (
            .O(N__78359),
            .I(N__78321));
    CEMux I__18397 (
            .O(N__78358),
            .I(N__78321));
    CEMux I__18396 (
            .O(N__78357),
            .I(N__78321));
    CEMux I__18395 (
            .O(N__78356),
            .I(N__78321));
    CEMux I__18394 (
            .O(N__78355),
            .I(N__78321));
    CEMux I__18393 (
            .O(N__78354),
            .I(N__78321));
    CEMux I__18392 (
            .O(N__78353),
            .I(N__78321));
    CEMux I__18391 (
            .O(N__78352),
            .I(N__78321));
    Glb2LocalMux I__18390 (
            .O(N__78349),
            .I(N__78321));
    Glb2LocalMux I__18389 (
            .O(N__78346),
            .I(N__78321));
    GlobalMux I__18388 (
            .O(N__78321),
            .I(N__78318));
    gio2CtrlBuf I__18387 (
            .O(N__78318),
            .I(\pid_side.N_478_g ));
    InMux I__18386 (
            .O(N__78315),
            .I(N__78308));
    InMux I__18385 (
            .O(N__78314),
            .I(N__78305));
    InMux I__18384 (
            .O(N__78313),
            .I(N__78298));
    InMux I__18383 (
            .O(N__78312),
            .I(N__78298));
    InMux I__18382 (
            .O(N__78311),
            .I(N__78298));
    LocalMux I__18381 (
            .O(N__78308),
            .I(\pid_side.error_d_regZ0Z_5 ));
    LocalMux I__18380 (
            .O(N__78305),
            .I(\pid_side.error_d_regZ0Z_5 ));
    LocalMux I__18379 (
            .O(N__78298),
            .I(\pid_side.error_d_regZ0Z_5 ));
    InMux I__18378 (
            .O(N__78291),
            .I(N__78285));
    InMux I__18377 (
            .O(N__78290),
            .I(N__78278));
    InMux I__18376 (
            .O(N__78289),
            .I(N__78278));
    InMux I__18375 (
            .O(N__78288),
            .I(N__78278));
    LocalMux I__18374 (
            .O(N__78285),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    LocalMux I__18373 (
            .O(N__78278),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    InMux I__18372 (
            .O(N__78273),
            .I(N__78270));
    LocalMux I__18371 (
            .O(N__78270),
            .I(N__78267));
    Sp12to4 I__18370 (
            .O(N__78267),
            .I(N__78263));
    InMux I__18369 (
            .O(N__78266),
            .I(N__78260));
    Span12Mux_v I__18368 (
            .O(N__78263),
            .I(N__78256));
    LocalMux I__18367 (
            .O(N__78260),
            .I(N__78253));
    InMux I__18366 (
            .O(N__78259),
            .I(N__78250));
    Odrv12 I__18365 (
            .O(N__78256),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    Odrv4 I__18364 (
            .O(N__78253),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    LocalMux I__18363 (
            .O(N__78250),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    InMux I__18362 (
            .O(N__78243),
            .I(N__78240));
    LocalMux I__18361 (
            .O(N__78240),
            .I(N__78237));
    Span4Mux_h I__18360 (
            .O(N__78237),
            .I(N__78234));
    Span4Mux_v I__18359 (
            .O(N__78234),
            .I(N__78231));
    Span4Mux_h I__18358 (
            .O(N__78231),
            .I(N__78224));
    InMux I__18357 (
            .O(N__78230),
            .I(N__78221));
    InMux I__18356 (
            .O(N__78229),
            .I(N__78216));
    InMux I__18355 (
            .O(N__78228),
            .I(N__78216));
    InMux I__18354 (
            .O(N__78227),
            .I(N__78213));
    Odrv4 I__18353 (
            .O(N__78224),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__18352 (
            .O(N__78221),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__18351 (
            .O(N__78216),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__18350 (
            .O(N__78213),
            .I(\ppm_encoder_1.N_221 ));
    InMux I__18349 (
            .O(N__78204),
            .I(N__78187));
    InMux I__18348 (
            .O(N__78203),
            .I(N__78187));
    InMux I__18347 (
            .O(N__78202),
            .I(N__78187));
    InMux I__18346 (
            .O(N__78201),
            .I(N__78187));
    InMux I__18345 (
            .O(N__78200),
            .I(N__78179));
    InMux I__18344 (
            .O(N__78199),
            .I(N__78169));
    InMux I__18343 (
            .O(N__78198),
            .I(N__78169));
    InMux I__18342 (
            .O(N__78197),
            .I(N__78169));
    InMux I__18341 (
            .O(N__78196),
            .I(N__78169));
    LocalMux I__18340 (
            .O(N__78187),
            .I(N__78166));
    InMux I__18339 (
            .O(N__78186),
            .I(N__78163));
    InMux I__18338 (
            .O(N__78185),
            .I(N__78154));
    InMux I__18337 (
            .O(N__78184),
            .I(N__78154));
    InMux I__18336 (
            .O(N__78183),
            .I(N__78154));
    InMux I__18335 (
            .O(N__78182),
            .I(N__78154));
    LocalMux I__18334 (
            .O(N__78179),
            .I(N__78151));
    InMux I__18333 (
            .O(N__78178),
            .I(N__78148));
    LocalMux I__18332 (
            .O(N__78169),
            .I(N__78145));
    Span4Mux_h I__18331 (
            .O(N__78166),
            .I(N__78138));
    LocalMux I__18330 (
            .O(N__78163),
            .I(N__78138));
    LocalMux I__18329 (
            .O(N__78154),
            .I(N__78138));
    Span4Mux_h I__18328 (
            .O(N__78151),
            .I(N__78135));
    LocalMux I__18327 (
            .O(N__78148),
            .I(N__78130));
    Span4Mux_h I__18326 (
            .O(N__78145),
            .I(N__78130));
    Span4Mux_h I__18325 (
            .O(N__78138),
            .I(N__78127));
    Span4Mux_v I__18324 (
            .O(N__78135),
            .I(N__78124));
    Sp12to4 I__18323 (
            .O(N__78130),
            .I(N__78121));
    Sp12to4 I__18322 (
            .O(N__78127),
            .I(N__78118));
    Sp12to4 I__18321 (
            .O(N__78124),
            .I(N__78113));
    Span12Mux_v I__18320 (
            .O(N__78121),
            .I(N__78113));
    Span12Mux_v I__18319 (
            .O(N__78118),
            .I(N__78110));
    Odrv12 I__18318 (
            .O(N__78113),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv12 I__18317 (
            .O(N__78110),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__18316 (
            .O(N__78105),
            .I(N__78102));
    LocalMux I__18315 (
            .O(N__78102),
            .I(N__78099));
    Odrv12 I__18314 (
            .O(N__78099),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__18313 (
            .O(N__78096),
            .I(N__78093));
    LocalMux I__18312 (
            .O(N__78093),
            .I(N__78090));
    Odrv4 I__18311 (
            .O(N__78090),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__18310 (
            .O(N__78087),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__18309 (
            .O(N__78084),
            .I(N__78081));
    LocalMux I__18308 (
            .O(N__78081),
            .I(N__78078));
    Span4Mux_h I__18307 (
            .O(N__78078),
            .I(N__78075));
    Span4Mux_v I__18306 (
            .O(N__78075),
            .I(N__78072));
    Span4Mux_v I__18305 (
            .O(N__78072),
            .I(N__78069));
    Span4Mux_h I__18304 (
            .O(N__78069),
            .I(N__78066));
    Odrv4 I__18303 (
            .O(N__78066),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ));
    CascadeMux I__18302 (
            .O(N__78063),
            .I(N__78060));
    InMux I__18301 (
            .O(N__78060),
            .I(N__78057));
    LocalMux I__18300 (
            .O(N__78057),
            .I(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ));
    InMux I__18299 (
            .O(N__78054),
            .I(N__78051));
    LocalMux I__18298 (
            .O(N__78051),
            .I(N__78048));
    Odrv4 I__18297 (
            .O(N__78048),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__18296 (
            .O(N__78045),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__18295 (
            .O(N__78042),
            .I(N__78039));
    LocalMux I__18294 (
            .O(N__78039),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__18293 (
            .O(N__78036),
            .I(N__78033));
    LocalMux I__18292 (
            .O(N__78033),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__18291 (
            .O(N__78030),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__18290 (
            .O(N__78027),
            .I(N__78024));
    LocalMux I__18289 (
            .O(N__78024),
            .I(N__78021));
    Span4Mux_v I__18288 (
            .O(N__78021),
            .I(N__78018));
    Sp12to4 I__18287 (
            .O(N__78018),
            .I(N__78015));
    Span12Mux_s11_h I__18286 (
            .O(N__78015),
            .I(N__78012));
    Odrv12 I__18285 (
            .O(N__78012),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__18284 (
            .O(N__78009),
            .I(N__78006));
    LocalMux I__18283 (
            .O(N__78006),
            .I(N__78003));
    Span4Mux_h I__18282 (
            .O(N__78003),
            .I(N__78000));
    Odrv4 I__18281 (
            .O(N__78000),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__18280 (
            .O(N__77997),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__18279 (
            .O(N__77994),
            .I(N__77991));
    LocalMux I__18278 (
            .O(N__77991),
            .I(N__77988));
    Span4Mux_v I__18277 (
            .O(N__77988),
            .I(N__77985));
    Span4Mux_h I__18276 (
            .O(N__77985),
            .I(N__77982));
    Odrv4 I__18275 (
            .O(N__77982),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__18274 (
            .O(N__77979),
            .I(N__77976));
    LocalMux I__18273 (
            .O(N__77976),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__18272 (
            .O(N__77973),
            .I(bfn_21_10_0_));
    InMux I__18271 (
            .O(N__77970),
            .I(N__77967));
    LocalMux I__18270 (
            .O(N__77967),
            .I(N__77964));
    Odrv4 I__18269 (
            .O(N__77964),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    CascadeMux I__18268 (
            .O(N__77961),
            .I(N__77958));
    InMux I__18267 (
            .O(N__77958),
            .I(N__77955));
    LocalMux I__18266 (
            .O(N__77955),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__18265 (
            .O(N__77952),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    CascadeMux I__18264 (
            .O(N__77949),
            .I(N__77945));
    CascadeMux I__18263 (
            .O(N__77948),
            .I(N__77942));
    InMux I__18262 (
            .O(N__77945),
            .I(N__77938));
    InMux I__18261 (
            .O(N__77942),
            .I(N__77935));
    InMux I__18260 (
            .O(N__77941),
            .I(N__77932));
    LocalMux I__18259 (
            .O(N__77938),
            .I(N__77929));
    LocalMux I__18258 (
            .O(N__77935),
            .I(N__77926));
    LocalMux I__18257 (
            .O(N__77932),
            .I(N__77923));
    Span4Mux_v I__18256 (
            .O(N__77929),
            .I(N__77918));
    Span4Mux_h I__18255 (
            .O(N__77926),
            .I(N__77918));
    Odrv4 I__18254 (
            .O(N__77923),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__18253 (
            .O(N__77918),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__18252 (
            .O(N__77913),
            .I(N__77910));
    LocalMux I__18251 (
            .O(N__77910),
            .I(N__77907));
    Span4Mux_v I__18250 (
            .O(N__77907),
            .I(N__77898));
    InMux I__18249 (
            .O(N__77906),
            .I(N__77893));
    InMux I__18248 (
            .O(N__77905),
            .I(N__77893));
    InMux I__18247 (
            .O(N__77904),
            .I(N__77884));
    InMux I__18246 (
            .O(N__77903),
            .I(N__77884));
    InMux I__18245 (
            .O(N__77902),
            .I(N__77884));
    InMux I__18244 (
            .O(N__77901),
            .I(N__77884));
    Odrv4 I__18243 (
            .O(N__77898),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    LocalMux I__18242 (
            .O(N__77893),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    LocalMux I__18241 (
            .O(N__77884),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    InMux I__18240 (
            .O(N__77877),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__18239 (
            .O(N__77874),
            .I(N__77871));
    LocalMux I__18238 (
            .O(N__77871),
            .I(N__77868));
    Odrv12 I__18237 (
            .O(N__77868),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__18236 (
            .O(N__77865),
            .I(N__77862));
    LocalMux I__18235 (
            .O(N__77862),
            .I(N__77859));
    Span4Mux_h I__18234 (
            .O(N__77859),
            .I(N__77856));
    Odrv4 I__18233 (
            .O(N__77856),
            .I(\pid_side.O_2_7 ));
    CascadeMux I__18232 (
            .O(N__77853),
            .I(N__77850));
    InMux I__18231 (
            .O(N__77850),
            .I(N__77847));
    LocalMux I__18230 (
            .O(N__77847),
            .I(N__77844));
    Span4Mux_h I__18229 (
            .O(N__77844),
            .I(N__77841));
    Odrv4 I__18228 (
            .O(N__77841),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__18227 (
            .O(N__77838),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__18226 (
            .O(N__77835),
            .I(N__77832));
    LocalMux I__18225 (
            .O(N__77832),
            .I(N__77829));
    Span4Mux_h I__18224 (
            .O(N__77829),
            .I(N__77826));
    Odrv4 I__18223 (
            .O(N__77826),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__18222 (
            .O(N__77823),
            .I(N__77820));
    LocalMux I__18221 (
            .O(N__77820),
            .I(N__77817));
    Span4Mux_v I__18220 (
            .O(N__77817),
            .I(N__77814));
    Odrv4 I__18219 (
            .O(N__77814),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__18218 (
            .O(N__77811),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__18217 (
            .O(N__77808),
            .I(N__77805));
    LocalMux I__18216 (
            .O(N__77805),
            .I(N__77802));
    Span12Mux_s10_h I__18215 (
            .O(N__77802),
            .I(N__77799));
    Span12Mux_v I__18214 (
            .O(N__77799),
            .I(N__77796));
    Odrv12 I__18213 (
            .O(N__77796),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ));
    CascadeMux I__18212 (
            .O(N__77793),
            .I(N__77790));
    InMux I__18211 (
            .O(N__77790),
            .I(N__77787));
    LocalMux I__18210 (
            .O(N__77787),
            .I(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ));
    InMux I__18209 (
            .O(N__77784),
            .I(N__77781));
    LocalMux I__18208 (
            .O(N__77781),
            .I(N__77778));
    Span4Mux_h I__18207 (
            .O(N__77778),
            .I(N__77775));
    Odrv4 I__18206 (
            .O(N__77775),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__18205 (
            .O(N__77772),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__18204 (
            .O(N__77769),
            .I(N__77766));
    LocalMux I__18203 (
            .O(N__77766),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    CascadeMux I__18202 (
            .O(N__77763),
            .I(N__77760));
    InMux I__18201 (
            .O(N__77760),
            .I(N__77757));
    LocalMux I__18200 (
            .O(N__77757),
            .I(N__77754));
    Span4Mux_h I__18199 (
            .O(N__77754),
            .I(N__77751));
    Odrv4 I__18198 (
            .O(N__77751),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__18197 (
            .O(N__77748),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__18196 (
            .O(N__77745),
            .I(N__77742));
    LocalMux I__18195 (
            .O(N__77742),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__18194 (
            .O(N__77739),
            .I(N__77736));
    LocalMux I__18193 (
            .O(N__77736),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__18192 (
            .O(N__77733),
            .I(bfn_21_9_0_));
    InMux I__18191 (
            .O(N__77730),
            .I(N__77727));
    LocalMux I__18190 (
            .O(N__77727),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__18189 (
            .O(N__77724),
            .I(N__77721));
    LocalMux I__18188 (
            .O(N__77721),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__18187 (
            .O(N__77718),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__18186 (
            .O(N__77715),
            .I(N__77712));
    LocalMux I__18185 (
            .O(N__77712),
            .I(N__77709));
    Span4Mux_h I__18184 (
            .O(N__77709),
            .I(N__77706));
    Odrv4 I__18183 (
            .O(N__77706),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__18182 (
            .O(N__77703),
            .I(N__77700));
    LocalMux I__18181 (
            .O(N__77700),
            .I(N__77697));
    Span4Mux_h I__18180 (
            .O(N__77697),
            .I(N__77694));
    Odrv4 I__18179 (
            .O(N__77694),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__18178 (
            .O(N__77691),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__18177 (
            .O(N__77688),
            .I(N__77685));
    LocalMux I__18176 (
            .O(N__77685),
            .I(N__77682));
    Odrv4 I__18175 (
            .O(N__77682),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__18174 (
            .O(N__77679),
            .I(N__77676));
    LocalMux I__18173 (
            .O(N__77676),
            .I(N__77673));
    Odrv4 I__18172 (
            .O(N__77673),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__18171 (
            .O(N__77670),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    CascadeMux I__18170 (
            .O(N__77667),
            .I(N__77650));
    CascadeMux I__18169 (
            .O(N__77666),
            .I(N__77643));
    CascadeMux I__18168 (
            .O(N__77665),
            .I(N__77597));
    CascadeMux I__18167 (
            .O(N__77664),
            .I(N__77594));
    InMux I__18166 (
            .O(N__77663),
            .I(N__77583));
    InMux I__18165 (
            .O(N__77662),
            .I(N__77580));
    InMux I__18164 (
            .O(N__77661),
            .I(N__77571));
    InMux I__18163 (
            .O(N__77660),
            .I(N__77571));
    InMux I__18162 (
            .O(N__77659),
            .I(N__77571));
    InMux I__18161 (
            .O(N__77658),
            .I(N__77571));
    InMux I__18160 (
            .O(N__77657),
            .I(N__77568));
    InMux I__18159 (
            .O(N__77656),
            .I(N__77563));
    InMux I__18158 (
            .O(N__77655),
            .I(N__77563));
    InMux I__18157 (
            .O(N__77654),
            .I(N__77560));
    InMux I__18156 (
            .O(N__77653),
            .I(N__77553));
    InMux I__18155 (
            .O(N__77650),
            .I(N__77553));
    InMux I__18154 (
            .O(N__77649),
            .I(N__77553));
    InMux I__18153 (
            .O(N__77648),
            .I(N__77546));
    InMux I__18152 (
            .O(N__77647),
            .I(N__77546));
    InMux I__18151 (
            .O(N__77646),
            .I(N__77546));
    InMux I__18150 (
            .O(N__77643),
            .I(N__77541));
    InMux I__18149 (
            .O(N__77642),
            .I(N__77541));
    InMux I__18148 (
            .O(N__77641),
            .I(N__77534));
    InMux I__18147 (
            .O(N__77640),
            .I(N__77534));
    InMux I__18146 (
            .O(N__77639),
            .I(N__77534));
    InMux I__18145 (
            .O(N__77638),
            .I(N__77525));
    InMux I__18144 (
            .O(N__77637),
            .I(N__77525));
    InMux I__18143 (
            .O(N__77636),
            .I(N__77525));
    InMux I__18142 (
            .O(N__77635),
            .I(N__77525));
    InMux I__18141 (
            .O(N__77634),
            .I(N__77522));
    InMux I__18140 (
            .O(N__77633),
            .I(N__77519));
    InMux I__18139 (
            .O(N__77632),
            .I(N__77516));
    InMux I__18138 (
            .O(N__77631),
            .I(N__77513));
    InMux I__18137 (
            .O(N__77630),
            .I(N__77510));
    InMux I__18136 (
            .O(N__77629),
            .I(N__77507));
    InMux I__18135 (
            .O(N__77628),
            .I(N__77500));
    InMux I__18134 (
            .O(N__77627),
            .I(N__77500));
    InMux I__18133 (
            .O(N__77626),
            .I(N__77500));
    InMux I__18132 (
            .O(N__77625),
            .I(N__77497));
    InMux I__18131 (
            .O(N__77624),
            .I(N__77492));
    InMux I__18130 (
            .O(N__77623),
            .I(N__77492));
    InMux I__18129 (
            .O(N__77622),
            .I(N__77487));
    InMux I__18128 (
            .O(N__77621),
            .I(N__77487));
    InMux I__18127 (
            .O(N__77620),
            .I(N__77484));
    InMux I__18126 (
            .O(N__77619),
            .I(N__77481));
    InMux I__18125 (
            .O(N__77618),
            .I(N__77478));
    InMux I__18124 (
            .O(N__77617),
            .I(N__77475));
    InMux I__18123 (
            .O(N__77616),
            .I(N__77472));
    InMux I__18122 (
            .O(N__77615),
            .I(N__77469));
    InMux I__18121 (
            .O(N__77614),
            .I(N__77462));
    InMux I__18120 (
            .O(N__77613),
            .I(N__77462));
    InMux I__18119 (
            .O(N__77612),
            .I(N__77462));
    InMux I__18118 (
            .O(N__77611),
            .I(N__77455));
    InMux I__18117 (
            .O(N__77610),
            .I(N__77455));
    InMux I__18116 (
            .O(N__77609),
            .I(N__77455));
    InMux I__18115 (
            .O(N__77608),
            .I(N__77452));
    InMux I__18114 (
            .O(N__77607),
            .I(N__77449));
    InMux I__18113 (
            .O(N__77606),
            .I(N__77446));
    InMux I__18112 (
            .O(N__77605),
            .I(N__77443));
    InMux I__18111 (
            .O(N__77604),
            .I(N__77440));
    InMux I__18110 (
            .O(N__77603),
            .I(N__77437));
    InMux I__18109 (
            .O(N__77602),
            .I(N__77434));
    InMux I__18108 (
            .O(N__77601),
            .I(N__77431));
    InMux I__18107 (
            .O(N__77600),
            .I(N__77422));
    InMux I__18106 (
            .O(N__77597),
            .I(N__77422));
    InMux I__18105 (
            .O(N__77594),
            .I(N__77422));
    InMux I__18104 (
            .O(N__77593),
            .I(N__77422));
    InMux I__18103 (
            .O(N__77592),
            .I(N__77415));
    InMux I__18102 (
            .O(N__77591),
            .I(N__77415));
    InMux I__18101 (
            .O(N__77590),
            .I(N__77415));
    InMux I__18100 (
            .O(N__77589),
            .I(N__77412));
    InMux I__18099 (
            .O(N__77588),
            .I(N__77409));
    InMux I__18098 (
            .O(N__77587),
            .I(N__77406));
    InMux I__18097 (
            .O(N__77586),
            .I(N__77403));
    LocalMux I__18096 (
            .O(N__77583),
            .I(N__77243));
    LocalMux I__18095 (
            .O(N__77580),
            .I(N__77240));
    LocalMux I__18094 (
            .O(N__77571),
            .I(N__77237));
    LocalMux I__18093 (
            .O(N__77568),
            .I(N__77234));
    LocalMux I__18092 (
            .O(N__77563),
            .I(N__77231));
    LocalMux I__18091 (
            .O(N__77560),
            .I(N__77228));
    LocalMux I__18090 (
            .O(N__77553),
            .I(N__77225));
    LocalMux I__18089 (
            .O(N__77546),
            .I(N__77222));
    LocalMux I__18088 (
            .O(N__77541),
            .I(N__77219));
    LocalMux I__18087 (
            .O(N__77534),
            .I(N__77216));
    LocalMux I__18086 (
            .O(N__77525),
            .I(N__77213));
    LocalMux I__18085 (
            .O(N__77522),
            .I(N__77210));
    LocalMux I__18084 (
            .O(N__77519),
            .I(N__77207));
    LocalMux I__18083 (
            .O(N__77516),
            .I(N__77204));
    LocalMux I__18082 (
            .O(N__77513),
            .I(N__77201));
    LocalMux I__18081 (
            .O(N__77510),
            .I(N__77198));
    LocalMux I__18080 (
            .O(N__77507),
            .I(N__77195));
    LocalMux I__18079 (
            .O(N__77500),
            .I(N__77192));
    LocalMux I__18078 (
            .O(N__77497),
            .I(N__77189));
    LocalMux I__18077 (
            .O(N__77492),
            .I(N__77186));
    LocalMux I__18076 (
            .O(N__77487),
            .I(N__77183));
    LocalMux I__18075 (
            .O(N__77484),
            .I(N__77180));
    LocalMux I__18074 (
            .O(N__77481),
            .I(N__77177));
    LocalMux I__18073 (
            .O(N__77478),
            .I(N__77174));
    LocalMux I__18072 (
            .O(N__77475),
            .I(N__77171));
    LocalMux I__18071 (
            .O(N__77472),
            .I(N__77168));
    LocalMux I__18070 (
            .O(N__77469),
            .I(N__77165));
    LocalMux I__18069 (
            .O(N__77462),
            .I(N__77162));
    LocalMux I__18068 (
            .O(N__77455),
            .I(N__77159));
    LocalMux I__18067 (
            .O(N__77452),
            .I(N__77156));
    LocalMux I__18066 (
            .O(N__77449),
            .I(N__77153));
    LocalMux I__18065 (
            .O(N__77446),
            .I(N__77150));
    LocalMux I__18064 (
            .O(N__77443),
            .I(N__77147));
    LocalMux I__18063 (
            .O(N__77440),
            .I(N__77144));
    LocalMux I__18062 (
            .O(N__77437),
            .I(N__77141));
    LocalMux I__18061 (
            .O(N__77434),
            .I(N__77138));
    LocalMux I__18060 (
            .O(N__77431),
            .I(N__77135));
    LocalMux I__18059 (
            .O(N__77422),
            .I(N__77132));
    LocalMux I__18058 (
            .O(N__77415),
            .I(N__77129));
    LocalMux I__18057 (
            .O(N__77412),
            .I(N__77126));
    LocalMux I__18056 (
            .O(N__77409),
            .I(N__77123));
    LocalMux I__18055 (
            .O(N__77406),
            .I(N__77120));
    LocalMux I__18054 (
            .O(N__77403),
            .I(N__77117));
    SRMux I__18053 (
            .O(N__77402),
            .I(N__76716));
    SRMux I__18052 (
            .O(N__77401),
            .I(N__76716));
    SRMux I__18051 (
            .O(N__77400),
            .I(N__76716));
    SRMux I__18050 (
            .O(N__77399),
            .I(N__76716));
    SRMux I__18049 (
            .O(N__77398),
            .I(N__76716));
    SRMux I__18048 (
            .O(N__77397),
            .I(N__76716));
    SRMux I__18047 (
            .O(N__77396),
            .I(N__76716));
    SRMux I__18046 (
            .O(N__77395),
            .I(N__76716));
    SRMux I__18045 (
            .O(N__77394),
            .I(N__76716));
    SRMux I__18044 (
            .O(N__77393),
            .I(N__76716));
    SRMux I__18043 (
            .O(N__77392),
            .I(N__76716));
    SRMux I__18042 (
            .O(N__77391),
            .I(N__76716));
    SRMux I__18041 (
            .O(N__77390),
            .I(N__76716));
    SRMux I__18040 (
            .O(N__77389),
            .I(N__76716));
    SRMux I__18039 (
            .O(N__77388),
            .I(N__76716));
    SRMux I__18038 (
            .O(N__77387),
            .I(N__76716));
    SRMux I__18037 (
            .O(N__77386),
            .I(N__76716));
    SRMux I__18036 (
            .O(N__77385),
            .I(N__76716));
    SRMux I__18035 (
            .O(N__77384),
            .I(N__76716));
    SRMux I__18034 (
            .O(N__77383),
            .I(N__76716));
    SRMux I__18033 (
            .O(N__77382),
            .I(N__76716));
    SRMux I__18032 (
            .O(N__77381),
            .I(N__76716));
    SRMux I__18031 (
            .O(N__77380),
            .I(N__76716));
    SRMux I__18030 (
            .O(N__77379),
            .I(N__76716));
    SRMux I__18029 (
            .O(N__77378),
            .I(N__76716));
    SRMux I__18028 (
            .O(N__77377),
            .I(N__76716));
    SRMux I__18027 (
            .O(N__77376),
            .I(N__76716));
    SRMux I__18026 (
            .O(N__77375),
            .I(N__76716));
    SRMux I__18025 (
            .O(N__77374),
            .I(N__76716));
    SRMux I__18024 (
            .O(N__77373),
            .I(N__76716));
    SRMux I__18023 (
            .O(N__77372),
            .I(N__76716));
    SRMux I__18022 (
            .O(N__77371),
            .I(N__76716));
    SRMux I__18021 (
            .O(N__77370),
            .I(N__76716));
    SRMux I__18020 (
            .O(N__77369),
            .I(N__76716));
    SRMux I__18019 (
            .O(N__77368),
            .I(N__76716));
    SRMux I__18018 (
            .O(N__77367),
            .I(N__76716));
    SRMux I__18017 (
            .O(N__77366),
            .I(N__76716));
    SRMux I__18016 (
            .O(N__77365),
            .I(N__76716));
    SRMux I__18015 (
            .O(N__77364),
            .I(N__76716));
    SRMux I__18014 (
            .O(N__77363),
            .I(N__76716));
    SRMux I__18013 (
            .O(N__77362),
            .I(N__76716));
    SRMux I__18012 (
            .O(N__77361),
            .I(N__76716));
    SRMux I__18011 (
            .O(N__77360),
            .I(N__76716));
    SRMux I__18010 (
            .O(N__77359),
            .I(N__76716));
    SRMux I__18009 (
            .O(N__77358),
            .I(N__76716));
    SRMux I__18008 (
            .O(N__77357),
            .I(N__76716));
    SRMux I__18007 (
            .O(N__77356),
            .I(N__76716));
    SRMux I__18006 (
            .O(N__77355),
            .I(N__76716));
    SRMux I__18005 (
            .O(N__77354),
            .I(N__76716));
    SRMux I__18004 (
            .O(N__77353),
            .I(N__76716));
    SRMux I__18003 (
            .O(N__77352),
            .I(N__76716));
    SRMux I__18002 (
            .O(N__77351),
            .I(N__76716));
    SRMux I__18001 (
            .O(N__77350),
            .I(N__76716));
    SRMux I__18000 (
            .O(N__77349),
            .I(N__76716));
    SRMux I__17999 (
            .O(N__77348),
            .I(N__76716));
    SRMux I__17998 (
            .O(N__77347),
            .I(N__76716));
    SRMux I__17997 (
            .O(N__77346),
            .I(N__76716));
    SRMux I__17996 (
            .O(N__77345),
            .I(N__76716));
    SRMux I__17995 (
            .O(N__77344),
            .I(N__76716));
    SRMux I__17994 (
            .O(N__77343),
            .I(N__76716));
    SRMux I__17993 (
            .O(N__77342),
            .I(N__76716));
    SRMux I__17992 (
            .O(N__77341),
            .I(N__76716));
    SRMux I__17991 (
            .O(N__77340),
            .I(N__76716));
    SRMux I__17990 (
            .O(N__77339),
            .I(N__76716));
    SRMux I__17989 (
            .O(N__77338),
            .I(N__76716));
    SRMux I__17988 (
            .O(N__77337),
            .I(N__76716));
    SRMux I__17987 (
            .O(N__77336),
            .I(N__76716));
    SRMux I__17986 (
            .O(N__77335),
            .I(N__76716));
    SRMux I__17985 (
            .O(N__77334),
            .I(N__76716));
    SRMux I__17984 (
            .O(N__77333),
            .I(N__76716));
    SRMux I__17983 (
            .O(N__77332),
            .I(N__76716));
    SRMux I__17982 (
            .O(N__77331),
            .I(N__76716));
    SRMux I__17981 (
            .O(N__77330),
            .I(N__76716));
    SRMux I__17980 (
            .O(N__77329),
            .I(N__76716));
    SRMux I__17979 (
            .O(N__77328),
            .I(N__76716));
    SRMux I__17978 (
            .O(N__77327),
            .I(N__76716));
    SRMux I__17977 (
            .O(N__77326),
            .I(N__76716));
    SRMux I__17976 (
            .O(N__77325),
            .I(N__76716));
    SRMux I__17975 (
            .O(N__77324),
            .I(N__76716));
    SRMux I__17974 (
            .O(N__77323),
            .I(N__76716));
    SRMux I__17973 (
            .O(N__77322),
            .I(N__76716));
    SRMux I__17972 (
            .O(N__77321),
            .I(N__76716));
    SRMux I__17971 (
            .O(N__77320),
            .I(N__76716));
    SRMux I__17970 (
            .O(N__77319),
            .I(N__76716));
    SRMux I__17969 (
            .O(N__77318),
            .I(N__76716));
    SRMux I__17968 (
            .O(N__77317),
            .I(N__76716));
    SRMux I__17967 (
            .O(N__77316),
            .I(N__76716));
    SRMux I__17966 (
            .O(N__77315),
            .I(N__76716));
    SRMux I__17965 (
            .O(N__77314),
            .I(N__76716));
    SRMux I__17964 (
            .O(N__77313),
            .I(N__76716));
    SRMux I__17963 (
            .O(N__77312),
            .I(N__76716));
    SRMux I__17962 (
            .O(N__77311),
            .I(N__76716));
    SRMux I__17961 (
            .O(N__77310),
            .I(N__76716));
    SRMux I__17960 (
            .O(N__77309),
            .I(N__76716));
    SRMux I__17959 (
            .O(N__77308),
            .I(N__76716));
    SRMux I__17958 (
            .O(N__77307),
            .I(N__76716));
    SRMux I__17957 (
            .O(N__77306),
            .I(N__76716));
    SRMux I__17956 (
            .O(N__77305),
            .I(N__76716));
    SRMux I__17955 (
            .O(N__77304),
            .I(N__76716));
    SRMux I__17954 (
            .O(N__77303),
            .I(N__76716));
    SRMux I__17953 (
            .O(N__77302),
            .I(N__76716));
    SRMux I__17952 (
            .O(N__77301),
            .I(N__76716));
    SRMux I__17951 (
            .O(N__77300),
            .I(N__76716));
    SRMux I__17950 (
            .O(N__77299),
            .I(N__76716));
    SRMux I__17949 (
            .O(N__77298),
            .I(N__76716));
    SRMux I__17948 (
            .O(N__77297),
            .I(N__76716));
    SRMux I__17947 (
            .O(N__77296),
            .I(N__76716));
    SRMux I__17946 (
            .O(N__77295),
            .I(N__76716));
    SRMux I__17945 (
            .O(N__77294),
            .I(N__76716));
    SRMux I__17944 (
            .O(N__77293),
            .I(N__76716));
    SRMux I__17943 (
            .O(N__77292),
            .I(N__76716));
    SRMux I__17942 (
            .O(N__77291),
            .I(N__76716));
    SRMux I__17941 (
            .O(N__77290),
            .I(N__76716));
    SRMux I__17940 (
            .O(N__77289),
            .I(N__76716));
    SRMux I__17939 (
            .O(N__77288),
            .I(N__76716));
    SRMux I__17938 (
            .O(N__77287),
            .I(N__76716));
    SRMux I__17937 (
            .O(N__77286),
            .I(N__76716));
    SRMux I__17936 (
            .O(N__77285),
            .I(N__76716));
    SRMux I__17935 (
            .O(N__77284),
            .I(N__76716));
    SRMux I__17934 (
            .O(N__77283),
            .I(N__76716));
    SRMux I__17933 (
            .O(N__77282),
            .I(N__76716));
    SRMux I__17932 (
            .O(N__77281),
            .I(N__76716));
    SRMux I__17931 (
            .O(N__77280),
            .I(N__76716));
    SRMux I__17930 (
            .O(N__77279),
            .I(N__76716));
    SRMux I__17929 (
            .O(N__77278),
            .I(N__76716));
    SRMux I__17928 (
            .O(N__77277),
            .I(N__76716));
    SRMux I__17927 (
            .O(N__77276),
            .I(N__76716));
    SRMux I__17926 (
            .O(N__77275),
            .I(N__76716));
    SRMux I__17925 (
            .O(N__77274),
            .I(N__76716));
    SRMux I__17924 (
            .O(N__77273),
            .I(N__76716));
    SRMux I__17923 (
            .O(N__77272),
            .I(N__76716));
    SRMux I__17922 (
            .O(N__77271),
            .I(N__76716));
    SRMux I__17921 (
            .O(N__77270),
            .I(N__76716));
    SRMux I__17920 (
            .O(N__77269),
            .I(N__76716));
    SRMux I__17919 (
            .O(N__77268),
            .I(N__76716));
    SRMux I__17918 (
            .O(N__77267),
            .I(N__76716));
    SRMux I__17917 (
            .O(N__77266),
            .I(N__76716));
    SRMux I__17916 (
            .O(N__77265),
            .I(N__76716));
    SRMux I__17915 (
            .O(N__77264),
            .I(N__76716));
    SRMux I__17914 (
            .O(N__77263),
            .I(N__76716));
    SRMux I__17913 (
            .O(N__77262),
            .I(N__76716));
    SRMux I__17912 (
            .O(N__77261),
            .I(N__76716));
    SRMux I__17911 (
            .O(N__77260),
            .I(N__76716));
    SRMux I__17910 (
            .O(N__77259),
            .I(N__76716));
    SRMux I__17909 (
            .O(N__77258),
            .I(N__76716));
    SRMux I__17908 (
            .O(N__77257),
            .I(N__76716));
    SRMux I__17907 (
            .O(N__77256),
            .I(N__76716));
    SRMux I__17906 (
            .O(N__77255),
            .I(N__76716));
    SRMux I__17905 (
            .O(N__77254),
            .I(N__76716));
    SRMux I__17904 (
            .O(N__77253),
            .I(N__76716));
    SRMux I__17903 (
            .O(N__77252),
            .I(N__76716));
    SRMux I__17902 (
            .O(N__77251),
            .I(N__76716));
    SRMux I__17901 (
            .O(N__77250),
            .I(N__76716));
    SRMux I__17900 (
            .O(N__77249),
            .I(N__76716));
    SRMux I__17899 (
            .O(N__77248),
            .I(N__76716));
    SRMux I__17898 (
            .O(N__77247),
            .I(N__76716));
    SRMux I__17897 (
            .O(N__77246),
            .I(N__76716));
    Glb2LocalMux I__17896 (
            .O(N__77243),
            .I(N__76716));
    Glb2LocalMux I__17895 (
            .O(N__77240),
            .I(N__76716));
    Glb2LocalMux I__17894 (
            .O(N__77237),
            .I(N__76716));
    Glb2LocalMux I__17893 (
            .O(N__77234),
            .I(N__76716));
    Glb2LocalMux I__17892 (
            .O(N__77231),
            .I(N__76716));
    Glb2LocalMux I__17891 (
            .O(N__77228),
            .I(N__76716));
    Glb2LocalMux I__17890 (
            .O(N__77225),
            .I(N__76716));
    Glb2LocalMux I__17889 (
            .O(N__77222),
            .I(N__76716));
    Glb2LocalMux I__17888 (
            .O(N__77219),
            .I(N__76716));
    Glb2LocalMux I__17887 (
            .O(N__77216),
            .I(N__76716));
    Glb2LocalMux I__17886 (
            .O(N__77213),
            .I(N__76716));
    Glb2LocalMux I__17885 (
            .O(N__77210),
            .I(N__76716));
    Glb2LocalMux I__17884 (
            .O(N__77207),
            .I(N__76716));
    Glb2LocalMux I__17883 (
            .O(N__77204),
            .I(N__76716));
    Glb2LocalMux I__17882 (
            .O(N__77201),
            .I(N__76716));
    Glb2LocalMux I__17881 (
            .O(N__77198),
            .I(N__76716));
    Glb2LocalMux I__17880 (
            .O(N__77195),
            .I(N__76716));
    Glb2LocalMux I__17879 (
            .O(N__77192),
            .I(N__76716));
    Glb2LocalMux I__17878 (
            .O(N__77189),
            .I(N__76716));
    Glb2LocalMux I__17877 (
            .O(N__77186),
            .I(N__76716));
    Glb2LocalMux I__17876 (
            .O(N__77183),
            .I(N__76716));
    Glb2LocalMux I__17875 (
            .O(N__77180),
            .I(N__76716));
    Glb2LocalMux I__17874 (
            .O(N__77177),
            .I(N__76716));
    Glb2LocalMux I__17873 (
            .O(N__77174),
            .I(N__76716));
    Glb2LocalMux I__17872 (
            .O(N__77171),
            .I(N__76716));
    Glb2LocalMux I__17871 (
            .O(N__77168),
            .I(N__76716));
    Glb2LocalMux I__17870 (
            .O(N__77165),
            .I(N__76716));
    Glb2LocalMux I__17869 (
            .O(N__77162),
            .I(N__76716));
    Glb2LocalMux I__17868 (
            .O(N__77159),
            .I(N__76716));
    Glb2LocalMux I__17867 (
            .O(N__77156),
            .I(N__76716));
    Glb2LocalMux I__17866 (
            .O(N__77153),
            .I(N__76716));
    Glb2LocalMux I__17865 (
            .O(N__77150),
            .I(N__76716));
    Glb2LocalMux I__17864 (
            .O(N__77147),
            .I(N__76716));
    Glb2LocalMux I__17863 (
            .O(N__77144),
            .I(N__76716));
    Glb2LocalMux I__17862 (
            .O(N__77141),
            .I(N__76716));
    Glb2LocalMux I__17861 (
            .O(N__77138),
            .I(N__76716));
    Glb2LocalMux I__17860 (
            .O(N__77135),
            .I(N__76716));
    Glb2LocalMux I__17859 (
            .O(N__77132),
            .I(N__76716));
    Glb2LocalMux I__17858 (
            .O(N__77129),
            .I(N__76716));
    Glb2LocalMux I__17857 (
            .O(N__77126),
            .I(N__76716));
    Glb2LocalMux I__17856 (
            .O(N__77123),
            .I(N__76716));
    Glb2LocalMux I__17855 (
            .O(N__77120),
            .I(N__76716));
    Glb2LocalMux I__17854 (
            .O(N__77117),
            .I(N__76716));
    GlobalMux I__17853 (
            .O(N__76716),
            .I(N__76713));
    gio2CtrlBuf I__17852 (
            .O(N__76713),
            .I(reset_system_g));
    IoInMux I__17851 (
            .O(N__76710),
            .I(N__76707));
    LocalMux I__17850 (
            .O(N__76707),
            .I(N__76704));
    Span4Mux_s1_v I__17849 (
            .O(N__76704),
            .I(N__76701));
    Odrv4 I__17848 (
            .O(N__76701),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__17847 (
            .O(N__76698),
            .I(N__76695));
    LocalMux I__17846 (
            .O(N__76695),
            .I(N__76690));
    InMux I__17845 (
            .O(N__76694),
            .I(N__76687));
    InMux I__17844 (
            .O(N__76693),
            .I(N__76684));
    Span4Mux_h I__17843 (
            .O(N__76690),
            .I(N__76681));
    LocalMux I__17842 (
            .O(N__76687),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__17841 (
            .O(N__76684),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv4 I__17840 (
            .O(N__76681),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__17839 (
            .O(N__76674),
            .I(N__76671));
    LocalMux I__17838 (
            .O(N__76671),
            .I(N__76667));
    InMux I__17837 (
            .O(N__76670),
            .I(N__76664));
    Span4Mux_h I__17836 (
            .O(N__76667),
            .I(N__76661));
    LocalMux I__17835 (
            .O(N__76664),
            .I(N__76658));
    Span4Mux_v I__17834 (
            .O(N__76661),
            .I(N__76654));
    Span4Mux_h I__17833 (
            .O(N__76658),
            .I(N__76651));
    InMux I__17832 (
            .O(N__76657),
            .I(N__76648));
    Odrv4 I__17831 (
            .O(N__76654),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__17830 (
            .O(N__76651),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__17829 (
            .O(N__76648),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    CascadeMux I__17828 (
            .O(N__76641),
            .I(N__76635));
    InMux I__17827 (
            .O(N__76640),
            .I(N__76601));
    InMux I__17826 (
            .O(N__76639),
            .I(N__76601));
    InMux I__17825 (
            .O(N__76638),
            .I(N__76601));
    InMux I__17824 (
            .O(N__76635),
            .I(N__76596));
    InMux I__17823 (
            .O(N__76634),
            .I(N__76596));
    InMux I__17822 (
            .O(N__76633),
            .I(N__76585));
    InMux I__17821 (
            .O(N__76632),
            .I(N__76585));
    InMux I__17820 (
            .O(N__76631),
            .I(N__76585));
    InMux I__17819 (
            .O(N__76630),
            .I(N__76585));
    InMux I__17818 (
            .O(N__76629),
            .I(N__76585));
    InMux I__17817 (
            .O(N__76628),
            .I(N__76576));
    InMux I__17816 (
            .O(N__76627),
            .I(N__76576));
    InMux I__17815 (
            .O(N__76626),
            .I(N__76576));
    InMux I__17814 (
            .O(N__76625),
            .I(N__76576));
    InMux I__17813 (
            .O(N__76624),
            .I(N__76569));
    InMux I__17812 (
            .O(N__76623),
            .I(N__76569));
    InMux I__17811 (
            .O(N__76622),
            .I(N__76569));
    InMux I__17810 (
            .O(N__76621),
            .I(N__76560));
    InMux I__17809 (
            .O(N__76620),
            .I(N__76555));
    InMux I__17808 (
            .O(N__76619),
            .I(N__76555));
    InMux I__17807 (
            .O(N__76618),
            .I(N__76548));
    InMux I__17806 (
            .O(N__76617),
            .I(N__76548));
    InMux I__17805 (
            .O(N__76616),
            .I(N__76548));
    InMux I__17804 (
            .O(N__76615),
            .I(N__76535));
    InMux I__17803 (
            .O(N__76614),
            .I(N__76535));
    InMux I__17802 (
            .O(N__76613),
            .I(N__76535));
    InMux I__17801 (
            .O(N__76612),
            .I(N__76535));
    InMux I__17800 (
            .O(N__76611),
            .I(N__76535));
    InMux I__17799 (
            .O(N__76610),
            .I(N__76535));
    CascadeMux I__17798 (
            .O(N__76609),
            .I(N__76531));
    InMux I__17797 (
            .O(N__76608),
            .I(N__76524));
    LocalMux I__17796 (
            .O(N__76601),
            .I(N__76521));
    LocalMux I__17795 (
            .O(N__76596),
            .I(N__76518));
    LocalMux I__17794 (
            .O(N__76585),
            .I(N__76511));
    LocalMux I__17793 (
            .O(N__76576),
            .I(N__76511));
    LocalMux I__17792 (
            .O(N__76569),
            .I(N__76511));
    InMux I__17791 (
            .O(N__76568),
            .I(N__76502));
    InMux I__17790 (
            .O(N__76567),
            .I(N__76502));
    InMux I__17789 (
            .O(N__76566),
            .I(N__76502));
    InMux I__17788 (
            .O(N__76565),
            .I(N__76502));
    InMux I__17787 (
            .O(N__76564),
            .I(N__76497));
    InMux I__17786 (
            .O(N__76563),
            .I(N__76497));
    LocalMux I__17785 (
            .O(N__76560),
            .I(N__76494));
    LocalMux I__17784 (
            .O(N__76555),
            .I(N__76481));
    LocalMux I__17783 (
            .O(N__76548),
            .I(N__76481));
    LocalMux I__17782 (
            .O(N__76535),
            .I(N__76481));
    InMux I__17781 (
            .O(N__76534),
            .I(N__76466));
    InMux I__17780 (
            .O(N__76531),
            .I(N__76466));
    InMux I__17779 (
            .O(N__76530),
            .I(N__76466));
    InMux I__17778 (
            .O(N__76529),
            .I(N__76466));
    CascadeMux I__17777 (
            .O(N__76528),
            .I(N__76463));
    InMux I__17776 (
            .O(N__76527),
            .I(N__76458));
    LocalMux I__17775 (
            .O(N__76524),
            .I(N__76454));
    Span4Mux_v I__17774 (
            .O(N__76521),
            .I(N__76445));
    Span4Mux_v I__17773 (
            .O(N__76518),
            .I(N__76445));
    Span4Mux_v I__17772 (
            .O(N__76511),
            .I(N__76445));
    LocalMux I__17771 (
            .O(N__76502),
            .I(N__76445));
    LocalMux I__17770 (
            .O(N__76497),
            .I(N__76440));
    Span4Mux_v I__17769 (
            .O(N__76494),
            .I(N__76440));
    InMux I__17768 (
            .O(N__76493),
            .I(N__76433));
    InMux I__17767 (
            .O(N__76492),
            .I(N__76433));
    InMux I__17766 (
            .O(N__76491),
            .I(N__76433));
    InMux I__17765 (
            .O(N__76490),
            .I(N__76426));
    InMux I__17764 (
            .O(N__76489),
            .I(N__76426));
    InMux I__17763 (
            .O(N__76488),
            .I(N__76426));
    Span4Mux_v I__17762 (
            .O(N__76481),
            .I(N__76423));
    InMux I__17761 (
            .O(N__76480),
            .I(N__76410));
    InMux I__17760 (
            .O(N__76479),
            .I(N__76410));
    InMux I__17759 (
            .O(N__76478),
            .I(N__76410));
    InMux I__17758 (
            .O(N__76477),
            .I(N__76410));
    InMux I__17757 (
            .O(N__76476),
            .I(N__76410));
    InMux I__17756 (
            .O(N__76475),
            .I(N__76410));
    LocalMux I__17755 (
            .O(N__76466),
            .I(N__76403));
    InMux I__17754 (
            .O(N__76463),
            .I(N__76395));
    InMux I__17753 (
            .O(N__76462),
            .I(N__76392));
    InMux I__17752 (
            .O(N__76461),
            .I(N__76389));
    LocalMux I__17751 (
            .O(N__76458),
            .I(N__76386));
    InMux I__17750 (
            .O(N__76457),
            .I(N__76383));
    Span4Mux_v I__17749 (
            .O(N__76454),
            .I(N__76376));
    Span4Mux_h I__17748 (
            .O(N__76445),
            .I(N__76376));
    Span4Mux_h I__17747 (
            .O(N__76440),
            .I(N__76376));
    LocalMux I__17746 (
            .O(N__76433),
            .I(N__76367));
    LocalMux I__17745 (
            .O(N__76426),
            .I(N__76367));
    Sp12to4 I__17744 (
            .O(N__76423),
            .I(N__76367));
    LocalMux I__17743 (
            .O(N__76410),
            .I(N__76367));
    InMux I__17742 (
            .O(N__76409),
            .I(N__76358));
    InMux I__17741 (
            .O(N__76408),
            .I(N__76358));
    InMux I__17740 (
            .O(N__76407),
            .I(N__76358));
    InMux I__17739 (
            .O(N__76406),
            .I(N__76358));
    Span12Mux_v I__17738 (
            .O(N__76403),
            .I(N__76355));
    InMux I__17737 (
            .O(N__76402),
            .I(N__76344));
    InMux I__17736 (
            .O(N__76401),
            .I(N__76344));
    InMux I__17735 (
            .O(N__76400),
            .I(N__76344));
    InMux I__17734 (
            .O(N__76399),
            .I(N__76344));
    InMux I__17733 (
            .O(N__76398),
            .I(N__76344));
    LocalMux I__17732 (
            .O(N__76395),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__17731 (
            .O(N__76392),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__17730 (
            .O(N__76389),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__17729 (
            .O(N__76386),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__17728 (
            .O(N__76383),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__17727 (
            .O(N__76376),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv12 I__17726 (
            .O(N__76367),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__17725 (
            .O(N__76358),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv12 I__17724 (
            .O(N__76355),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__17723 (
            .O(N__76344),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    InMux I__17722 (
            .O(N__76323),
            .I(N__76320));
    LocalMux I__17721 (
            .O(N__76320),
            .I(N__76316));
    InMux I__17720 (
            .O(N__76319),
            .I(N__76313));
    Span4Mux_v I__17719 (
            .O(N__76316),
            .I(N__76310));
    LocalMux I__17718 (
            .O(N__76313),
            .I(N__76307));
    Span4Mux_h I__17717 (
            .O(N__76310),
            .I(N__76301));
    Span4Mux_h I__17716 (
            .O(N__76307),
            .I(N__76301));
    InMux I__17715 (
            .O(N__76306),
            .I(N__76298));
    Odrv4 I__17714 (
            .O(N__76301),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__17713 (
            .O(N__76298),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    CascadeMux I__17712 (
            .O(N__76293),
            .I(N__76288));
    CascadeMux I__17711 (
            .O(N__76292),
            .I(N__76280));
    CascadeMux I__17710 (
            .O(N__76291),
            .I(N__76273));
    InMux I__17709 (
            .O(N__76288),
            .I(N__76264));
    InMux I__17708 (
            .O(N__76287),
            .I(N__76264));
    CascadeMux I__17707 (
            .O(N__76286),
            .I(N__76259));
    CascadeMux I__17706 (
            .O(N__76285),
            .I(N__76256));
    CascadeMux I__17705 (
            .O(N__76284),
            .I(N__76251));
    CascadeMux I__17704 (
            .O(N__76283),
            .I(N__76247));
    InMux I__17703 (
            .O(N__76280),
            .I(N__76242));
    InMux I__17702 (
            .O(N__76279),
            .I(N__76237));
    InMux I__17701 (
            .O(N__76278),
            .I(N__76237));
    InMux I__17700 (
            .O(N__76277),
            .I(N__76234));
    InMux I__17699 (
            .O(N__76276),
            .I(N__76227));
    InMux I__17698 (
            .O(N__76273),
            .I(N__76227));
    InMux I__17697 (
            .O(N__76272),
            .I(N__76227));
    InMux I__17696 (
            .O(N__76271),
            .I(N__76221));
    InMux I__17695 (
            .O(N__76270),
            .I(N__76214));
    InMux I__17694 (
            .O(N__76269),
            .I(N__76214));
    LocalMux I__17693 (
            .O(N__76264),
            .I(N__76211));
    InMux I__17692 (
            .O(N__76263),
            .I(N__76200));
    InMux I__17691 (
            .O(N__76262),
            .I(N__76200));
    InMux I__17690 (
            .O(N__76259),
            .I(N__76200));
    InMux I__17689 (
            .O(N__76256),
            .I(N__76200));
    InMux I__17688 (
            .O(N__76255),
            .I(N__76200));
    InMux I__17687 (
            .O(N__76254),
            .I(N__76195));
    InMux I__17686 (
            .O(N__76251),
            .I(N__76195));
    InMux I__17685 (
            .O(N__76250),
            .I(N__76188));
    InMux I__17684 (
            .O(N__76247),
            .I(N__76188));
    InMux I__17683 (
            .O(N__76246),
            .I(N__76188));
    InMux I__17682 (
            .O(N__76245),
            .I(N__76185));
    LocalMux I__17681 (
            .O(N__76242),
            .I(N__76176));
    LocalMux I__17680 (
            .O(N__76237),
            .I(N__76176));
    LocalMux I__17679 (
            .O(N__76234),
            .I(N__76176));
    LocalMux I__17678 (
            .O(N__76227),
            .I(N__76176));
    CascadeMux I__17677 (
            .O(N__76226),
            .I(N__76171));
    CascadeMux I__17676 (
            .O(N__76225),
            .I(N__76167));
    InMux I__17675 (
            .O(N__76224),
            .I(N__76163));
    LocalMux I__17674 (
            .O(N__76221),
            .I(N__76160));
    CascadeMux I__17673 (
            .O(N__76220),
            .I(N__76152));
    CascadeMux I__17672 (
            .O(N__76219),
            .I(N__76148));
    LocalMux I__17671 (
            .O(N__76214),
            .I(N__76144));
    Sp12to4 I__17670 (
            .O(N__76211),
            .I(N__76133));
    LocalMux I__17669 (
            .O(N__76200),
            .I(N__76133));
    LocalMux I__17668 (
            .O(N__76195),
            .I(N__76133));
    LocalMux I__17667 (
            .O(N__76188),
            .I(N__76133));
    LocalMux I__17666 (
            .O(N__76185),
            .I(N__76133));
    Span4Mux_v I__17665 (
            .O(N__76176),
            .I(N__76130));
    InMux I__17664 (
            .O(N__76175),
            .I(N__76125));
    InMux I__17663 (
            .O(N__76174),
            .I(N__76125));
    InMux I__17662 (
            .O(N__76171),
            .I(N__76118));
    InMux I__17661 (
            .O(N__76170),
            .I(N__76118));
    InMux I__17660 (
            .O(N__76167),
            .I(N__76118));
    InMux I__17659 (
            .O(N__76166),
            .I(N__76115));
    LocalMux I__17658 (
            .O(N__76163),
            .I(N__76110));
    Sp12to4 I__17657 (
            .O(N__76160),
            .I(N__76110));
    InMux I__17656 (
            .O(N__76159),
            .I(N__76107));
    InMux I__17655 (
            .O(N__76158),
            .I(N__76098));
    InMux I__17654 (
            .O(N__76157),
            .I(N__76098));
    InMux I__17653 (
            .O(N__76156),
            .I(N__76098));
    InMux I__17652 (
            .O(N__76155),
            .I(N__76098));
    InMux I__17651 (
            .O(N__76152),
            .I(N__76094));
    InMux I__17650 (
            .O(N__76151),
            .I(N__76091));
    InMux I__17649 (
            .O(N__76148),
            .I(N__76088));
    InMux I__17648 (
            .O(N__76147),
            .I(N__76085));
    Span4Mux_v I__17647 (
            .O(N__76144),
            .I(N__76082));
    Span12Mux_v I__17646 (
            .O(N__76133),
            .I(N__76079));
    Sp12to4 I__17645 (
            .O(N__76130),
            .I(N__76064));
    LocalMux I__17644 (
            .O(N__76125),
            .I(N__76064));
    LocalMux I__17643 (
            .O(N__76118),
            .I(N__76064));
    LocalMux I__17642 (
            .O(N__76115),
            .I(N__76064));
    Span12Mux_v I__17641 (
            .O(N__76110),
            .I(N__76064));
    LocalMux I__17640 (
            .O(N__76107),
            .I(N__76064));
    LocalMux I__17639 (
            .O(N__76098),
            .I(N__76064));
    InMux I__17638 (
            .O(N__76097),
            .I(N__76061));
    LocalMux I__17637 (
            .O(N__76094),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__17636 (
            .O(N__76091),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__17635 (
            .O(N__76088),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__17634 (
            .O(N__76085),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__17633 (
            .O(N__76082),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv12 I__17632 (
            .O(N__76079),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv12 I__17631 (
            .O(N__76064),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__17630 (
            .O(N__76061),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    InMux I__17629 (
            .O(N__76044),
            .I(N__76041));
    LocalMux I__17628 (
            .O(N__76041),
            .I(N__76038));
    Span4Mux_h I__17627 (
            .O(N__76038),
            .I(N__76035));
    Odrv4 I__17626 (
            .O(N__76035),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ));
    CascadeMux I__17625 (
            .O(N__76032),
            .I(N__76029));
    InMux I__17624 (
            .O(N__76029),
            .I(N__76026));
    LocalMux I__17623 (
            .O(N__76026),
            .I(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ));
    InMux I__17622 (
            .O(N__76023),
            .I(N__76020));
    LocalMux I__17621 (
            .O(N__76020),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__17620 (
            .O(N__76017),
            .I(N__76014));
    LocalMux I__17619 (
            .O(N__76014),
            .I(N__76011));
    Span4Mux_v I__17618 (
            .O(N__76011),
            .I(N__76008));
    Span4Mux_h I__17617 (
            .O(N__76008),
            .I(N__76005));
    Odrv4 I__17616 (
            .O(N__76005),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__17615 (
            .O(N__76002),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__17614 (
            .O(N__75999),
            .I(N__75996));
    LocalMux I__17613 (
            .O(N__75996),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ));
    CascadeMux I__17612 (
            .O(N__75993),
            .I(N__75990));
    InMux I__17611 (
            .O(N__75990),
            .I(N__75987));
    LocalMux I__17610 (
            .O(N__75987),
            .I(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ));
    InMux I__17609 (
            .O(N__75984),
            .I(N__75981));
    LocalMux I__17608 (
            .O(N__75981),
            .I(N__75978));
    Span4Mux_v I__17607 (
            .O(N__75978),
            .I(N__75975));
    Odrv4 I__17606 (
            .O(N__75975),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__17605 (
            .O(N__75972),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__17604 (
            .O(N__75969),
            .I(N__75966));
    LocalMux I__17603 (
            .O(N__75966),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__17602 (
            .O(N__75963),
            .I(N__75960));
    LocalMux I__17601 (
            .O(N__75960),
            .I(N__75957));
    Span4Mux_v I__17600 (
            .O(N__75957),
            .I(N__75954));
    Odrv4 I__17599 (
            .O(N__75954),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__17598 (
            .O(N__75951),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__17597 (
            .O(N__75948),
            .I(N__75945));
    LocalMux I__17596 (
            .O(N__75945),
            .I(N__75942));
    Odrv4 I__17595 (
            .O(N__75942),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__17594 (
            .O(N__75939),
            .I(N__75936));
    LocalMux I__17593 (
            .O(N__75936),
            .I(\pid_side.N_1881_i ));
    CascadeMux I__17592 (
            .O(N__75933),
            .I(\pid_side.N_1881_i_cascade_ ));
    InMux I__17591 (
            .O(N__75930),
            .I(N__75927));
    LocalMux I__17590 (
            .O(N__75927),
            .I(N__75923));
    InMux I__17589 (
            .O(N__75926),
            .I(N__75920));
    Span4Mux_h I__17588 (
            .O(N__75923),
            .I(N__75915));
    LocalMux I__17587 (
            .O(N__75920),
            .I(N__75915));
    Odrv4 I__17586 (
            .O(N__75915),
            .I(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ));
    InMux I__17585 (
            .O(N__75912),
            .I(N__75906));
    InMux I__17584 (
            .O(N__75911),
            .I(N__75906));
    LocalMux I__17583 (
            .O(N__75906),
            .I(N__75903));
    Odrv4 I__17582 (
            .O(N__75903),
            .I(\pid_side.N_1887_i ));
    InMux I__17581 (
            .O(N__75900),
            .I(N__75897));
    LocalMux I__17580 (
            .O(N__75897),
            .I(N__75894));
    Span4Mux_h I__17579 (
            .O(N__75894),
            .I(N__75890));
    InMux I__17578 (
            .O(N__75893),
            .I(N__75887));
    Span4Mux_h I__17577 (
            .O(N__75890),
            .I(N__75884));
    LocalMux I__17576 (
            .O(N__75887),
            .I(N__75881));
    Odrv4 I__17575 (
            .O(N__75884),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ));
    Odrv12 I__17574 (
            .O(N__75881),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ));
    InMux I__17573 (
            .O(N__75876),
            .I(N__75873));
    LocalMux I__17572 (
            .O(N__75873),
            .I(N__75870));
    Span4Mux_v I__17571 (
            .O(N__75870),
            .I(N__75867));
    Span4Mux_h I__17570 (
            .O(N__75867),
            .I(N__75864));
    Odrv4 I__17569 (
            .O(N__75864),
            .I(\pid_front.O_6 ));
    InMux I__17568 (
            .O(N__75861),
            .I(N__75852));
    InMux I__17567 (
            .O(N__75860),
            .I(N__75852));
    InMux I__17566 (
            .O(N__75859),
            .I(N__75852));
    LocalMux I__17565 (
            .O(N__75852),
            .I(N__75849));
    Span12Mux_h I__17564 (
            .O(N__75849),
            .I(N__75846));
    Odrv12 I__17563 (
            .O(N__75846),
            .I(\pid_front.error_d_regZ0Z_4 ));
    InMux I__17562 (
            .O(N__75843),
            .I(N__75840));
    LocalMux I__17561 (
            .O(N__75840),
            .I(N__75837));
    Span4Mux_v I__17560 (
            .O(N__75837),
            .I(N__75834));
    Span4Mux_h I__17559 (
            .O(N__75834),
            .I(N__75831));
    Odrv4 I__17558 (
            .O(N__75831),
            .I(\pid_front.O_4 ));
    InMux I__17557 (
            .O(N__75828),
            .I(N__75819));
    InMux I__17556 (
            .O(N__75827),
            .I(N__75819));
    InMux I__17555 (
            .O(N__75826),
            .I(N__75819));
    LocalMux I__17554 (
            .O(N__75819),
            .I(N__75816));
    Span4Mux_h I__17553 (
            .O(N__75816),
            .I(N__75813));
    Span4Mux_h I__17552 (
            .O(N__75813),
            .I(N__75810));
    Odrv4 I__17551 (
            .O(N__75810),
            .I(\pid_front.error_d_regZ0Z_2 ));
    InMux I__17550 (
            .O(N__75807),
            .I(N__75804));
    LocalMux I__17549 (
            .O(N__75804),
            .I(N__75801));
    Span4Mux_v I__17548 (
            .O(N__75801),
            .I(N__75798));
    Span4Mux_h I__17547 (
            .O(N__75798),
            .I(N__75795));
    Odrv4 I__17546 (
            .O(N__75795),
            .I(\pid_front.O_11 ));
    InMux I__17545 (
            .O(N__75792),
            .I(N__75785));
    InMux I__17544 (
            .O(N__75791),
            .I(N__75785));
    InMux I__17543 (
            .O(N__75790),
            .I(N__75780));
    LocalMux I__17542 (
            .O(N__75785),
            .I(N__75777));
    InMux I__17541 (
            .O(N__75784),
            .I(N__75772));
    InMux I__17540 (
            .O(N__75783),
            .I(N__75772));
    LocalMux I__17539 (
            .O(N__75780),
            .I(N__75769));
    Span4Mux_v I__17538 (
            .O(N__75777),
            .I(N__75764));
    LocalMux I__17537 (
            .O(N__75772),
            .I(N__75764));
    Span4Mux_h I__17536 (
            .O(N__75769),
            .I(N__75761));
    Span4Mux_h I__17535 (
            .O(N__75764),
            .I(N__75758));
    Span4Mux_h I__17534 (
            .O(N__75761),
            .I(N__75755));
    Span4Mux_h I__17533 (
            .O(N__75758),
            .I(N__75752));
    Odrv4 I__17532 (
            .O(N__75755),
            .I(\pid_front.error_d_regZ0Z_9 ));
    Odrv4 I__17531 (
            .O(N__75752),
            .I(\pid_front.error_d_regZ0Z_9 ));
    InMux I__17530 (
            .O(N__75747),
            .I(N__75744));
    LocalMux I__17529 (
            .O(N__75744),
            .I(N__75741));
    Span4Mux_h I__17528 (
            .O(N__75741),
            .I(N__75738));
    Span4Mux_h I__17527 (
            .O(N__75738),
            .I(N__75735));
    Odrv4 I__17526 (
            .O(N__75735),
            .I(\pid_front.O_13 ));
    InMux I__17525 (
            .O(N__75732),
            .I(N__75727));
    InMux I__17524 (
            .O(N__75731),
            .I(N__75722));
    InMux I__17523 (
            .O(N__75730),
            .I(N__75722));
    LocalMux I__17522 (
            .O(N__75727),
            .I(N__75719));
    LocalMux I__17521 (
            .O(N__75722),
            .I(N__75716));
    Span4Mux_v I__17520 (
            .O(N__75719),
            .I(N__75711));
    Span4Mux_h I__17519 (
            .O(N__75716),
            .I(N__75711));
    Span4Mux_h I__17518 (
            .O(N__75711),
            .I(N__75708));
    Span4Mux_h I__17517 (
            .O(N__75708),
            .I(N__75705));
    Odrv4 I__17516 (
            .O(N__75705),
            .I(\pid_front.error_d_regZ0Z_11 ));
    InMux I__17515 (
            .O(N__75702),
            .I(N__75699));
    LocalMux I__17514 (
            .O(N__75699),
            .I(N__75696));
    Span4Mux_v I__17513 (
            .O(N__75696),
            .I(N__75693));
    Span4Mux_h I__17512 (
            .O(N__75693),
            .I(N__75690));
    Odrv4 I__17511 (
            .O(N__75690),
            .I(\pid_front.O_5 ));
    InMux I__17510 (
            .O(N__75687),
            .I(N__75678));
    InMux I__17509 (
            .O(N__75686),
            .I(N__75678));
    InMux I__17508 (
            .O(N__75685),
            .I(N__75678));
    LocalMux I__17507 (
            .O(N__75678),
            .I(N__75675));
    Span4Mux_h I__17506 (
            .O(N__75675),
            .I(N__75672));
    Sp12to4 I__17505 (
            .O(N__75672),
            .I(N__75669));
    Span12Mux_v I__17504 (
            .O(N__75669),
            .I(N__75666));
    Odrv12 I__17503 (
            .O(N__75666),
            .I(\pid_front.error_d_regZ0Z_3 ));
    CascadeMux I__17502 (
            .O(N__75663),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2_cascade_ ));
    InMux I__17501 (
            .O(N__75660),
            .I(N__75656));
    InMux I__17500 (
            .O(N__75659),
            .I(N__75653));
    LocalMux I__17499 (
            .O(N__75656),
            .I(N__75648));
    LocalMux I__17498 (
            .O(N__75653),
            .I(N__75648));
    Span4Mux_h I__17497 (
            .O(N__75648),
            .I(N__75645));
    Odrv4 I__17496 (
            .O(N__75645),
            .I(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ));
    InMux I__17495 (
            .O(N__75642),
            .I(N__75636));
    InMux I__17494 (
            .O(N__75641),
            .I(N__75636));
    LocalMux I__17493 (
            .O(N__75636),
            .I(N__75631));
    InMux I__17492 (
            .O(N__75635),
            .I(N__75626));
    InMux I__17491 (
            .O(N__75634),
            .I(N__75626));
    Odrv4 I__17490 (
            .O(N__75631),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    LocalMux I__17489 (
            .O(N__75626),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    InMux I__17488 (
            .O(N__75621),
            .I(N__75615));
    InMux I__17487 (
            .O(N__75620),
            .I(N__75608));
    InMux I__17486 (
            .O(N__75619),
            .I(N__75608));
    InMux I__17485 (
            .O(N__75618),
            .I(N__75608));
    LocalMux I__17484 (
            .O(N__75615),
            .I(N__75603));
    LocalMux I__17483 (
            .O(N__75608),
            .I(N__75603));
    Odrv4 I__17482 (
            .O(N__75603),
            .I(\pid_side.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__17481 (
            .O(N__75600),
            .I(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ));
    InMux I__17480 (
            .O(N__75597),
            .I(N__75594));
    LocalMux I__17479 (
            .O(N__75594),
            .I(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ));
    InMux I__17478 (
            .O(N__75591),
            .I(N__75585));
    InMux I__17477 (
            .O(N__75590),
            .I(N__75585));
    LocalMux I__17476 (
            .O(N__75585),
            .I(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ));
    InMux I__17475 (
            .O(N__75582),
            .I(N__75579));
    LocalMux I__17474 (
            .O(N__75579),
            .I(N__75575));
    CascadeMux I__17473 (
            .O(N__75578),
            .I(N__75572));
    Span4Mux_v I__17472 (
            .O(N__75575),
            .I(N__75569));
    InMux I__17471 (
            .O(N__75572),
            .I(N__75566));
    Odrv4 I__17470 (
            .O(N__75569),
            .I(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ));
    LocalMux I__17469 (
            .O(N__75566),
            .I(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ));
    CascadeMux I__17468 (
            .O(N__75561),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ));
    InMux I__17467 (
            .O(N__75558),
            .I(N__75555));
    LocalMux I__17466 (
            .O(N__75555),
            .I(N__75552));
    Span4Mux_h I__17465 (
            .O(N__75552),
            .I(N__75549));
    Odrv4 I__17464 (
            .O(N__75549),
            .I(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ));
    InMux I__17463 (
            .O(N__75546),
            .I(N__75539));
    InMux I__17462 (
            .O(N__75545),
            .I(N__75539));
    InMux I__17461 (
            .O(N__75544),
            .I(N__75536));
    LocalMux I__17460 (
            .O(N__75539),
            .I(N__75533));
    LocalMux I__17459 (
            .O(N__75536),
            .I(N__75530));
    Span12Mux_s10_h I__17458 (
            .O(N__75533),
            .I(N__75527));
    Odrv4 I__17457 (
            .O(N__75530),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ));
    Odrv12 I__17456 (
            .O(N__75527),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ));
    InMux I__17455 (
            .O(N__75522),
            .I(N__75519));
    LocalMux I__17454 (
            .O(N__75519),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ));
    CascadeMux I__17453 (
            .O(N__75516),
            .I(N__75513));
    InMux I__17452 (
            .O(N__75513),
            .I(N__75509));
    InMux I__17451 (
            .O(N__75512),
            .I(N__75506));
    LocalMux I__17450 (
            .O(N__75509),
            .I(N__75503));
    LocalMux I__17449 (
            .O(N__75506),
            .I(N__75498));
    Span4Mux_h I__17448 (
            .O(N__75503),
            .I(N__75498));
    Odrv4 I__17447 (
            .O(N__75498),
            .I(\pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ));
    CascadeMux I__17446 (
            .O(N__75495),
            .I(N__75492));
    InMux I__17445 (
            .O(N__75492),
            .I(N__75486));
    InMux I__17444 (
            .O(N__75491),
            .I(N__75486));
    LocalMux I__17443 (
            .O(N__75486),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ));
    InMux I__17442 (
            .O(N__75483),
            .I(N__75480));
    LocalMux I__17441 (
            .O(N__75480),
            .I(N__75477));
    Odrv4 I__17440 (
            .O(N__75477),
            .I(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ));
    CascadeMux I__17439 (
            .O(N__75474),
            .I(N__75470));
    InMux I__17438 (
            .O(N__75473),
            .I(N__75461));
    InMux I__17437 (
            .O(N__75470),
            .I(N__75461));
    InMux I__17436 (
            .O(N__75469),
            .I(N__75461));
    InMux I__17435 (
            .O(N__75468),
            .I(N__75458));
    LocalMux I__17434 (
            .O(N__75461),
            .I(N__75455));
    LocalMux I__17433 (
            .O(N__75458),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    Odrv4 I__17432 (
            .O(N__75455),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    InMux I__17431 (
            .O(N__75450),
            .I(N__75438));
    InMux I__17430 (
            .O(N__75449),
            .I(N__75438));
    InMux I__17429 (
            .O(N__75448),
            .I(N__75438));
    InMux I__17428 (
            .O(N__75447),
            .I(N__75438));
    LocalMux I__17427 (
            .O(N__75438),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    CascadeMux I__17426 (
            .O(N__75435),
            .I(\pid_side.N_1893_i_cascade_ ));
    InMux I__17425 (
            .O(N__75432),
            .I(N__75429));
    LocalMux I__17424 (
            .O(N__75429),
            .I(N__75426));
    Span4Mux_h I__17423 (
            .O(N__75426),
            .I(N__75423));
    Span4Mux_h I__17422 (
            .O(N__75423),
            .I(N__75420));
    Odrv4 I__17421 (
            .O(N__75420),
            .I(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ));
    CascadeMux I__17420 (
            .O(N__75417),
            .I(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ));
    InMux I__17419 (
            .O(N__75414),
            .I(N__75411));
    LocalMux I__17418 (
            .O(N__75411),
            .I(N__75406));
    InMux I__17417 (
            .O(N__75410),
            .I(N__75403));
    InMux I__17416 (
            .O(N__75409),
            .I(N__75400));
    Span4Mux_h I__17415 (
            .O(N__75406),
            .I(N__75397));
    LocalMux I__17414 (
            .O(N__75403),
            .I(N__75394));
    LocalMux I__17413 (
            .O(N__75400),
            .I(N__75389));
    Span4Mux_h I__17412 (
            .O(N__75397),
            .I(N__75389));
    Odrv4 I__17411 (
            .O(N__75394),
            .I(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ));
    Odrv4 I__17410 (
            .O(N__75389),
            .I(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ));
    InMux I__17409 (
            .O(N__75384),
            .I(N__75381));
    LocalMux I__17408 (
            .O(N__75381),
            .I(N__75378));
    Span4Mux_h I__17407 (
            .O(N__75378),
            .I(N__75375));
    Odrv4 I__17406 (
            .O(N__75375),
            .I(\pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ));
    CascadeMux I__17405 (
            .O(N__75372),
            .I(N__75369));
    InMux I__17404 (
            .O(N__75369),
            .I(N__75365));
    CascadeMux I__17403 (
            .O(N__75368),
            .I(N__75361));
    LocalMux I__17402 (
            .O(N__75365),
            .I(N__75358));
    InMux I__17401 (
            .O(N__75364),
            .I(N__75355));
    InMux I__17400 (
            .O(N__75361),
            .I(N__75352));
    Span4Mux_v I__17399 (
            .O(N__75358),
            .I(N__75349));
    LocalMux I__17398 (
            .O(N__75355),
            .I(N__75346));
    LocalMux I__17397 (
            .O(N__75352),
            .I(N__75343));
    Span4Mux_h I__17396 (
            .O(N__75349),
            .I(N__75340));
    Span4Mux_h I__17395 (
            .O(N__75346),
            .I(N__75335));
    Span4Mux_v I__17394 (
            .O(N__75343),
            .I(N__75335));
    Odrv4 I__17393 (
            .O(N__75340),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    Odrv4 I__17392 (
            .O(N__75335),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    InMux I__17391 (
            .O(N__75330),
            .I(N__75327));
    LocalMux I__17390 (
            .O(N__75327),
            .I(N__75324));
    Span4Mux_h I__17389 (
            .O(N__75324),
            .I(N__75321));
    Odrv4 I__17388 (
            .O(N__75321),
            .I(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ));
    InMux I__17387 (
            .O(N__75318),
            .I(N__75315));
    LocalMux I__17386 (
            .O(N__75315),
            .I(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ));
    InMux I__17385 (
            .O(N__75312),
            .I(N__75309));
    LocalMux I__17384 (
            .O(N__75309),
            .I(N__75305));
    InMux I__17383 (
            .O(N__75308),
            .I(N__75302));
    Span4Mux_h I__17382 (
            .O(N__75305),
            .I(N__75299));
    LocalMux I__17381 (
            .O(N__75302),
            .I(N__75296));
    Odrv4 I__17380 (
            .O(N__75299),
            .I(\pid_side.error_p_regZ0Z_2 ));
    Odrv12 I__17379 (
            .O(N__75296),
            .I(\pid_side.error_p_regZ0Z_2 ));
    InMux I__17378 (
            .O(N__75291),
            .I(N__75288));
    LocalMux I__17377 (
            .O(N__75288),
            .I(N__75284));
    InMux I__17376 (
            .O(N__75287),
            .I(N__75281));
    Span4Mux_h I__17375 (
            .O(N__75284),
            .I(N__75278));
    LocalMux I__17374 (
            .O(N__75281),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    Odrv4 I__17373 (
            .O(N__75278),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    InMux I__17372 (
            .O(N__75273),
            .I(N__75270));
    LocalMux I__17371 (
            .O(N__75270),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    CascadeMux I__17370 (
            .O(N__75267),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ));
    InMux I__17369 (
            .O(N__75264),
            .I(N__75261));
    LocalMux I__17368 (
            .O(N__75261),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ));
    InMux I__17367 (
            .O(N__75258),
            .I(N__75255));
    LocalMux I__17366 (
            .O(N__75255),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ));
    CascadeMux I__17365 (
            .O(N__75252),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ));
    InMux I__17364 (
            .O(N__75249),
            .I(N__75242));
    InMux I__17363 (
            .O(N__75248),
            .I(N__75242));
    InMux I__17362 (
            .O(N__75247),
            .I(N__75239));
    LocalMux I__17361 (
            .O(N__75242),
            .I(N__75236));
    LocalMux I__17360 (
            .O(N__75239),
            .I(N__75233));
    Span4Mux_h I__17359 (
            .O(N__75236),
            .I(N__75230));
    Span4Mux_v I__17358 (
            .O(N__75233),
            .I(N__75227));
    Span4Mux_h I__17357 (
            .O(N__75230),
            .I(N__75224));
    Odrv4 I__17356 (
            .O(N__75227),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ));
    Odrv4 I__17355 (
            .O(N__75224),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ));
    CascadeMux I__17354 (
            .O(N__75219),
            .I(N__75216));
    InMux I__17353 (
            .O(N__75216),
            .I(N__75213));
    LocalMux I__17352 (
            .O(N__75213),
            .I(N__75210));
    Odrv4 I__17351 (
            .O(N__75210),
            .I(\pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ));
    CascadeMux I__17350 (
            .O(N__75207),
            .I(N__75203));
    InMux I__17349 (
            .O(N__75206),
            .I(N__75195));
    InMux I__17348 (
            .O(N__75203),
            .I(N__75195));
    InMux I__17347 (
            .O(N__75202),
            .I(N__75195));
    LocalMux I__17346 (
            .O(N__75195),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    InMux I__17345 (
            .O(N__75192),
            .I(N__75189));
    LocalMux I__17344 (
            .O(N__75189),
            .I(N__75186));
    Span4Mux_h I__17343 (
            .O(N__75186),
            .I(N__75183));
    Odrv4 I__17342 (
            .O(N__75183),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ));
    CascadeMux I__17341 (
            .O(N__75180),
            .I(N__75177));
    InMux I__17340 (
            .O(N__75177),
            .I(N__75173));
    InMux I__17339 (
            .O(N__75176),
            .I(N__75170));
    LocalMux I__17338 (
            .O(N__75173),
            .I(N__75167));
    LocalMux I__17337 (
            .O(N__75170),
            .I(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ));
    Odrv12 I__17336 (
            .O(N__75167),
            .I(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ));
    CascadeMux I__17335 (
            .O(N__75162),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ));
    InMux I__17334 (
            .O(N__75159),
            .I(N__75154));
    InMux I__17333 (
            .O(N__75158),
            .I(N__75151));
    InMux I__17332 (
            .O(N__75157),
            .I(N__75148));
    LocalMux I__17331 (
            .O(N__75154),
            .I(N__75145));
    LocalMux I__17330 (
            .O(N__75151),
            .I(N__75142));
    LocalMux I__17329 (
            .O(N__75148),
            .I(N__75139));
    Span4Mux_v I__17328 (
            .O(N__75145),
            .I(N__75134));
    Span4Mux_h I__17327 (
            .O(N__75142),
            .I(N__75134));
    Span4Mux_v I__17326 (
            .O(N__75139),
            .I(N__75129));
    Span4Mux_h I__17325 (
            .O(N__75134),
            .I(N__75129));
    Odrv4 I__17324 (
            .O(N__75129),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ));
    InMux I__17323 (
            .O(N__75126),
            .I(N__75123));
    LocalMux I__17322 (
            .O(N__75123),
            .I(N__75120));
    Odrv4 I__17321 (
            .O(N__75120),
            .I(\pid_side.error_p_reg_esr_RNIT9E37Z0Z_7 ));
    InMux I__17320 (
            .O(N__75117),
            .I(N__75114));
    LocalMux I__17319 (
            .O(N__75114),
            .I(N__75111));
    Odrv4 I__17318 (
            .O(N__75111),
            .I(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10 ));
    CascadeMux I__17317 (
            .O(N__75108),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ));
    CascadeMux I__17316 (
            .O(N__75105),
            .I(N__75102));
    InMux I__17315 (
            .O(N__75102),
            .I(N__75099));
    LocalMux I__17314 (
            .O(N__75099),
            .I(N__75096));
    Odrv4 I__17313 (
            .O(N__75096),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ));
    InMux I__17312 (
            .O(N__75093),
            .I(N__75090));
    LocalMux I__17311 (
            .O(N__75090),
            .I(N__75087));
    Odrv4 I__17310 (
            .O(N__75087),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ));
    CascadeMux I__17309 (
            .O(N__75084),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ));
    InMux I__17308 (
            .O(N__75081),
            .I(N__75077));
    InMux I__17307 (
            .O(N__75080),
            .I(N__75073));
    LocalMux I__17306 (
            .O(N__75077),
            .I(N__75070));
    InMux I__17305 (
            .O(N__75076),
            .I(N__75067));
    LocalMux I__17304 (
            .O(N__75073),
            .I(N__75062));
    Span4Mux_h I__17303 (
            .O(N__75070),
            .I(N__75062));
    LocalMux I__17302 (
            .O(N__75067),
            .I(N__75059));
    Span4Mux_h I__17301 (
            .O(N__75062),
            .I(N__75056));
    Odrv4 I__17300 (
            .O(N__75059),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    Odrv4 I__17299 (
            .O(N__75056),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    InMux I__17298 (
            .O(N__75051),
            .I(N__75048));
    LocalMux I__17297 (
            .O(N__75048),
            .I(N__75044));
    InMux I__17296 (
            .O(N__75047),
            .I(N__75041));
    Odrv4 I__17295 (
            .O(N__75044),
            .I(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ));
    LocalMux I__17294 (
            .O(N__75041),
            .I(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ));
    CascadeMux I__17293 (
            .O(N__75036),
            .I(\pid_side.un1_pid_prereg_66_0_cascade_ ));
    InMux I__17292 (
            .O(N__75033),
            .I(N__75030));
    LocalMux I__17291 (
            .O(N__75030),
            .I(N__75027));
    Odrv4 I__17290 (
            .O(N__75027),
            .I(\pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ));
    InMux I__17289 (
            .O(N__75024),
            .I(N__75021));
    LocalMux I__17288 (
            .O(N__75021),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ));
    InMux I__17287 (
            .O(N__75018),
            .I(N__75012));
    InMux I__17286 (
            .O(N__75017),
            .I(N__75012));
    LocalMux I__17285 (
            .O(N__75012),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ));
    CascadeMux I__17284 (
            .O(N__75009),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ));
    InMux I__17283 (
            .O(N__75006),
            .I(N__74997));
    InMux I__17282 (
            .O(N__75005),
            .I(N__74997));
    InMux I__17281 (
            .O(N__75004),
            .I(N__74997));
    LocalMux I__17280 (
            .O(N__74997),
            .I(N__74993));
    InMux I__17279 (
            .O(N__74996),
            .I(N__74990));
    Span4Mux_h I__17278 (
            .O(N__74993),
            .I(N__74987));
    LocalMux I__17277 (
            .O(N__74990),
            .I(N__74984));
    Span4Mux_h I__17276 (
            .O(N__74987),
            .I(N__74981));
    Odrv4 I__17275 (
            .O(N__74984),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ));
    Odrv4 I__17274 (
            .O(N__74981),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ));
    CascadeMux I__17273 (
            .O(N__74976),
            .I(N__74973));
    InMux I__17272 (
            .O(N__74973),
            .I(N__74969));
    InMux I__17271 (
            .O(N__74972),
            .I(N__74966));
    LocalMux I__17270 (
            .O(N__74969),
            .I(N__74963));
    LocalMux I__17269 (
            .O(N__74966),
            .I(N__74960));
    Odrv12 I__17268 (
            .O(N__74963),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ));
    Odrv4 I__17267 (
            .O(N__74960),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ));
    InMux I__17266 (
            .O(N__74955),
            .I(N__74952));
    LocalMux I__17265 (
            .O(N__74952),
            .I(\pid_side.N_1869_i ));
    CascadeMux I__17264 (
            .O(N__74949),
            .I(\pid_side.N_1869_i_cascade_ ));
    InMux I__17263 (
            .O(N__74946),
            .I(N__74943));
    LocalMux I__17262 (
            .O(N__74943),
            .I(N__74940));
    Span4Mux_h I__17261 (
            .O(N__74940),
            .I(N__74937));
    Odrv4 I__17260 (
            .O(N__74937),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__17259 (
            .O(N__74934),
            .I(N__74930));
    InMux I__17258 (
            .O(N__74933),
            .I(N__74927));
    LocalMux I__17257 (
            .O(N__74930),
            .I(N__74924));
    LocalMux I__17256 (
            .O(N__74927),
            .I(N__74921));
    Span4Mux_v I__17255 (
            .O(N__74924),
            .I(N__74918));
    Span4Mux_v I__17254 (
            .O(N__74921),
            .I(N__74915));
    Span4Mux_h I__17253 (
            .O(N__74918),
            .I(N__74912));
    Span4Mux_h I__17252 (
            .O(N__74915),
            .I(N__74909));
    Odrv4 I__17251 (
            .O(N__74912),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    Odrv4 I__17250 (
            .O(N__74909),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    InMux I__17249 (
            .O(N__74904),
            .I(N__74900));
    InMux I__17248 (
            .O(N__74903),
            .I(N__74895));
    LocalMux I__17247 (
            .O(N__74900),
            .I(N__74891));
    InMux I__17246 (
            .O(N__74899),
            .I(N__74886));
    InMux I__17245 (
            .O(N__74898),
            .I(N__74886));
    LocalMux I__17244 (
            .O(N__74895),
            .I(N__74883));
    CascadeMux I__17243 (
            .O(N__74894),
            .I(N__74880));
    Span4Mux_h I__17242 (
            .O(N__74891),
            .I(N__74874));
    LocalMux I__17241 (
            .O(N__74886),
            .I(N__74874));
    Span4Mux_h I__17240 (
            .O(N__74883),
            .I(N__74870));
    InMux I__17239 (
            .O(N__74880),
            .I(N__74865));
    InMux I__17238 (
            .O(N__74879),
            .I(N__74865));
    Span4Mux_v I__17237 (
            .O(N__74874),
            .I(N__74862));
    InMux I__17236 (
            .O(N__74873),
            .I(N__74859));
    Span4Mux_h I__17235 (
            .O(N__74870),
            .I(N__74849));
    LocalMux I__17234 (
            .O(N__74865),
            .I(N__74846));
    Span4Mux_h I__17233 (
            .O(N__74862),
            .I(N__74841));
    LocalMux I__17232 (
            .O(N__74859),
            .I(N__74841));
    InMux I__17231 (
            .O(N__74858),
            .I(N__74836));
    InMux I__17230 (
            .O(N__74857),
            .I(N__74836));
    InMux I__17229 (
            .O(N__74856),
            .I(N__74831));
    InMux I__17228 (
            .O(N__74855),
            .I(N__74831));
    InMux I__17227 (
            .O(N__74854),
            .I(N__74828));
    InMux I__17226 (
            .O(N__74853),
            .I(N__74823));
    InMux I__17225 (
            .O(N__74852),
            .I(N__74823));
    Odrv4 I__17224 (
            .O(N__74849),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv12 I__17223 (
            .O(N__74846),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__17222 (
            .O(N__74841),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__17221 (
            .O(N__74836),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__17220 (
            .O(N__74831),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__17219 (
            .O(N__74828),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__17218 (
            .O(N__74823),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    CascadeMux I__17217 (
            .O(N__74808),
            .I(N__74804));
    InMux I__17216 (
            .O(N__74807),
            .I(N__74796));
    InMux I__17215 (
            .O(N__74804),
            .I(N__74796));
    InMux I__17214 (
            .O(N__74803),
            .I(N__74796));
    LocalMux I__17213 (
            .O(N__74796),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    CascadeMux I__17212 (
            .O(N__74793),
            .I(N__74790));
    InMux I__17211 (
            .O(N__74790),
            .I(N__74782));
    CascadeMux I__17210 (
            .O(N__74789),
            .I(N__74779));
    InMux I__17209 (
            .O(N__74788),
            .I(N__74776));
    InMux I__17208 (
            .O(N__74787),
            .I(N__74771));
    InMux I__17207 (
            .O(N__74786),
            .I(N__74771));
    CascadeMux I__17206 (
            .O(N__74785),
            .I(N__74767));
    LocalMux I__17205 (
            .O(N__74782),
            .I(N__74763));
    InMux I__17204 (
            .O(N__74779),
            .I(N__74760));
    LocalMux I__17203 (
            .O(N__74776),
            .I(N__74754));
    LocalMux I__17202 (
            .O(N__74771),
            .I(N__74754));
    InMux I__17201 (
            .O(N__74770),
            .I(N__74749));
    InMux I__17200 (
            .O(N__74767),
            .I(N__74749));
    CascadeMux I__17199 (
            .O(N__74766),
            .I(N__74745));
    Span4Mux_v I__17198 (
            .O(N__74763),
            .I(N__74739));
    LocalMux I__17197 (
            .O(N__74760),
            .I(N__74736));
    InMux I__17196 (
            .O(N__74759),
            .I(N__74733));
    Span4Mux_v I__17195 (
            .O(N__74754),
            .I(N__74727));
    LocalMux I__17194 (
            .O(N__74749),
            .I(N__74727));
    InMux I__17193 (
            .O(N__74748),
            .I(N__74724));
    InMux I__17192 (
            .O(N__74745),
            .I(N__74721));
    CascadeMux I__17191 (
            .O(N__74744),
            .I(N__74718));
    CascadeMux I__17190 (
            .O(N__74743),
            .I(N__74715));
    CascadeMux I__17189 (
            .O(N__74742),
            .I(N__74711));
    Span4Mux_h I__17188 (
            .O(N__74739),
            .I(N__74706));
    Span4Mux_v I__17187 (
            .O(N__74736),
            .I(N__74706));
    LocalMux I__17186 (
            .O(N__74733),
            .I(N__74703));
    InMux I__17185 (
            .O(N__74732),
            .I(N__74697));
    Span4Mux_h I__17184 (
            .O(N__74727),
            .I(N__74694));
    LocalMux I__17183 (
            .O(N__74724),
            .I(N__74689));
    LocalMux I__17182 (
            .O(N__74721),
            .I(N__74689));
    InMux I__17181 (
            .O(N__74718),
            .I(N__74684));
    InMux I__17180 (
            .O(N__74715),
            .I(N__74684));
    InMux I__17179 (
            .O(N__74714),
            .I(N__74679));
    InMux I__17178 (
            .O(N__74711),
            .I(N__74679));
    Span4Mux_h I__17177 (
            .O(N__74706),
            .I(N__74674));
    Span4Mux_h I__17176 (
            .O(N__74703),
            .I(N__74674));
    InMux I__17175 (
            .O(N__74702),
            .I(N__74667));
    InMux I__17174 (
            .O(N__74701),
            .I(N__74667));
    InMux I__17173 (
            .O(N__74700),
            .I(N__74667));
    LocalMux I__17172 (
            .O(N__74697),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__17171 (
            .O(N__74694),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__17170 (
            .O(N__74689),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__17169 (
            .O(N__74684),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__17168 (
            .O(N__74679),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__17167 (
            .O(N__74674),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__17166 (
            .O(N__74667),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__17165 (
            .O(N__74652),
            .I(N__74649));
    LocalMux I__17164 (
            .O(N__74649),
            .I(N__74646));
    Span4Mux_v I__17163 (
            .O(N__74646),
            .I(N__74642));
    InMux I__17162 (
            .O(N__74645),
            .I(N__74639));
    Span4Mux_h I__17161 (
            .O(N__74642),
            .I(N__74634));
    LocalMux I__17160 (
            .O(N__74639),
            .I(N__74634));
    Span4Mux_h I__17159 (
            .O(N__74634),
            .I(N__74631));
    Span4Mux_h I__17158 (
            .O(N__74631),
            .I(N__74628));
    Odrv4 I__17157 (
            .O(N__74628),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__17156 (
            .O(N__74625),
            .I(N__74622));
    LocalMux I__17155 (
            .O(N__74622),
            .I(N__74619));
    Span4Mux_h I__17154 (
            .O(N__74619),
            .I(N__74616));
    Odrv4 I__17153 (
            .O(N__74616),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__17152 (
            .O(N__74613),
            .I(N__74610));
    LocalMux I__17151 (
            .O(N__74610),
            .I(N__74607));
    Odrv4 I__17150 (
            .O(N__74607),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__17149 (
            .O(N__74604),
            .I(N__74599));
    InMux I__17148 (
            .O(N__74603),
            .I(N__74594));
    InMux I__17147 (
            .O(N__74602),
            .I(N__74594));
    LocalMux I__17146 (
            .O(N__74599),
            .I(N__74591));
    LocalMux I__17145 (
            .O(N__74594),
            .I(N__74588));
    Span4Mux_h I__17144 (
            .O(N__74591),
            .I(N__74585));
    Span4Mux_h I__17143 (
            .O(N__74588),
            .I(N__74582));
    Span4Mux_v I__17142 (
            .O(N__74585),
            .I(N__74579));
    Span4Mux_v I__17141 (
            .O(N__74582),
            .I(N__74576));
    Odrv4 I__17140 (
            .O(N__74579),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    Odrv4 I__17139 (
            .O(N__74576),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__17138 (
            .O(N__74571),
            .I(N__74565));
    CascadeMux I__17137 (
            .O(N__74570),
            .I(N__74557));
    CascadeMux I__17136 (
            .O(N__74569),
            .I(N__74554));
    CascadeMux I__17135 (
            .O(N__74568),
            .I(N__74551));
    LocalMux I__17134 (
            .O(N__74565),
            .I(N__74547));
    CascadeMux I__17133 (
            .O(N__74564),
            .I(N__74544));
    CascadeMux I__17132 (
            .O(N__74563),
            .I(N__74541));
    CascadeMux I__17131 (
            .O(N__74562),
            .I(N__74537));
    InMux I__17130 (
            .O(N__74561),
            .I(N__74532));
    InMux I__17129 (
            .O(N__74560),
            .I(N__74532));
    InMux I__17128 (
            .O(N__74557),
            .I(N__74529));
    InMux I__17127 (
            .O(N__74554),
            .I(N__74524));
    InMux I__17126 (
            .O(N__74551),
            .I(N__74524));
    InMux I__17125 (
            .O(N__74550),
            .I(N__74521));
    Span4Mux_v I__17124 (
            .O(N__74547),
            .I(N__74518));
    InMux I__17123 (
            .O(N__74544),
            .I(N__74513));
    InMux I__17122 (
            .O(N__74541),
            .I(N__74513));
    InMux I__17121 (
            .O(N__74540),
            .I(N__74508));
    InMux I__17120 (
            .O(N__74537),
            .I(N__74508));
    LocalMux I__17119 (
            .O(N__74532),
            .I(N__74496));
    LocalMux I__17118 (
            .O(N__74529),
            .I(N__74496));
    LocalMux I__17117 (
            .O(N__74524),
            .I(N__74496));
    LocalMux I__17116 (
            .O(N__74521),
            .I(N__74493));
    Span4Mux_h I__17115 (
            .O(N__74518),
            .I(N__74486));
    LocalMux I__17114 (
            .O(N__74513),
            .I(N__74486));
    LocalMux I__17113 (
            .O(N__74508),
            .I(N__74486));
    InMux I__17112 (
            .O(N__74507),
            .I(N__74483));
    CascadeMux I__17111 (
            .O(N__74506),
            .I(N__74480));
    CascadeMux I__17110 (
            .O(N__74505),
            .I(N__74477));
    CascadeMux I__17109 (
            .O(N__74504),
            .I(N__74474));
    CascadeMux I__17108 (
            .O(N__74503),
            .I(N__74470));
    Span4Mux_v I__17107 (
            .O(N__74496),
            .I(N__74464));
    Span4Mux_v I__17106 (
            .O(N__74493),
            .I(N__74464));
    Span4Mux_v I__17105 (
            .O(N__74486),
            .I(N__74461));
    LocalMux I__17104 (
            .O(N__74483),
            .I(N__74458));
    InMux I__17103 (
            .O(N__74480),
            .I(N__74453));
    InMux I__17102 (
            .O(N__74477),
            .I(N__74453));
    InMux I__17101 (
            .O(N__74474),
            .I(N__74450));
    InMux I__17100 (
            .O(N__74473),
            .I(N__74445));
    InMux I__17099 (
            .O(N__74470),
            .I(N__74445));
    InMux I__17098 (
            .O(N__74469),
            .I(N__74442));
    Odrv4 I__17097 (
            .O(N__74464),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__17096 (
            .O(N__74461),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__17095 (
            .O(N__74458),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__17094 (
            .O(N__74453),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__17093 (
            .O(N__74450),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__17092 (
            .O(N__74445),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__17091 (
            .O(N__74442),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    CascadeMux I__17090 (
            .O(N__74427),
            .I(N__74423));
    InMux I__17089 (
            .O(N__74426),
            .I(N__74403));
    InMux I__17088 (
            .O(N__74423),
            .I(N__74403));
    InMux I__17087 (
            .O(N__74422),
            .I(N__74403));
    CascadeMux I__17086 (
            .O(N__74421),
            .I(N__74400));
    InMux I__17085 (
            .O(N__74420),
            .I(N__74395));
    InMux I__17084 (
            .O(N__74419),
            .I(N__74395));
    InMux I__17083 (
            .O(N__74418),
            .I(N__74386));
    InMux I__17082 (
            .O(N__74417),
            .I(N__74386));
    InMux I__17081 (
            .O(N__74416),
            .I(N__74386));
    InMux I__17080 (
            .O(N__74415),
            .I(N__74386));
    InMux I__17079 (
            .O(N__74414),
            .I(N__74379));
    InMux I__17078 (
            .O(N__74413),
            .I(N__74379));
    InMux I__17077 (
            .O(N__74412),
            .I(N__74371));
    InMux I__17076 (
            .O(N__74411),
            .I(N__74371));
    InMux I__17075 (
            .O(N__74410),
            .I(N__74371));
    LocalMux I__17074 (
            .O(N__74403),
            .I(N__74368));
    InMux I__17073 (
            .O(N__74400),
            .I(N__74365));
    LocalMux I__17072 (
            .O(N__74395),
            .I(N__74362));
    LocalMux I__17071 (
            .O(N__74386),
            .I(N__74359));
    InMux I__17070 (
            .O(N__74385),
            .I(N__74354));
    InMux I__17069 (
            .O(N__74384),
            .I(N__74354));
    LocalMux I__17068 (
            .O(N__74379),
            .I(N__74351));
    InMux I__17067 (
            .O(N__74378),
            .I(N__74348));
    LocalMux I__17066 (
            .O(N__74371),
            .I(N__74343));
    Span4Mux_v I__17065 (
            .O(N__74368),
            .I(N__74343));
    LocalMux I__17064 (
            .O(N__74365),
            .I(N__74334));
    Span4Mux_h I__17063 (
            .O(N__74362),
            .I(N__74334));
    Span4Mux_v I__17062 (
            .O(N__74359),
            .I(N__74334));
    LocalMux I__17061 (
            .O(N__74354),
            .I(N__74334));
    Span4Mux_h I__17060 (
            .O(N__74351),
            .I(N__74331));
    LocalMux I__17059 (
            .O(N__74348),
            .I(N__74326));
    Span4Mux_h I__17058 (
            .O(N__74343),
            .I(N__74326));
    Span4Mux_h I__17057 (
            .O(N__74334),
            .I(N__74323));
    Odrv4 I__17056 (
            .O(N__74331),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__17055 (
            .O(N__74326),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__17054 (
            .O(N__74323),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__17053 (
            .O(N__74316),
            .I(N__74313));
    LocalMux I__17052 (
            .O(N__74313),
            .I(N__74310));
    Odrv4 I__17051 (
            .O(N__74310),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__17050 (
            .O(N__74307),
            .I(N__74304));
    LocalMux I__17049 (
            .O(N__74304),
            .I(N__74300));
    InMux I__17048 (
            .O(N__74303),
            .I(N__74296));
    Span4Mux_v I__17047 (
            .O(N__74300),
            .I(N__74293));
    InMux I__17046 (
            .O(N__74299),
            .I(N__74290));
    LocalMux I__17045 (
            .O(N__74296),
            .I(N__74287));
    Span4Mux_v I__17044 (
            .O(N__74293),
            .I(N__74282));
    LocalMux I__17043 (
            .O(N__74290),
            .I(N__74282));
    Odrv4 I__17042 (
            .O(N__74287),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    Odrv4 I__17041 (
            .O(N__74282),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    InMux I__17040 (
            .O(N__74277),
            .I(N__74274));
    LocalMux I__17039 (
            .O(N__74274),
            .I(N__74271));
    Span4Mux_h I__17038 (
            .O(N__74271),
            .I(N__74268));
    Span4Mux_h I__17037 (
            .O(N__74268),
            .I(N__74265));
    Odrv4 I__17036 (
            .O(N__74265),
            .I(\pid_side.O_2_6 ));
    InMux I__17035 (
            .O(N__74262),
            .I(N__74256));
    InMux I__17034 (
            .O(N__74261),
            .I(N__74256));
    LocalMux I__17033 (
            .O(N__74256),
            .I(N__74253));
    Span4Mux_v I__17032 (
            .O(N__74253),
            .I(N__74250));
    Span4Mux_h I__17031 (
            .O(N__74250),
            .I(N__74247));
    Odrv4 I__17030 (
            .O(N__74247),
            .I(\pid_side.error_p_regZ0Z_3 ));
    InMux I__17029 (
            .O(N__74244),
            .I(N__74241));
    LocalMux I__17028 (
            .O(N__74241),
            .I(N__74238));
    Span4Mux_h I__17027 (
            .O(N__74238),
            .I(N__74235));
    Span4Mux_h I__17026 (
            .O(N__74235),
            .I(N__74232));
    Odrv4 I__17025 (
            .O(N__74232),
            .I(\pid_side.O_2_5 ));
    InMux I__17024 (
            .O(N__74229),
            .I(N__74226));
    LocalMux I__17023 (
            .O(N__74226),
            .I(N__74222));
    InMux I__17022 (
            .O(N__74225),
            .I(N__74219));
    Span4Mux_v I__17021 (
            .O(N__74222),
            .I(N__74216));
    LocalMux I__17020 (
            .O(N__74219),
            .I(N__74213));
    Span4Mux_h I__17019 (
            .O(N__74216),
            .I(N__74207));
    Span4Mux_h I__17018 (
            .O(N__74213),
            .I(N__74207));
    InMux I__17017 (
            .O(N__74212),
            .I(N__74204));
    Odrv4 I__17016 (
            .O(N__74207),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__17015 (
            .O(N__74204),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__17014 (
            .O(N__74199),
            .I(N__74196));
    LocalMux I__17013 (
            .O(N__74196),
            .I(N__74193));
    Span4Mux_v I__17012 (
            .O(N__74193),
            .I(N__74188));
    InMux I__17011 (
            .O(N__74192),
            .I(N__74183));
    InMux I__17010 (
            .O(N__74191),
            .I(N__74183));
    Odrv4 I__17009 (
            .O(N__74188),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__17008 (
            .O(N__74183),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    InMux I__17007 (
            .O(N__74178),
            .I(N__74169));
    InMux I__17006 (
            .O(N__74177),
            .I(N__74169));
    CascadeMux I__17005 (
            .O(N__74176),
            .I(N__74165));
    CascadeMux I__17004 (
            .O(N__74175),
            .I(N__74161));
    CascadeMux I__17003 (
            .O(N__74174),
            .I(N__74158));
    LocalMux I__17002 (
            .O(N__74169),
            .I(N__74155));
    CascadeMux I__17001 (
            .O(N__74168),
            .I(N__74151));
    InMux I__17000 (
            .O(N__74165),
            .I(N__74145));
    InMux I__16999 (
            .O(N__74164),
            .I(N__74145));
    InMux I__16998 (
            .O(N__74161),
            .I(N__74140));
    InMux I__16997 (
            .O(N__74158),
            .I(N__74140));
    Span4Mux_v I__16996 (
            .O(N__74155),
            .I(N__74137));
    InMux I__16995 (
            .O(N__74154),
            .I(N__74134));
    InMux I__16994 (
            .O(N__74151),
            .I(N__74129));
    InMux I__16993 (
            .O(N__74150),
            .I(N__74129));
    LocalMux I__16992 (
            .O(N__74145),
            .I(N__74126));
    LocalMux I__16991 (
            .O(N__74140),
            .I(N__74117));
    Sp12to4 I__16990 (
            .O(N__74137),
            .I(N__74117));
    LocalMux I__16989 (
            .O(N__74134),
            .I(N__74117));
    LocalMux I__16988 (
            .O(N__74129),
            .I(N__74117));
    Span12Mux_v I__16987 (
            .O(N__74126),
            .I(N__74114));
    Odrv12 I__16986 (
            .O(N__74117),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    Odrv12 I__16985 (
            .O(N__74114),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    InMux I__16984 (
            .O(N__74109),
            .I(N__74105));
    InMux I__16983 (
            .O(N__74108),
            .I(N__74102));
    LocalMux I__16982 (
            .O(N__74105),
            .I(N__74099));
    LocalMux I__16981 (
            .O(N__74102),
            .I(N__74096));
    Span4Mux_h I__16980 (
            .O(N__74099),
            .I(N__74092));
    Span4Mux_h I__16979 (
            .O(N__74096),
            .I(N__74089));
    InMux I__16978 (
            .O(N__74095),
            .I(N__74086));
    Odrv4 I__16977 (
            .O(N__74092),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__16976 (
            .O(N__74089),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__16975 (
            .O(N__74086),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    InMux I__16974 (
            .O(N__74079),
            .I(N__74076));
    LocalMux I__16973 (
            .O(N__74076),
            .I(N__74073));
    Odrv4 I__16972 (
            .O(N__74073),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__16971 (
            .O(N__74070),
            .I(N__74066));
    CascadeMux I__16970 (
            .O(N__74069),
            .I(N__74063));
    LocalMux I__16969 (
            .O(N__74066),
            .I(N__74060));
    InMux I__16968 (
            .O(N__74063),
            .I(N__74057));
    Span4Mux_h I__16967 (
            .O(N__74060),
            .I(N__74054));
    LocalMux I__16966 (
            .O(N__74057),
            .I(N__74051));
    Odrv4 I__16965 (
            .O(N__74054),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    Odrv12 I__16964 (
            .O(N__74051),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    InMux I__16963 (
            .O(N__74046),
            .I(N__74037));
    InMux I__16962 (
            .O(N__74045),
            .I(N__74037));
    InMux I__16961 (
            .O(N__74044),
            .I(N__74037));
    LocalMux I__16960 (
            .O(N__74037),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__16959 (
            .O(N__74034),
            .I(N__74031));
    LocalMux I__16958 (
            .O(N__74031),
            .I(N__74027));
    InMux I__16957 (
            .O(N__74030),
            .I(N__74023));
    Span12Mux_h I__16956 (
            .O(N__74027),
            .I(N__74020));
    InMux I__16955 (
            .O(N__74026),
            .I(N__74017));
    LocalMux I__16954 (
            .O(N__74023),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv12 I__16953 (
            .O(N__74020),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    LocalMux I__16952 (
            .O(N__74017),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    InMux I__16951 (
            .O(N__74010),
            .I(N__74007));
    LocalMux I__16950 (
            .O(N__74007),
            .I(N__74004));
    Span4Mux_h I__16949 (
            .O(N__74004),
            .I(N__74001));
    Span4Mux_h I__16948 (
            .O(N__74001),
            .I(N__73998));
    Odrv4 I__16947 (
            .O(N__73998),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__16946 (
            .O(N__73995),
            .I(N__73992));
    LocalMux I__16945 (
            .O(N__73992),
            .I(N__73989));
    Odrv4 I__16944 (
            .O(N__73989),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__16943 (
            .O(N__73986),
            .I(N__73983));
    LocalMux I__16942 (
            .O(N__73983),
            .I(N__73980));
    Span4Mux_v I__16941 (
            .O(N__73980),
            .I(N__73977));
    Span4Mux_h I__16940 (
            .O(N__73977),
            .I(N__73972));
    InMux I__16939 (
            .O(N__73976),
            .I(N__73969));
    InMux I__16938 (
            .O(N__73975),
            .I(N__73966));
    Odrv4 I__16937 (
            .O(N__73972),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    LocalMux I__16936 (
            .O(N__73969),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    LocalMux I__16935 (
            .O(N__73966),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    CascadeMux I__16934 (
            .O(N__73959),
            .I(N__73955));
    InMux I__16933 (
            .O(N__73958),
            .I(N__73952));
    InMux I__16932 (
            .O(N__73955),
            .I(N__73949));
    LocalMux I__16931 (
            .O(N__73952),
            .I(N__73946));
    LocalMux I__16930 (
            .O(N__73949),
            .I(N__73943));
    Odrv12 I__16929 (
            .O(N__73946),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    Odrv4 I__16928 (
            .O(N__73943),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    CascadeMux I__16927 (
            .O(N__73938),
            .I(\ppm_encoder_1.un1_init_pulses_0_1_cascade_ ));
    InMux I__16926 (
            .O(N__73935),
            .I(N__73930));
    InMux I__16925 (
            .O(N__73934),
            .I(N__73927));
    CascadeMux I__16924 (
            .O(N__73933),
            .I(N__73924));
    LocalMux I__16923 (
            .O(N__73930),
            .I(N__73920));
    LocalMux I__16922 (
            .O(N__73927),
            .I(N__73917));
    InMux I__16921 (
            .O(N__73924),
            .I(N__73914));
    InMux I__16920 (
            .O(N__73923),
            .I(N__73911));
    Span4Mux_h I__16919 (
            .O(N__73920),
            .I(N__73908));
    Span4Mux_h I__16918 (
            .O(N__73917),
            .I(N__73905));
    LocalMux I__16917 (
            .O(N__73914),
            .I(N__73900));
    LocalMux I__16916 (
            .O(N__73911),
            .I(N__73900));
    Span4Mux_v I__16915 (
            .O(N__73908),
            .I(N__73897));
    Odrv4 I__16914 (
            .O(N__73905),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv12 I__16913 (
            .O(N__73900),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__16912 (
            .O(N__73897),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__16911 (
            .O(N__73890),
            .I(N__73887));
    LocalMux I__16910 (
            .O(N__73887),
            .I(N__73884));
    Span4Mux_h I__16909 (
            .O(N__73884),
            .I(N__73881));
    Odrv4 I__16908 (
            .O(N__73881),
            .I(\ppm_encoder_1.un1_init_pulses_11_0 ));
    InMux I__16907 (
            .O(N__73878),
            .I(N__73874));
    InMux I__16906 (
            .O(N__73877),
            .I(N__73871));
    LocalMux I__16905 (
            .O(N__73874),
            .I(N__73867));
    LocalMux I__16904 (
            .O(N__73871),
            .I(N__73864));
    InMux I__16903 (
            .O(N__73870),
            .I(N__73861));
    Span4Mux_h I__16902 (
            .O(N__73867),
            .I(N__73858));
    Span4Mux_h I__16901 (
            .O(N__73864),
            .I(N__73855));
    LocalMux I__16900 (
            .O(N__73861),
            .I(N__73852));
    Span4Mux_h I__16899 (
            .O(N__73858),
            .I(N__73847));
    Span4Mux_v I__16898 (
            .O(N__73855),
            .I(N__73847));
    Odrv12 I__16897 (
            .O(N__73852),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__16896 (
            .O(N__73847),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__16895 (
            .O(N__73842),
            .I(N__73839));
    LocalMux I__16894 (
            .O(N__73839),
            .I(N__73836));
    Span4Mux_h I__16893 (
            .O(N__73836),
            .I(N__73833));
    Odrv4 I__16892 (
            .O(N__73833),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__16891 (
            .O(N__73830),
            .I(N__73827));
    LocalMux I__16890 (
            .O(N__73827),
            .I(N__73824));
    Span12Mux_h I__16889 (
            .O(N__73824),
            .I(N__73819));
    InMux I__16888 (
            .O(N__73823),
            .I(N__73816));
    InMux I__16887 (
            .O(N__73822),
            .I(N__73813));
    Span12Mux_v I__16886 (
            .O(N__73819),
            .I(N__73810));
    LocalMux I__16885 (
            .O(N__73816),
            .I(N__73805));
    LocalMux I__16884 (
            .O(N__73813),
            .I(N__73805));
    Odrv12 I__16883 (
            .O(N__73810),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    Odrv4 I__16882 (
            .O(N__73805),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    InMux I__16881 (
            .O(N__73800),
            .I(N__73797));
    LocalMux I__16880 (
            .O(N__73797),
            .I(N__73794));
    Span4Mux_h I__16879 (
            .O(N__73794),
            .I(N__73791));
    Odrv4 I__16878 (
            .O(N__73791),
            .I(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ));
    InMux I__16877 (
            .O(N__73788),
            .I(N__73784));
    InMux I__16876 (
            .O(N__73787),
            .I(N__73781));
    LocalMux I__16875 (
            .O(N__73784),
            .I(N__73778));
    LocalMux I__16874 (
            .O(N__73781),
            .I(N__73775));
    Span4Mux_h I__16873 (
            .O(N__73778),
            .I(N__73772));
    Span4Mux_v I__16872 (
            .O(N__73775),
            .I(N__73764));
    Span4Mux_h I__16871 (
            .O(N__73772),
            .I(N__73764));
    InMux I__16870 (
            .O(N__73771),
            .I(N__73761));
    InMux I__16869 (
            .O(N__73770),
            .I(N__73756));
    InMux I__16868 (
            .O(N__73769),
            .I(N__73756));
    Span4Mux_h I__16867 (
            .O(N__73764),
            .I(N__73751));
    LocalMux I__16866 (
            .O(N__73761),
            .I(N__73751));
    LocalMux I__16865 (
            .O(N__73756),
            .I(N__73747));
    Span4Mux_v I__16864 (
            .O(N__73751),
            .I(N__73744));
    InMux I__16863 (
            .O(N__73750),
            .I(N__73741));
    Span4Mux_h I__16862 (
            .O(N__73747),
            .I(N__73732));
    Span4Mux_h I__16861 (
            .O(N__73744),
            .I(N__73732));
    LocalMux I__16860 (
            .O(N__73741),
            .I(N__73732));
    InMux I__16859 (
            .O(N__73740),
            .I(N__73729));
    InMux I__16858 (
            .O(N__73739),
            .I(N__73722));
    Span4Mux_v I__16857 (
            .O(N__73732),
            .I(N__73718));
    LocalMux I__16856 (
            .O(N__73729),
            .I(N__73714));
    InMux I__16855 (
            .O(N__73728),
            .I(N__73711));
    InMux I__16854 (
            .O(N__73727),
            .I(N__73708));
    InMux I__16853 (
            .O(N__73726),
            .I(N__73705));
    InMux I__16852 (
            .O(N__73725),
            .I(N__73702));
    LocalMux I__16851 (
            .O(N__73722),
            .I(N__73699));
    InMux I__16850 (
            .O(N__73721),
            .I(N__73696));
    Span4Mux_v I__16849 (
            .O(N__73718),
            .I(N__73693));
    InMux I__16848 (
            .O(N__73717),
            .I(N__73689));
    Span4Mux_v I__16847 (
            .O(N__73714),
            .I(N__73686));
    LocalMux I__16846 (
            .O(N__73711),
            .I(N__73683));
    LocalMux I__16845 (
            .O(N__73708),
            .I(N__73680));
    LocalMux I__16844 (
            .O(N__73705),
            .I(N__73677));
    LocalMux I__16843 (
            .O(N__73702),
            .I(N__73674));
    Span4Mux_v I__16842 (
            .O(N__73699),
            .I(N__73671));
    LocalMux I__16841 (
            .O(N__73696),
            .I(N__73666));
    Span4Mux_v I__16840 (
            .O(N__73693),
            .I(N__73666));
    InMux I__16839 (
            .O(N__73692),
            .I(N__73663));
    LocalMux I__16838 (
            .O(N__73689),
            .I(N__73659));
    Span4Mux_h I__16837 (
            .O(N__73686),
            .I(N__73654));
    Span4Mux_h I__16836 (
            .O(N__73683),
            .I(N__73654));
    Span4Mux_v I__16835 (
            .O(N__73680),
            .I(N__73649));
    Span4Mux_v I__16834 (
            .O(N__73677),
            .I(N__73649));
    Sp12to4 I__16833 (
            .O(N__73674),
            .I(N__73646));
    Sp12to4 I__16832 (
            .O(N__73671),
            .I(N__73643));
    Span4Mux_h I__16831 (
            .O(N__73666),
            .I(N__73640));
    LocalMux I__16830 (
            .O(N__73663),
            .I(N__73637));
    InMux I__16829 (
            .O(N__73662),
            .I(N__73634));
    Span4Mux_h I__16828 (
            .O(N__73659),
            .I(N__73631));
    Span4Mux_v I__16827 (
            .O(N__73654),
            .I(N__73628));
    Sp12to4 I__16826 (
            .O(N__73649),
            .I(N__73623));
    Span12Mux_v I__16825 (
            .O(N__73646),
            .I(N__73623));
    Span12Mux_s8_h I__16824 (
            .O(N__73643),
            .I(N__73620));
    Span4Mux_h I__16823 (
            .O(N__73640),
            .I(N__73615));
    Span4Mux_v I__16822 (
            .O(N__73637),
            .I(N__73615));
    LocalMux I__16821 (
            .O(N__73634),
            .I(uart_pc_data_1));
    Odrv4 I__16820 (
            .O(N__73631),
            .I(uart_pc_data_1));
    Odrv4 I__16819 (
            .O(N__73628),
            .I(uart_pc_data_1));
    Odrv12 I__16818 (
            .O(N__73623),
            .I(uart_pc_data_1));
    Odrv12 I__16817 (
            .O(N__73620),
            .I(uart_pc_data_1));
    Odrv4 I__16816 (
            .O(N__73615),
            .I(uart_pc_data_1));
    CascadeMux I__16815 (
            .O(N__73602),
            .I(N__73596));
    InMux I__16814 (
            .O(N__73601),
            .I(N__73587));
    CascadeMux I__16813 (
            .O(N__73600),
            .I(N__73584));
    CascadeMux I__16812 (
            .O(N__73599),
            .I(N__73581));
    InMux I__16811 (
            .O(N__73596),
            .I(N__73575));
    InMux I__16810 (
            .O(N__73595),
            .I(N__73575));
    InMux I__16809 (
            .O(N__73594),
            .I(N__73569));
    InMux I__16808 (
            .O(N__73593),
            .I(N__73564));
    InMux I__16807 (
            .O(N__73592),
            .I(N__73561));
    InMux I__16806 (
            .O(N__73591),
            .I(N__73556));
    InMux I__16805 (
            .O(N__73590),
            .I(N__73556));
    LocalMux I__16804 (
            .O(N__73587),
            .I(N__73553));
    InMux I__16803 (
            .O(N__73584),
            .I(N__73548));
    InMux I__16802 (
            .O(N__73581),
            .I(N__73548));
    InMux I__16801 (
            .O(N__73580),
            .I(N__73545));
    LocalMux I__16800 (
            .O(N__73575),
            .I(N__73541));
    InMux I__16799 (
            .O(N__73574),
            .I(N__73536));
    InMux I__16798 (
            .O(N__73573),
            .I(N__73536));
    InMux I__16797 (
            .O(N__73572),
            .I(N__73532));
    LocalMux I__16796 (
            .O(N__73569),
            .I(N__73529));
    InMux I__16795 (
            .O(N__73568),
            .I(N__73524));
    InMux I__16794 (
            .O(N__73567),
            .I(N__73524));
    LocalMux I__16793 (
            .O(N__73564),
            .I(N__73521));
    LocalMux I__16792 (
            .O(N__73561),
            .I(N__73518));
    LocalMux I__16791 (
            .O(N__73556),
            .I(N__73515));
    Span4Mux_v I__16790 (
            .O(N__73553),
            .I(N__73508));
    LocalMux I__16789 (
            .O(N__73548),
            .I(N__73508));
    LocalMux I__16788 (
            .O(N__73545),
            .I(N__73508));
    InMux I__16787 (
            .O(N__73544),
            .I(N__73500));
    Span4Mux_h I__16786 (
            .O(N__73541),
            .I(N__73495));
    LocalMux I__16785 (
            .O(N__73536),
            .I(N__73495));
    InMux I__16784 (
            .O(N__73535),
            .I(N__73492));
    LocalMux I__16783 (
            .O(N__73532),
            .I(N__73489));
    Span12Mux_s10_h I__16782 (
            .O(N__73529),
            .I(N__73484));
    LocalMux I__16781 (
            .O(N__73524),
            .I(N__73481));
    Span4Mux_h I__16780 (
            .O(N__73521),
            .I(N__73472));
    Span4Mux_v I__16779 (
            .O(N__73518),
            .I(N__73472));
    Span4Mux_v I__16778 (
            .O(N__73515),
            .I(N__73472));
    Span4Mux_h I__16777 (
            .O(N__73508),
            .I(N__73472));
    InMux I__16776 (
            .O(N__73507),
            .I(N__73465));
    InMux I__16775 (
            .O(N__73506),
            .I(N__73465));
    InMux I__16774 (
            .O(N__73505),
            .I(N__73465));
    InMux I__16773 (
            .O(N__73504),
            .I(N__73462));
    InMux I__16772 (
            .O(N__73503),
            .I(N__73459));
    LocalMux I__16771 (
            .O(N__73500),
            .I(N__73454));
    Span4Mux_h I__16770 (
            .O(N__73495),
            .I(N__73454));
    LocalMux I__16769 (
            .O(N__73492),
            .I(N__73449));
    Span4Mux_v I__16768 (
            .O(N__73489),
            .I(N__73449));
    InMux I__16767 (
            .O(N__73488),
            .I(N__73446));
    InMux I__16766 (
            .O(N__73487),
            .I(N__73443));
    Span12Mux_v I__16765 (
            .O(N__73484),
            .I(N__73438));
    Span12Mux_h I__16764 (
            .O(N__73481),
            .I(N__73438));
    Span4Mux_h I__16763 (
            .O(N__73472),
            .I(N__73435));
    LocalMux I__16762 (
            .O(N__73465),
            .I(N__73424));
    LocalMux I__16761 (
            .O(N__73462),
            .I(N__73424));
    LocalMux I__16760 (
            .O(N__73459),
            .I(N__73424));
    Span4Mux_h I__16759 (
            .O(N__73454),
            .I(N__73424));
    Span4Mux_h I__16758 (
            .O(N__73449),
            .I(N__73424));
    LocalMux I__16757 (
            .O(N__73446),
            .I(xy_ki_1));
    LocalMux I__16756 (
            .O(N__73443),
            .I(xy_ki_1));
    Odrv12 I__16755 (
            .O(N__73438),
            .I(xy_ki_1));
    Odrv4 I__16754 (
            .O(N__73435),
            .I(xy_ki_1));
    Odrv4 I__16753 (
            .O(N__73424),
            .I(xy_ki_1));
    CEMux I__16752 (
            .O(N__73413),
            .I(N__73408));
    CEMux I__16751 (
            .O(N__73412),
            .I(N__73405));
    CEMux I__16750 (
            .O(N__73411),
            .I(N__73399));
    LocalMux I__16749 (
            .O(N__73408),
            .I(N__73396));
    LocalMux I__16748 (
            .O(N__73405),
            .I(N__73393));
    CEMux I__16747 (
            .O(N__73404),
            .I(N__73390));
    CEMux I__16746 (
            .O(N__73403),
            .I(N__73387));
    CEMux I__16745 (
            .O(N__73402),
            .I(N__73384));
    LocalMux I__16744 (
            .O(N__73399),
            .I(N__73380));
    Span4Mux_v I__16743 (
            .O(N__73396),
            .I(N__73377));
    Span4Mux_v I__16742 (
            .O(N__73393),
            .I(N__73372));
    LocalMux I__16741 (
            .O(N__73390),
            .I(N__73372));
    LocalMux I__16740 (
            .O(N__73387),
            .I(N__73369));
    LocalMux I__16739 (
            .O(N__73384),
            .I(N__73366));
    CEMux I__16738 (
            .O(N__73383),
            .I(N__73363));
    Span4Mux_v I__16737 (
            .O(N__73380),
            .I(N__73360));
    Span4Mux_v I__16736 (
            .O(N__73377),
            .I(N__73357));
    Span4Mux_v I__16735 (
            .O(N__73372),
            .I(N__73354));
    Span4Mux_h I__16734 (
            .O(N__73369),
            .I(N__73349));
    Span4Mux_v I__16733 (
            .O(N__73366),
            .I(N__73349));
    LocalMux I__16732 (
            .O(N__73363),
            .I(N__73346));
    Span4Mux_v I__16731 (
            .O(N__73360),
            .I(N__73341));
    Span4Mux_v I__16730 (
            .O(N__73357),
            .I(N__73341));
    Span4Mux_h I__16729 (
            .O(N__73354),
            .I(N__73336));
    Span4Mux_v I__16728 (
            .O(N__73349),
            .I(N__73336));
    Span4Mux_h I__16727 (
            .O(N__73346),
            .I(N__73333));
    Span4Mux_h I__16726 (
            .O(N__73341),
            .I(N__73330));
    Span4Mux_v I__16725 (
            .O(N__73336),
            .I(N__73327));
    Span4Mux_h I__16724 (
            .O(N__73333),
            .I(N__73324));
    Odrv4 I__16723 (
            .O(N__73330),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__16722 (
            .O(N__73327),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__16721 (
            .O(N__73324),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    CascadeMux I__16720 (
            .O(N__73317),
            .I(\pid_side.g0_3_1_cascade_ ));
    InMux I__16719 (
            .O(N__73314),
            .I(N__73311));
    LocalMux I__16718 (
            .O(N__73311),
            .I(\pid_side.N_28_1_0 ));
    InMux I__16717 (
            .O(N__73308),
            .I(N__73300));
    CascadeMux I__16716 (
            .O(N__73307),
            .I(N__73296));
    CascadeMux I__16715 (
            .O(N__73306),
            .I(N__73292));
    CascadeMux I__16714 (
            .O(N__73305),
            .I(N__73289));
    CascadeMux I__16713 (
            .O(N__73304),
            .I(N__73283));
    CascadeMux I__16712 (
            .O(N__73303),
            .I(N__73280));
    LocalMux I__16711 (
            .O(N__73300),
            .I(N__73277));
    CascadeMux I__16710 (
            .O(N__73299),
            .I(N__73274));
    InMux I__16709 (
            .O(N__73296),
            .I(N__73271));
    InMux I__16708 (
            .O(N__73295),
            .I(N__73266));
    InMux I__16707 (
            .O(N__73292),
            .I(N__73266));
    InMux I__16706 (
            .O(N__73289),
            .I(N__73263));
    InMux I__16705 (
            .O(N__73288),
            .I(N__73258));
    InMux I__16704 (
            .O(N__73287),
            .I(N__73258));
    InMux I__16703 (
            .O(N__73286),
            .I(N__73255));
    InMux I__16702 (
            .O(N__73283),
            .I(N__73251));
    InMux I__16701 (
            .O(N__73280),
            .I(N__73248));
    Span4Mux_v I__16700 (
            .O(N__73277),
            .I(N__73245));
    InMux I__16699 (
            .O(N__73274),
            .I(N__73242));
    LocalMux I__16698 (
            .O(N__73271),
            .I(N__73237));
    LocalMux I__16697 (
            .O(N__73266),
            .I(N__73237));
    LocalMux I__16696 (
            .O(N__73263),
            .I(N__73234));
    LocalMux I__16695 (
            .O(N__73258),
            .I(N__73229));
    LocalMux I__16694 (
            .O(N__73255),
            .I(N__73229));
    InMux I__16693 (
            .O(N__73254),
            .I(N__73224));
    LocalMux I__16692 (
            .O(N__73251),
            .I(N__73221));
    LocalMux I__16691 (
            .O(N__73248),
            .I(N__73214));
    Span4Mux_h I__16690 (
            .O(N__73245),
            .I(N__73214));
    LocalMux I__16689 (
            .O(N__73242),
            .I(N__73214));
    Span4Mux_v I__16688 (
            .O(N__73237),
            .I(N__73207));
    Span4Mux_v I__16687 (
            .O(N__73234),
            .I(N__73207));
    Span4Mux_v I__16686 (
            .O(N__73229),
            .I(N__73207));
    InMux I__16685 (
            .O(N__73228),
            .I(N__73202));
    InMux I__16684 (
            .O(N__73227),
            .I(N__73199));
    LocalMux I__16683 (
            .O(N__73224),
            .I(N__73194));
    Span4Mux_h I__16682 (
            .O(N__73221),
            .I(N__73194));
    Span4Mux_h I__16681 (
            .O(N__73214),
            .I(N__73191));
    Span4Mux_h I__16680 (
            .O(N__73207),
            .I(N__73188));
    InMux I__16679 (
            .O(N__73206),
            .I(N__73183));
    InMux I__16678 (
            .O(N__73205),
            .I(N__73183));
    LocalMux I__16677 (
            .O(N__73202),
            .I(xy_ki_fast_1));
    LocalMux I__16676 (
            .O(N__73199),
            .I(xy_ki_fast_1));
    Odrv4 I__16675 (
            .O(N__73194),
            .I(xy_ki_fast_1));
    Odrv4 I__16674 (
            .O(N__73191),
            .I(xy_ki_fast_1));
    Odrv4 I__16673 (
            .O(N__73188),
            .I(xy_ki_fast_1));
    LocalMux I__16672 (
            .O(N__73183),
            .I(xy_ki_fast_1));
    InMux I__16671 (
            .O(N__73170),
            .I(N__73167));
    LocalMux I__16670 (
            .O(N__73167),
            .I(N__73162));
    InMux I__16669 (
            .O(N__73166),
            .I(N__73155));
    InMux I__16668 (
            .O(N__73165),
            .I(N__73151));
    Span4Mux_s2_h I__16667 (
            .O(N__73162),
            .I(N__73148));
    InMux I__16666 (
            .O(N__73161),
            .I(N__73145));
    InMux I__16665 (
            .O(N__73160),
            .I(N__73140));
    InMux I__16664 (
            .O(N__73159),
            .I(N__73140));
    InMux I__16663 (
            .O(N__73158),
            .I(N__73137));
    LocalMux I__16662 (
            .O(N__73155),
            .I(N__73133));
    InMux I__16661 (
            .O(N__73154),
            .I(N__73130));
    LocalMux I__16660 (
            .O(N__73151),
            .I(N__73127));
    Span4Mux_v I__16659 (
            .O(N__73148),
            .I(N__73124));
    LocalMux I__16658 (
            .O(N__73145),
            .I(N__73121));
    LocalMux I__16657 (
            .O(N__73140),
            .I(N__73118));
    LocalMux I__16656 (
            .O(N__73137),
            .I(N__73115));
    InMux I__16655 (
            .O(N__73136),
            .I(N__73112));
    Span4Mux_h I__16654 (
            .O(N__73133),
            .I(N__73109));
    LocalMux I__16653 (
            .O(N__73130),
            .I(N__73104));
    Span12Mux_s7_h I__16652 (
            .O(N__73127),
            .I(N__73104));
    Span4Mux_h I__16651 (
            .O(N__73124),
            .I(N__73101));
    Span4Mux_v I__16650 (
            .O(N__73121),
            .I(N__73096));
    Span4Mux_v I__16649 (
            .O(N__73118),
            .I(N__73096));
    Span4Mux_v I__16648 (
            .O(N__73115),
            .I(N__73091));
    LocalMux I__16647 (
            .O(N__73112),
            .I(N__73091));
    Odrv4 I__16646 (
            .O(N__73109),
            .I(\pid_side.error_2 ));
    Odrv12 I__16645 (
            .O(N__73104),
            .I(\pid_side.error_2 ));
    Odrv4 I__16644 (
            .O(N__73101),
            .I(\pid_side.error_2 ));
    Odrv4 I__16643 (
            .O(N__73096),
            .I(\pid_side.error_2 ));
    Odrv4 I__16642 (
            .O(N__73091),
            .I(\pid_side.error_2 ));
    InMux I__16641 (
            .O(N__73080),
            .I(N__73077));
    LocalMux I__16640 (
            .O(N__73077),
            .I(\pid_side.m11_0_ns_1_0 ));
    InMux I__16639 (
            .O(N__73074),
            .I(N__73071));
    LocalMux I__16638 (
            .O(N__73071),
            .I(N__73065));
    InMux I__16637 (
            .O(N__73070),
            .I(N__73062));
    InMux I__16636 (
            .O(N__73069),
            .I(N__73059));
    InMux I__16635 (
            .O(N__73068),
            .I(N__73056));
    Span4Mux_v I__16634 (
            .O(N__73065),
            .I(N__73046));
    LocalMux I__16633 (
            .O(N__73062),
            .I(N__73046));
    LocalMux I__16632 (
            .O(N__73059),
            .I(N__73043));
    LocalMux I__16631 (
            .O(N__73056),
            .I(N__73040));
    InMux I__16630 (
            .O(N__73055),
            .I(N__73037));
    InMux I__16629 (
            .O(N__73054),
            .I(N__73034));
    InMux I__16628 (
            .O(N__73053),
            .I(N__73031));
    InMux I__16627 (
            .O(N__73052),
            .I(N__73026));
    InMux I__16626 (
            .O(N__73051),
            .I(N__73026));
    Span4Mux_v I__16625 (
            .O(N__73046),
            .I(N__73023));
    Span4Mux_v I__16624 (
            .O(N__73043),
            .I(N__73012));
    Span4Mux_h I__16623 (
            .O(N__73040),
            .I(N__73012));
    LocalMux I__16622 (
            .O(N__73037),
            .I(N__73012));
    LocalMux I__16621 (
            .O(N__73034),
            .I(N__73012));
    LocalMux I__16620 (
            .O(N__73031),
            .I(N__73012));
    LocalMux I__16619 (
            .O(N__73026),
            .I(N__73009));
    Span4Mux_h I__16618 (
            .O(N__73023),
            .I(N__73004));
    Span4Mux_v I__16617 (
            .O(N__73012),
            .I(N__73004));
    Odrv12 I__16616 (
            .O(N__73009),
            .I(\pid_side.error_3 ));
    Odrv4 I__16615 (
            .O(N__73004),
            .I(\pid_side.error_3 ));
    CascadeMux I__16614 (
            .O(N__72999),
            .I(N__72995));
    CascadeMux I__16613 (
            .O(N__72998),
            .I(N__72985));
    InMux I__16612 (
            .O(N__72995),
            .I(N__72978));
    InMux I__16611 (
            .O(N__72994),
            .I(N__72973));
    InMux I__16610 (
            .O(N__72993),
            .I(N__72973));
    InMux I__16609 (
            .O(N__72992),
            .I(N__72968));
    InMux I__16608 (
            .O(N__72991),
            .I(N__72965));
    InMux I__16607 (
            .O(N__72990),
            .I(N__72960));
    InMux I__16606 (
            .O(N__72989),
            .I(N__72960));
    InMux I__16605 (
            .O(N__72988),
            .I(N__72951));
    InMux I__16604 (
            .O(N__72985),
            .I(N__72951));
    InMux I__16603 (
            .O(N__72984),
            .I(N__72951));
    InMux I__16602 (
            .O(N__72983),
            .I(N__72948));
    InMux I__16601 (
            .O(N__72982),
            .I(N__72943));
    InMux I__16600 (
            .O(N__72981),
            .I(N__72943));
    LocalMux I__16599 (
            .O(N__72978),
            .I(N__72940));
    LocalMux I__16598 (
            .O(N__72973),
            .I(N__72937));
    InMux I__16597 (
            .O(N__72972),
            .I(N__72934));
    InMux I__16596 (
            .O(N__72971),
            .I(N__72931));
    LocalMux I__16595 (
            .O(N__72968),
            .I(N__72928));
    LocalMux I__16594 (
            .O(N__72965),
            .I(N__72923));
    LocalMux I__16593 (
            .O(N__72960),
            .I(N__72923));
    InMux I__16592 (
            .O(N__72959),
            .I(N__72919));
    CascadeMux I__16591 (
            .O(N__72958),
            .I(N__72915));
    LocalMux I__16590 (
            .O(N__72951),
            .I(N__72912));
    LocalMux I__16589 (
            .O(N__72948),
            .I(N__72909));
    LocalMux I__16588 (
            .O(N__72943),
            .I(N__72904));
    Span4Mux_v I__16587 (
            .O(N__72940),
            .I(N__72901));
    Span4Mux_v I__16586 (
            .O(N__72937),
            .I(N__72898));
    LocalMux I__16585 (
            .O(N__72934),
            .I(N__72895));
    LocalMux I__16584 (
            .O(N__72931),
            .I(N__72888));
    Span4Mux_v I__16583 (
            .O(N__72928),
            .I(N__72888));
    Span4Mux_h I__16582 (
            .O(N__72923),
            .I(N__72888));
    CascadeMux I__16581 (
            .O(N__72922),
            .I(N__72880));
    LocalMux I__16580 (
            .O(N__72919),
            .I(N__72877));
    InMux I__16579 (
            .O(N__72918),
            .I(N__72872));
    InMux I__16578 (
            .O(N__72915),
            .I(N__72872));
    Span4Mux_v I__16577 (
            .O(N__72912),
            .I(N__72867));
    Span4Mux_v I__16576 (
            .O(N__72909),
            .I(N__72867));
    InMux I__16575 (
            .O(N__72908),
            .I(N__72864));
    InMux I__16574 (
            .O(N__72907),
            .I(N__72861));
    Span4Mux_v I__16573 (
            .O(N__72904),
            .I(N__72854));
    Span4Mux_h I__16572 (
            .O(N__72901),
            .I(N__72854));
    Span4Mux_h I__16571 (
            .O(N__72898),
            .I(N__72854));
    Span4Mux_v I__16570 (
            .O(N__72895),
            .I(N__72849));
    Span4Mux_h I__16569 (
            .O(N__72888),
            .I(N__72849));
    InMux I__16568 (
            .O(N__72887),
            .I(N__72840));
    InMux I__16567 (
            .O(N__72886),
            .I(N__72840));
    InMux I__16566 (
            .O(N__72885),
            .I(N__72840));
    InMux I__16565 (
            .O(N__72884),
            .I(N__72840));
    InMux I__16564 (
            .O(N__72883),
            .I(N__72835));
    InMux I__16563 (
            .O(N__72880),
            .I(N__72835));
    Span4Mux_h I__16562 (
            .O(N__72877),
            .I(N__72830));
    LocalMux I__16561 (
            .O(N__72872),
            .I(N__72830));
    Span4Mux_h I__16560 (
            .O(N__72867),
            .I(N__72825));
    LocalMux I__16559 (
            .O(N__72864),
            .I(N__72825));
    LocalMux I__16558 (
            .O(N__72861),
            .I(xy_ki_1_rep1));
    Odrv4 I__16557 (
            .O(N__72854),
            .I(xy_ki_1_rep1));
    Odrv4 I__16556 (
            .O(N__72849),
            .I(xy_ki_1_rep1));
    LocalMux I__16555 (
            .O(N__72840),
            .I(xy_ki_1_rep1));
    LocalMux I__16554 (
            .O(N__72835),
            .I(xy_ki_1_rep1));
    Odrv4 I__16553 (
            .O(N__72830),
            .I(xy_ki_1_rep1));
    Odrv4 I__16552 (
            .O(N__72825),
            .I(xy_ki_1_rep1));
    CascadeMux I__16551 (
            .O(N__72810),
            .I(N__72807));
    InMux I__16550 (
            .O(N__72807),
            .I(N__72804));
    LocalMux I__16549 (
            .O(N__72804),
            .I(\pid_side.m30_1_ns_1_0 ));
    InMux I__16548 (
            .O(N__72801),
            .I(N__72798));
    LocalMux I__16547 (
            .O(N__72798),
            .I(N__72794));
    InMux I__16546 (
            .O(N__72797),
            .I(N__72791));
    Span4Mux_v I__16545 (
            .O(N__72794),
            .I(N__72782));
    LocalMux I__16544 (
            .O(N__72791),
            .I(N__72779));
    InMux I__16543 (
            .O(N__72790),
            .I(N__72776));
    InMux I__16542 (
            .O(N__72789),
            .I(N__72773));
    InMux I__16541 (
            .O(N__72788),
            .I(N__72770));
    InMux I__16540 (
            .O(N__72787),
            .I(N__72766));
    InMux I__16539 (
            .O(N__72786),
            .I(N__72763));
    InMux I__16538 (
            .O(N__72785),
            .I(N__72760));
    Span4Mux_v I__16537 (
            .O(N__72782),
            .I(N__72757));
    Span4Mux_s2_h I__16536 (
            .O(N__72779),
            .I(N__72754));
    LocalMux I__16535 (
            .O(N__72776),
            .I(N__72747));
    LocalMux I__16534 (
            .O(N__72773),
            .I(N__72747));
    LocalMux I__16533 (
            .O(N__72770),
            .I(N__72747));
    InMux I__16532 (
            .O(N__72769),
            .I(N__72744));
    LocalMux I__16531 (
            .O(N__72766),
            .I(N__72737));
    LocalMux I__16530 (
            .O(N__72763),
            .I(N__72737));
    LocalMux I__16529 (
            .O(N__72760),
            .I(N__72737));
    Sp12to4 I__16528 (
            .O(N__72757),
            .I(N__72734));
    Span4Mux_h I__16527 (
            .O(N__72754),
            .I(N__72731));
    Span4Mux_v I__16526 (
            .O(N__72747),
            .I(N__72726));
    LocalMux I__16525 (
            .O(N__72744),
            .I(N__72726));
    Span4Mux_v I__16524 (
            .O(N__72737),
            .I(N__72723));
    Odrv12 I__16523 (
            .O(N__72734),
            .I(\pid_side.error_4 ));
    Odrv4 I__16522 (
            .O(N__72731),
            .I(\pid_side.error_4 ));
    Odrv4 I__16521 (
            .O(N__72726),
            .I(\pid_side.error_4 ));
    Odrv4 I__16520 (
            .O(N__72723),
            .I(\pid_side.error_4 ));
    InMux I__16519 (
            .O(N__72714),
            .I(N__72711));
    LocalMux I__16518 (
            .O(N__72711),
            .I(\pid_side.N_15_0_0 ));
    CascadeMux I__16517 (
            .O(N__72708),
            .I(N__72704));
    CascadeMux I__16516 (
            .O(N__72707),
            .I(N__72700));
    InMux I__16515 (
            .O(N__72704),
            .I(N__72692));
    InMux I__16514 (
            .O(N__72703),
            .I(N__72689));
    InMux I__16513 (
            .O(N__72700),
            .I(N__72686));
    CascadeMux I__16512 (
            .O(N__72699),
            .I(N__72683));
    CascadeMux I__16511 (
            .O(N__72698),
            .I(N__72680));
    InMux I__16510 (
            .O(N__72697),
            .I(N__72668));
    InMux I__16509 (
            .O(N__72696),
            .I(N__72668));
    InMux I__16508 (
            .O(N__72695),
            .I(N__72668));
    LocalMux I__16507 (
            .O(N__72692),
            .I(N__72665));
    LocalMux I__16506 (
            .O(N__72689),
            .I(N__72660));
    LocalMux I__16505 (
            .O(N__72686),
            .I(N__72657));
    InMux I__16504 (
            .O(N__72683),
            .I(N__72652));
    InMux I__16503 (
            .O(N__72680),
            .I(N__72652));
    InMux I__16502 (
            .O(N__72679),
            .I(N__72649));
    InMux I__16501 (
            .O(N__72678),
            .I(N__72644));
    InMux I__16500 (
            .O(N__72677),
            .I(N__72644));
    InMux I__16499 (
            .O(N__72676),
            .I(N__72639));
    InMux I__16498 (
            .O(N__72675),
            .I(N__72639));
    LocalMux I__16497 (
            .O(N__72668),
            .I(N__72634));
    Span4Mux_v I__16496 (
            .O(N__72665),
            .I(N__72634));
    InMux I__16495 (
            .O(N__72664),
            .I(N__72631));
    InMux I__16494 (
            .O(N__72663),
            .I(N__72628));
    Span4Mux_v I__16493 (
            .O(N__72660),
            .I(N__72621));
    Span4Mux_v I__16492 (
            .O(N__72657),
            .I(N__72621));
    LocalMux I__16491 (
            .O(N__72652),
            .I(N__72621));
    LocalMux I__16490 (
            .O(N__72649),
            .I(N__72616));
    LocalMux I__16489 (
            .O(N__72644),
            .I(N__72616));
    LocalMux I__16488 (
            .O(N__72639),
            .I(N__72613));
    Span4Mux_h I__16487 (
            .O(N__72634),
            .I(N__72608));
    LocalMux I__16486 (
            .O(N__72631),
            .I(N__72608));
    LocalMux I__16485 (
            .O(N__72628),
            .I(N__72605));
    Span4Mux_h I__16484 (
            .O(N__72621),
            .I(N__72598));
    Span4Mux_v I__16483 (
            .O(N__72616),
            .I(N__72598));
    Span4Mux_h I__16482 (
            .O(N__72613),
            .I(N__72598));
    Span4Mux_v I__16481 (
            .O(N__72608),
            .I(N__72595));
    Odrv4 I__16480 (
            .O(N__72605),
            .I(xy_ki_0_rep1));
    Odrv4 I__16479 (
            .O(N__72598),
            .I(xy_ki_0_rep1));
    Odrv4 I__16478 (
            .O(N__72595),
            .I(xy_ki_0_rep1));
    InMux I__16477 (
            .O(N__72588),
            .I(N__72585));
    LocalMux I__16476 (
            .O(N__72585),
            .I(N__72577));
    InMux I__16475 (
            .O(N__72584),
            .I(N__72574));
    InMux I__16474 (
            .O(N__72583),
            .I(N__72570));
    InMux I__16473 (
            .O(N__72582),
            .I(N__72566));
    InMux I__16472 (
            .O(N__72581),
            .I(N__72563));
    InMux I__16471 (
            .O(N__72580),
            .I(N__72560));
    Span4Mux_s2_h I__16470 (
            .O(N__72577),
            .I(N__72557));
    LocalMux I__16469 (
            .O(N__72574),
            .I(N__72554));
    InMux I__16468 (
            .O(N__72573),
            .I(N__72551));
    LocalMux I__16467 (
            .O(N__72570),
            .I(N__72548));
    InMux I__16466 (
            .O(N__72569),
            .I(N__72545));
    LocalMux I__16465 (
            .O(N__72566),
            .I(N__72538));
    LocalMux I__16464 (
            .O(N__72563),
            .I(N__72538));
    LocalMux I__16463 (
            .O(N__72560),
            .I(N__72538));
    Span4Mux_h I__16462 (
            .O(N__72557),
            .I(N__72535));
    Span12Mux_s7_h I__16461 (
            .O(N__72554),
            .I(N__72526));
    LocalMux I__16460 (
            .O(N__72551),
            .I(N__72526));
    Span12Mux_s6_v I__16459 (
            .O(N__72548),
            .I(N__72526));
    LocalMux I__16458 (
            .O(N__72545),
            .I(N__72526));
    Span4Mux_v I__16457 (
            .O(N__72538),
            .I(N__72523));
    Odrv4 I__16456 (
            .O(N__72535),
            .I(\pid_side.error_5 ));
    Odrv12 I__16455 (
            .O(N__72526),
            .I(\pid_side.error_5 ));
    Odrv4 I__16454 (
            .O(N__72523),
            .I(\pid_side.error_5 ));
    InMux I__16453 (
            .O(N__72516),
            .I(N__72513));
    LocalMux I__16452 (
            .O(N__72513),
            .I(N__72509));
    InMux I__16451 (
            .O(N__72512),
            .I(N__72506));
    Span4Mux_s2_h I__16450 (
            .O(N__72509),
            .I(N__72498));
    LocalMux I__16449 (
            .O(N__72506),
            .I(N__72495));
    InMux I__16448 (
            .O(N__72505),
            .I(N__72492));
    InMux I__16447 (
            .O(N__72504),
            .I(N__72489));
    InMux I__16446 (
            .O(N__72503),
            .I(N__72485));
    InMux I__16445 (
            .O(N__72502),
            .I(N__72482));
    InMux I__16444 (
            .O(N__72501),
            .I(N__72479));
    Span4Mux_v I__16443 (
            .O(N__72498),
            .I(N__72476));
    Span4Mux_s2_h I__16442 (
            .O(N__72495),
            .I(N__72473));
    LocalMux I__16441 (
            .O(N__72492),
            .I(N__72468));
    LocalMux I__16440 (
            .O(N__72489),
            .I(N__72468));
    InMux I__16439 (
            .O(N__72488),
            .I(N__72465));
    LocalMux I__16438 (
            .O(N__72485),
            .I(N__72458));
    LocalMux I__16437 (
            .O(N__72482),
            .I(N__72458));
    LocalMux I__16436 (
            .O(N__72479),
            .I(N__72458));
    Span4Mux_h I__16435 (
            .O(N__72476),
            .I(N__72455));
    Span4Mux_h I__16434 (
            .O(N__72473),
            .I(N__72452));
    Span4Mux_v I__16433 (
            .O(N__72468),
            .I(N__72447));
    LocalMux I__16432 (
            .O(N__72465),
            .I(N__72447));
    Span4Mux_v I__16431 (
            .O(N__72458),
            .I(N__72444));
    Odrv4 I__16430 (
            .O(N__72455),
            .I(\pid_side.error_6 ));
    Odrv4 I__16429 (
            .O(N__72452),
            .I(\pid_side.error_6 ));
    Odrv4 I__16428 (
            .O(N__72447),
            .I(\pid_side.error_6 ));
    Odrv4 I__16427 (
            .O(N__72444),
            .I(\pid_side.error_6 ));
    InMux I__16426 (
            .O(N__72435),
            .I(N__72432));
    LocalMux I__16425 (
            .O(N__72432),
            .I(N__72427));
    InMux I__16424 (
            .O(N__72431),
            .I(N__72422));
    CascadeMux I__16423 (
            .O(N__72430),
            .I(N__72418));
    Span4Mux_s0_h I__16422 (
            .O(N__72427),
            .I(N__72415));
    InMux I__16421 (
            .O(N__72426),
            .I(N__72412));
    InMux I__16420 (
            .O(N__72425),
            .I(N__72407));
    LocalMux I__16419 (
            .O(N__72422),
            .I(N__72404));
    InMux I__16418 (
            .O(N__72421),
            .I(N__72399));
    InMux I__16417 (
            .O(N__72418),
            .I(N__72399));
    Span4Mux_v I__16416 (
            .O(N__72415),
            .I(N__72396));
    LocalMux I__16415 (
            .O(N__72412),
            .I(N__72393));
    InMux I__16414 (
            .O(N__72411),
            .I(N__72390));
    InMux I__16413 (
            .O(N__72410),
            .I(N__72387));
    LocalMux I__16412 (
            .O(N__72407),
            .I(N__72384));
    Span4Mux_v I__16411 (
            .O(N__72404),
            .I(N__72381));
    LocalMux I__16410 (
            .O(N__72399),
            .I(N__72378));
    Span4Mux_v I__16409 (
            .O(N__72396),
            .I(N__72375));
    Span4Mux_h I__16408 (
            .O(N__72393),
            .I(N__72370));
    LocalMux I__16407 (
            .O(N__72390),
            .I(N__72370));
    LocalMux I__16406 (
            .O(N__72387),
            .I(N__72367));
    Span4Mux_h I__16405 (
            .O(N__72384),
            .I(N__72356));
    Span4Mux_h I__16404 (
            .O(N__72381),
            .I(N__72356));
    Span4Mux_v I__16403 (
            .O(N__72378),
            .I(N__72356));
    Span4Mux_h I__16402 (
            .O(N__72375),
            .I(N__72356));
    Span4Mux_v I__16401 (
            .O(N__72370),
            .I(N__72356));
    Odrv12 I__16400 (
            .O(N__72367),
            .I(\pid_side.error_8 ));
    Odrv4 I__16399 (
            .O(N__72356),
            .I(\pid_side.error_8 ));
    InMux I__16398 (
            .O(N__72351),
            .I(N__72348));
    LocalMux I__16397 (
            .O(N__72348),
            .I(N__72341));
    InMux I__16396 (
            .O(N__72347),
            .I(N__72338));
    InMux I__16395 (
            .O(N__72346),
            .I(N__72332));
    InMux I__16394 (
            .O(N__72345),
            .I(N__72329));
    InMux I__16393 (
            .O(N__72344),
            .I(N__72326));
    Span4Mux_v I__16392 (
            .O(N__72341),
            .I(N__72321));
    LocalMux I__16391 (
            .O(N__72338),
            .I(N__72321));
    InMux I__16390 (
            .O(N__72337),
            .I(N__72318));
    InMux I__16389 (
            .O(N__72336),
            .I(N__72315));
    InMux I__16388 (
            .O(N__72335),
            .I(N__72312));
    LocalMux I__16387 (
            .O(N__72332),
            .I(N__72307));
    LocalMux I__16386 (
            .O(N__72329),
            .I(N__72307));
    LocalMux I__16385 (
            .O(N__72326),
            .I(N__72304));
    Span4Mux_v I__16384 (
            .O(N__72321),
            .I(N__72301));
    LocalMux I__16383 (
            .O(N__72318),
            .I(N__72294));
    LocalMux I__16382 (
            .O(N__72315),
            .I(N__72294));
    LocalMux I__16381 (
            .O(N__72312),
            .I(N__72294));
    Span4Mux_v I__16380 (
            .O(N__72307),
            .I(N__72289));
    Span4Mux_h I__16379 (
            .O(N__72304),
            .I(N__72289));
    Span4Mux_h I__16378 (
            .O(N__72301),
            .I(N__72284));
    Span4Mux_v I__16377 (
            .O(N__72294),
            .I(N__72284));
    Odrv4 I__16376 (
            .O(N__72289),
            .I(\pid_side.error_7 ));
    Odrv4 I__16375 (
            .O(N__72284),
            .I(\pid_side.error_7 ));
    CascadeMux I__16374 (
            .O(N__72279),
            .I(\pid_side.g0_i_m4_1_cascade_ ));
    CascadeMux I__16373 (
            .O(N__72276),
            .I(N__72266));
    InMux I__16372 (
            .O(N__72275),
            .I(N__72261));
    InMux I__16371 (
            .O(N__72274),
            .I(N__72261));
    CascadeMux I__16370 (
            .O(N__72273),
            .I(N__72257));
    InMux I__16369 (
            .O(N__72272),
            .I(N__72254));
    CascadeMux I__16368 (
            .O(N__72271),
            .I(N__72250));
    CascadeMux I__16367 (
            .O(N__72270),
            .I(N__72247));
    CascadeMux I__16366 (
            .O(N__72269),
            .I(N__72241));
    InMux I__16365 (
            .O(N__72266),
            .I(N__72238));
    LocalMux I__16364 (
            .O(N__72261),
            .I(N__72235));
    InMux I__16363 (
            .O(N__72260),
            .I(N__72230));
    InMux I__16362 (
            .O(N__72257),
            .I(N__72230));
    LocalMux I__16361 (
            .O(N__72254),
            .I(N__72227));
    InMux I__16360 (
            .O(N__72253),
            .I(N__72222));
    InMux I__16359 (
            .O(N__72250),
            .I(N__72222));
    InMux I__16358 (
            .O(N__72247),
            .I(N__72215));
    InMux I__16357 (
            .O(N__72246),
            .I(N__72212));
    InMux I__16356 (
            .O(N__72245),
            .I(N__72204));
    InMux I__16355 (
            .O(N__72244),
            .I(N__72204));
    InMux I__16354 (
            .O(N__72241),
            .I(N__72201));
    LocalMux I__16353 (
            .O(N__72238),
            .I(N__72198));
    Span4Mux_v I__16352 (
            .O(N__72235),
            .I(N__72193));
    LocalMux I__16351 (
            .O(N__72230),
            .I(N__72193));
    Span4Mux_v I__16350 (
            .O(N__72227),
            .I(N__72188));
    LocalMux I__16349 (
            .O(N__72222),
            .I(N__72188));
    CascadeMux I__16348 (
            .O(N__72221),
            .I(N__72184));
    CascadeMux I__16347 (
            .O(N__72220),
            .I(N__72181));
    CascadeMux I__16346 (
            .O(N__72219),
            .I(N__72175));
    InMux I__16345 (
            .O(N__72218),
            .I(N__72172));
    LocalMux I__16344 (
            .O(N__72215),
            .I(N__72169));
    LocalMux I__16343 (
            .O(N__72212),
            .I(N__72166));
    InMux I__16342 (
            .O(N__72211),
            .I(N__72163));
    InMux I__16341 (
            .O(N__72210),
            .I(N__72160));
    InMux I__16340 (
            .O(N__72209),
            .I(N__72157));
    LocalMux I__16339 (
            .O(N__72204),
            .I(N__72152));
    LocalMux I__16338 (
            .O(N__72201),
            .I(N__72152));
    Span4Mux_h I__16337 (
            .O(N__72198),
            .I(N__72145));
    Span4Mux_v I__16336 (
            .O(N__72193),
            .I(N__72145));
    Span4Mux_v I__16335 (
            .O(N__72188),
            .I(N__72145));
    InMux I__16334 (
            .O(N__72187),
            .I(N__72140));
    InMux I__16333 (
            .O(N__72184),
            .I(N__72140));
    InMux I__16332 (
            .O(N__72181),
            .I(N__72137));
    InMux I__16331 (
            .O(N__72180),
            .I(N__72134));
    InMux I__16330 (
            .O(N__72179),
            .I(N__72127));
    InMux I__16329 (
            .O(N__72178),
            .I(N__72127));
    InMux I__16328 (
            .O(N__72175),
            .I(N__72127));
    LocalMux I__16327 (
            .O(N__72172),
            .I(xy_ki_1_rep2));
    Odrv4 I__16326 (
            .O(N__72169),
            .I(xy_ki_1_rep2));
    Odrv4 I__16325 (
            .O(N__72166),
            .I(xy_ki_1_rep2));
    LocalMux I__16324 (
            .O(N__72163),
            .I(xy_ki_1_rep2));
    LocalMux I__16323 (
            .O(N__72160),
            .I(xy_ki_1_rep2));
    LocalMux I__16322 (
            .O(N__72157),
            .I(xy_ki_1_rep2));
    Odrv4 I__16321 (
            .O(N__72152),
            .I(xy_ki_1_rep2));
    Odrv4 I__16320 (
            .O(N__72145),
            .I(xy_ki_1_rep2));
    LocalMux I__16319 (
            .O(N__72140),
            .I(xy_ki_1_rep2));
    LocalMux I__16318 (
            .O(N__72137),
            .I(xy_ki_1_rep2));
    LocalMux I__16317 (
            .O(N__72134),
            .I(xy_ki_1_rep2));
    LocalMux I__16316 (
            .O(N__72127),
            .I(xy_ki_1_rep2));
    InMux I__16315 (
            .O(N__72102),
            .I(N__72099));
    LocalMux I__16314 (
            .O(N__72099),
            .I(N__72096));
    Odrv4 I__16313 (
            .O(N__72096),
            .I(\pid_side.N_9_1 ));
    InMux I__16312 (
            .O(N__72093),
            .I(N__72089));
    InMux I__16311 (
            .O(N__72092),
            .I(N__72086));
    LocalMux I__16310 (
            .O(N__72089),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    LocalMux I__16309 (
            .O(N__72086),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    InMux I__16308 (
            .O(N__72081),
            .I(N__72078));
    LocalMux I__16307 (
            .O(N__72078),
            .I(N__72075));
    Odrv4 I__16306 (
            .O(N__72075),
            .I(drone_H_disp_side_i_8));
    CascadeMux I__16305 (
            .O(N__72072),
            .I(N__72067));
    InMux I__16304 (
            .O(N__72071),
            .I(N__72060));
    InMux I__16303 (
            .O(N__72070),
            .I(N__72060));
    InMux I__16302 (
            .O(N__72067),
            .I(N__72060));
    LocalMux I__16301 (
            .O(N__72060),
            .I(N__72057));
    Span4Mux_h I__16300 (
            .O(N__72057),
            .I(N__72051));
    InMux I__16299 (
            .O(N__72056),
            .I(N__72044));
    InMux I__16298 (
            .O(N__72055),
            .I(N__72044));
    InMux I__16297 (
            .O(N__72054),
            .I(N__72044));
    Span4Mux_h I__16296 (
            .O(N__72051),
            .I(N__72037));
    LocalMux I__16295 (
            .O(N__72044),
            .I(N__72037));
    InMux I__16294 (
            .O(N__72043),
            .I(N__72032));
    InMux I__16293 (
            .O(N__72042),
            .I(N__72032));
    Span4Mux_v I__16292 (
            .O(N__72037),
            .I(N__72029));
    LocalMux I__16291 (
            .O(N__72032),
            .I(N__72026));
    Span4Mux_v I__16290 (
            .O(N__72029),
            .I(N__72022));
    Span4Mux_v I__16289 (
            .O(N__72026),
            .I(N__72019));
    InMux I__16288 (
            .O(N__72025),
            .I(N__72016));
    Span4Mux_h I__16287 (
            .O(N__72022),
            .I(N__72013));
    Span4Mux_h I__16286 (
            .O(N__72019),
            .I(N__72008));
    LocalMux I__16285 (
            .O(N__72016),
            .I(N__72008));
    Span4Mux_h I__16284 (
            .O(N__72013),
            .I(N__72003));
    Span4Mux_h I__16283 (
            .O(N__72008),
            .I(N__72003));
    Odrv4 I__16282 (
            .O(N__72003),
            .I(uart_drone_data_0));
    InMux I__16281 (
            .O(N__72000),
            .I(N__71996));
    InMux I__16280 (
            .O(N__71999),
            .I(N__71993));
    LocalMux I__16279 (
            .O(N__71996),
            .I(N__71990));
    LocalMux I__16278 (
            .O(N__71993),
            .I(dron_frame_decoder_1_source_H_disp_side_fast_0));
    Odrv4 I__16277 (
            .O(N__71990),
            .I(dron_frame_decoder_1_source_H_disp_side_fast_0));
    CascadeMux I__16276 (
            .O(N__71985),
            .I(N__71980));
    CascadeMux I__16275 (
            .O(N__71984),
            .I(N__71973));
    InMux I__16274 (
            .O(N__71983),
            .I(N__71961));
    InMux I__16273 (
            .O(N__71980),
            .I(N__71961));
    InMux I__16272 (
            .O(N__71979),
            .I(N__71961));
    InMux I__16271 (
            .O(N__71978),
            .I(N__71961));
    InMux I__16270 (
            .O(N__71977),
            .I(N__71947));
    InMux I__16269 (
            .O(N__71976),
            .I(N__71947));
    InMux I__16268 (
            .O(N__71973),
            .I(N__71947));
    InMux I__16267 (
            .O(N__71972),
            .I(N__71947));
    CascadeMux I__16266 (
            .O(N__71971),
            .I(N__71943));
    CascadeMux I__16265 (
            .O(N__71970),
            .I(N__71940));
    LocalMux I__16264 (
            .O(N__71961),
            .I(N__71936));
    InMux I__16263 (
            .O(N__71960),
            .I(N__71927));
    InMux I__16262 (
            .O(N__71959),
            .I(N__71927));
    InMux I__16261 (
            .O(N__71958),
            .I(N__71927));
    InMux I__16260 (
            .O(N__71957),
            .I(N__71927));
    CascadeMux I__16259 (
            .O(N__71956),
            .I(N__71924));
    LocalMux I__16258 (
            .O(N__71947),
            .I(N__71921));
    InMux I__16257 (
            .O(N__71946),
            .I(N__71912));
    InMux I__16256 (
            .O(N__71943),
            .I(N__71912));
    InMux I__16255 (
            .O(N__71940),
            .I(N__71912));
    InMux I__16254 (
            .O(N__71939),
            .I(N__71912));
    Span4Mux_h I__16253 (
            .O(N__71936),
            .I(N__71908));
    LocalMux I__16252 (
            .O(N__71927),
            .I(N__71905));
    InMux I__16251 (
            .O(N__71924),
            .I(N__71902));
    Span4Mux_h I__16250 (
            .O(N__71921),
            .I(N__71897));
    LocalMux I__16249 (
            .O(N__71912),
            .I(N__71897));
    CascadeMux I__16248 (
            .O(N__71911),
            .I(N__71894));
    Span4Mux_v I__16247 (
            .O(N__71908),
            .I(N__71888));
    Span4Mux_h I__16246 (
            .O(N__71905),
            .I(N__71888));
    LocalMux I__16245 (
            .O(N__71902),
            .I(N__71885));
    Span4Mux_h I__16244 (
            .O(N__71897),
            .I(N__71882));
    InMux I__16243 (
            .O(N__71894),
            .I(N__71877));
    InMux I__16242 (
            .O(N__71893),
            .I(N__71877));
    Span4Mux_h I__16241 (
            .O(N__71888),
            .I(N__71872));
    Span4Mux_v I__16240 (
            .O(N__71885),
            .I(N__71867));
    Span4Mux_h I__16239 (
            .O(N__71882),
            .I(N__71867));
    LocalMux I__16238 (
            .O(N__71877),
            .I(N__71864));
    InMux I__16237 (
            .O(N__71876),
            .I(N__71859));
    InMux I__16236 (
            .O(N__71875),
            .I(N__71859));
    Span4Mux_h I__16235 (
            .O(N__71872),
            .I(N__71856));
    Span4Mux_v I__16234 (
            .O(N__71867),
            .I(N__71851));
    Span4Mux_v I__16233 (
            .O(N__71864),
            .I(N__71851));
    LocalMux I__16232 (
            .O(N__71859),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    Odrv4 I__16231 (
            .O(N__71856),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    Odrv4 I__16230 (
            .O(N__71851),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    CascadeMux I__16229 (
            .O(N__71844),
            .I(N__71839));
    CascadeMux I__16228 (
            .O(N__71843),
            .I(N__71834));
    CascadeMux I__16227 (
            .O(N__71842),
            .I(N__71830));
    InMux I__16226 (
            .O(N__71839),
            .I(N__71827));
    InMux I__16225 (
            .O(N__71838),
            .I(N__71824));
    InMux I__16224 (
            .O(N__71837),
            .I(N__71821));
    InMux I__16223 (
            .O(N__71834),
            .I(N__71818));
    InMux I__16222 (
            .O(N__71833),
            .I(N__71813));
    InMux I__16221 (
            .O(N__71830),
            .I(N__71813));
    LocalMux I__16220 (
            .O(N__71827),
            .I(N__71810));
    LocalMux I__16219 (
            .O(N__71824),
            .I(N__71805));
    LocalMux I__16218 (
            .O(N__71821),
            .I(N__71805));
    LocalMux I__16217 (
            .O(N__71818),
            .I(N__71802));
    LocalMux I__16216 (
            .O(N__71813),
            .I(N__71799));
    Span4Mux_h I__16215 (
            .O(N__71810),
            .I(N__71791));
    Span4Mux_h I__16214 (
            .O(N__71805),
            .I(N__71791));
    Span4Mux_h I__16213 (
            .O(N__71802),
            .I(N__71791));
    Span4Mux_h I__16212 (
            .O(N__71799),
            .I(N__71788));
    InMux I__16211 (
            .O(N__71798),
            .I(N__71785));
    Sp12to4 I__16210 (
            .O(N__71791),
            .I(N__71782));
    Span4Mux_h I__16209 (
            .O(N__71788),
            .I(N__71777));
    LocalMux I__16208 (
            .O(N__71785),
            .I(N__71777));
    Span12Mux_v I__16207 (
            .O(N__71782),
            .I(N__71774));
    Span4Mux_v I__16206 (
            .O(N__71777),
            .I(N__71771));
    Odrv12 I__16205 (
            .O(N__71774),
            .I(uart_drone_data_2));
    Odrv4 I__16204 (
            .O(N__71771),
            .I(uart_drone_data_2));
    CascadeMux I__16203 (
            .O(N__71766),
            .I(N__71762));
    CascadeMux I__16202 (
            .O(N__71765),
            .I(N__71757));
    InMux I__16201 (
            .O(N__71762),
            .I(N__71742));
    InMux I__16200 (
            .O(N__71761),
            .I(N__71742));
    InMux I__16199 (
            .O(N__71760),
            .I(N__71742));
    InMux I__16198 (
            .O(N__71757),
            .I(N__71742));
    InMux I__16197 (
            .O(N__71756),
            .I(N__71733));
    InMux I__16196 (
            .O(N__71755),
            .I(N__71733));
    InMux I__16195 (
            .O(N__71754),
            .I(N__71733));
    InMux I__16194 (
            .O(N__71753),
            .I(N__71733));
    CascadeMux I__16193 (
            .O(N__71752),
            .I(N__71730));
    CascadeMux I__16192 (
            .O(N__71751),
            .I(N__71725));
    LocalMux I__16191 (
            .O(N__71742),
            .I(N__71721));
    LocalMux I__16190 (
            .O(N__71733),
            .I(N__71718));
    InMux I__16189 (
            .O(N__71730),
            .I(N__71709));
    InMux I__16188 (
            .O(N__71729),
            .I(N__71709));
    InMux I__16187 (
            .O(N__71728),
            .I(N__71709));
    InMux I__16186 (
            .O(N__71725),
            .I(N__71709));
    InMux I__16185 (
            .O(N__71724),
            .I(N__71706));
    Span4Mux_v I__16184 (
            .O(N__71721),
            .I(N__71699));
    Span4Mux_v I__16183 (
            .O(N__71718),
            .I(N__71699));
    LocalMux I__16182 (
            .O(N__71709),
            .I(N__71699));
    LocalMux I__16181 (
            .O(N__71706),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_1_0 ));
    Odrv4 I__16180 (
            .O(N__71699),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_1_0 ));
    InMux I__16179 (
            .O(N__71694),
            .I(N__71688));
    InMux I__16178 (
            .O(N__71693),
            .I(N__71688));
    LocalMux I__16177 (
            .O(N__71688),
            .I(\dron_frame_decoder_1.drone_H_disp_side_10 ));
    InMux I__16176 (
            .O(N__71685),
            .I(N__71682));
    LocalMux I__16175 (
            .O(N__71682),
            .I(N__71679));
    Odrv4 I__16174 (
            .O(N__71679),
            .I(drone_H_disp_side_i_10));
    InMux I__16173 (
            .O(N__71676),
            .I(N__71672));
    InMux I__16172 (
            .O(N__71675),
            .I(N__71665));
    LocalMux I__16171 (
            .O(N__71672),
            .I(N__71662));
    InMux I__16170 (
            .O(N__71671),
            .I(N__71654));
    InMux I__16169 (
            .O(N__71670),
            .I(N__71654));
    CascadeMux I__16168 (
            .O(N__71669),
            .I(N__71651));
    InMux I__16167 (
            .O(N__71668),
            .I(N__71648));
    LocalMux I__16166 (
            .O(N__71665),
            .I(N__71645));
    Span4Mux_s2_h I__16165 (
            .O(N__71662),
            .I(N__71642));
    InMux I__16164 (
            .O(N__71661),
            .I(N__71637));
    InMux I__16163 (
            .O(N__71660),
            .I(N__71637));
    InMux I__16162 (
            .O(N__71659),
            .I(N__71634));
    LocalMux I__16161 (
            .O(N__71654),
            .I(N__71631));
    InMux I__16160 (
            .O(N__71651),
            .I(N__71628));
    LocalMux I__16159 (
            .O(N__71648),
            .I(N__71625));
    Span4Mux_s2_h I__16158 (
            .O(N__71645),
            .I(N__71622));
    Span4Mux_v I__16157 (
            .O(N__71642),
            .I(N__71619));
    LocalMux I__16156 (
            .O(N__71637),
            .I(N__71610));
    LocalMux I__16155 (
            .O(N__71634),
            .I(N__71610));
    Span4Mux_h I__16154 (
            .O(N__71631),
            .I(N__71610));
    LocalMux I__16153 (
            .O(N__71628),
            .I(N__71610));
    Span4Mux_h I__16152 (
            .O(N__71625),
            .I(N__71605));
    Span4Mux_h I__16151 (
            .O(N__71622),
            .I(N__71605));
    Span4Mux_h I__16150 (
            .O(N__71619),
            .I(N__71602));
    Span4Mux_v I__16149 (
            .O(N__71610),
            .I(N__71599));
    Odrv4 I__16148 (
            .O(N__71605),
            .I(\pid_side.error_1 ));
    Odrv4 I__16147 (
            .O(N__71602),
            .I(\pid_side.error_1 ));
    Odrv4 I__16146 (
            .O(N__71599),
            .I(\pid_side.error_1 ));
    InMux I__16145 (
            .O(N__71592),
            .I(N__71589));
    LocalMux I__16144 (
            .O(N__71589),
            .I(\pid_side.N_12_1_0 ));
    InMux I__16143 (
            .O(N__71586),
            .I(N__71579));
    InMux I__16142 (
            .O(N__71585),
            .I(N__71574));
    InMux I__16141 (
            .O(N__71584),
            .I(N__71571));
    InMux I__16140 (
            .O(N__71583),
            .I(N__71566));
    InMux I__16139 (
            .O(N__71582),
            .I(N__71566));
    LocalMux I__16138 (
            .O(N__71579),
            .I(N__71563));
    InMux I__16137 (
            .O(N__71578),
            .I(N__71560));
    CascadeMux I__16136 (
            .O(N__71577),
            .I(N__71554));
    LocalMux I__16135 (
            .O(N__71574),
            .I(N__71549));
    LocalMux I__16134 (
            .O(N__71571),
            .I(N__71546));
    LocalMux I__16133 (
            .O(N__71566),
            .I(N__71543));
    Span4Mux_v I__16132 (
            .O(N__71563),
            .I(N__71538));
    LocalMux I__16131 (
            .O(N__71560),
            .I(N__71535));
    InMux I__16130 (
            .O(N__71559),
            .I(N__71532));
    InMux I__16129 (
            .O(N__71558),
            .I(N__71527));
    InMux I__16128 (
            .O(N__71557),
            .I(N__71527));
    InMux I__16127 (
            .O(N__71554),
            .I(N__71518));
    InMux I__16126 (
            .O(N__71553),
            .I(N__71518));
    InMux I__16125 (
            .O(N__71552),
            .I(N__71518));
    Span4Mux_v I__16124 (
            .O(N__71549),
            .I(N__71511));
    Span4Mux_v I__16123 (
            .O(N__71546),
            .I(N__71511));
    Span4Mux_v I__16122 (
            .O(N__71543),
            .I(N__71511));
    InMux I__16121 (
            .O(N__71542),
            .I(N__71508));
    InMux I__16120 (
            .O(N__71541),
            .I(N__71505));
    Span4Mux_h I__16119 (
            .O(N__71538),
            .I(N__71496));
    Span4Mux_v I__16118 (
            .O(N__71535),
            .I(N__71496));
    LocalMux I__16117 (
            .O(N__71532),
            .I(N__71496));
    LocalMux I__16116 (
            .O(N__71527),
            .I(N__71496));
    InMux I__16115 (
            .O(N__71526),
            .I(N__71491));
    InMux I__16114 (
            .O(N__71525),
            .I(N__71491));
    LocalMux I__16113 (
            .O(N__71518),
            .I(N__71488));
    Span4Mux_h I__16112 (
            .O(N__71511),
            .I(N__71485));
    LocalMux I__16111 (
            .O(N__71508),
            .I(N__71476));
    LocalMux I__16110 (
            .O(N__71505),
            .I(N__71476));
    Span4Mux_h I__16109 (
            .O(N__71496),
            .I(N__71476));
    LocalMux I__16108 (
            .O(N__71491),
            .I(N__71476));
    Odrv4 I__16107 (
            .O(N__71488),
            .I(xy_ki_0_rep2));
    Odrv4 I__16106 (
            .O(N__71485),
            .I(xy_ki_0_rep2));
    Odrv4 I__16105 (
            .O(N__71476),
            .I(xy_ki_0_rep2));
    CascadeMux I__16104 (
            .O(N__71469),
            .I(N__71464));
    CascadeMux I__16103 (
            .O(N__71468),
            .I(N__71458));
    CascadeMux I__16102 (
            .O(N__71467),
            .I(N__71455));
    InMux I__16101 (
            .O(N__71464),
            .I(N__71444));
    InMux I__16100 (
            .O(N__71463),
            .I(N__71437));
    InMux I__16099 (
            .O(N__71462),
            .I(N__71437));
    InMux I__16098 (
            .O(N__71461),
            .I(N__71437));
    InMux I__16097 (
            .O(N__71458),
            .I(N__71434));
    InMux I__16096 (
            .O(N__71455),
            .I(N__71431));
    InMux I__16095 (
            .O(N__71454),
            .I(N__71428));
    InMux I__16094 (
            .O(N__71453),
            .I(N__71423));
    InMux I__16093 (
            .O(N__71452),
            .I(N__71423));
    InMux I__16092 (
            .O(N__71451),
            .I(N__71420));
    InMux I__16091 (
            .O(N__71450),
            .I(N__71417));
    InMux I__16090 (
            .O(N__71449),
            .I(N__71412));
    InMux I__16089 (
            .O(N__71448),
            .I(N__71412));
    InMux I__16088 (
            .O(N__71447),
            .I(N__71409));
    LocalMux I__16087 (
            .O(N__71444),
            .I(N__71404));
    LocalMux I__16086 (
            .O(N__71437),
            .I(N__71404));
    LocalMux I__16085 (
            .O(N__71434),
            .I(N__71399));
    LocalMux I__16084 (
            .O(N__71431),
            .I(N__71399));
    LocalMux I__16083 (
            .O(N__71428),
            .I(N__71394));
    LocalMux I__16082 (
            .O(N__71423),
            .I(N__71389));
    LocalMux I__16081 (
            .O(N__71420),
            .I(N__71389));
    LocalMux I__16080 (
            .O(N__71417),
            .I(N__71384));
    LocalMux I__16079 (
            .O(N__71412),
            .I(N__71384));
    LocalMux I__16078 (
            .O(N__71409),
            .I(N__71381));
    Span4Mux_v I__16077 (
            .O(N__71404),
            .I(N__71376));
    Span4Mux_v I__16076 (
            .O(N__71399),
            .I(N__71376));
    InMux I__16075 (
            .O(N__71398),
            .I(N__71371));
    InMux I__16074 (
            .O(N__71397),
            .I(N__71371));
    Span4Mux_h I__16073 (
            .O(N__71394),
            .I(N__71368));
    Span4Mux_h I__16072 (
            .O(N__71389),
            .I(N__71365));
    Span4Mux_v I__16071 (
            .O(N__71384),
            .I(N__71360));
    Span4Mux_h I__16070 (
            .O(N__71381),
            .I(N__71360));
    Span4Mux_h I__16069 (
            .O(N__71376),
            .I(N__71357));
    LocalMux I__16068 (
            .O(N__71371),
            .I(N__71354));
    Span4Mux_h I__16067 (
            .O(N__71368),
            .I(N__71349));
    Span4Mux_h I__16066 (
            .O(N__71365),
            .I(N__71349));
    Span4Mux_h I__16065 (
            .O(N__71360),
            .I(N__71346));
    Odrv4 I__16064 (
            .O(N__71357),
            .I(xy_ki_fast_0));
    Odrv12 I__16063 (
            .O(N__71354),
            .I(xy_ki_fast_0));
    Odrv4 I__16062 (
            .O(N__71349),
            .I(xy_ki_fast_0));
    Odrv4 I__16061 (
            .O(N__71346),
            .I(xy_ki_fast_0));
    InMux I__16060 (
            .O(N__71337),
            .I(N__71334));
    LocalMux I__16059 (
            .O(N__71334),
            .I(\pid_side.m87_0_ns_1 ));
    InMux I__16058 (
            .O(N__71331),
            .I(N__71327));
    InMux I__16057 (
            .O(N__71330),
            .I(N__71323));
    LocalMux I__16056 (
            .O(N__71327),
            .I(N__71320));
    InMux I__16055 (
            .O(N__71326),
            .I(N__71317));
    LocalMux I__16054 (
            .O(N__71323),
            .I(N__71314));
    Span4Mux_s2_h I__16053 (
            .O(N__71320),
            .I(N__71311));
    LocalMux I__16052 (
            .O(N__71317),
            .I(N__71305));
    Span4Mux_s2_h I__16051 (
            .O(N__71314),
            .I(N__71299));
    Span4Mux_v I__16050 (
            .O(N__71311),
            .I(N__71296));
    InMux I__16049 (
            .O(N__71310),
            .I(N__71291));
    InMux I__16048 (
            .O(N__71309),
            .I(N__71291));
    InMux I__16047 (
            .O(N__71308),
            .I(N__71288));
    Span4Mux_v I__16046 (
            .O(N__71305),
            .I(N__71285));
    InMux I__16045 (
            .O(N__71304),
            .I(N__71282));
    InMux I__16044 (
            .O(N__71303),
            .I(N__71277));
    InMux I__16043 (
            .O(N__71302),
            .I(N__71277));
    Span4Mux_h I__16042 (
            .O(N__71299),
            .I(N__71274));
    Span4Mux_h I__16041 (
            .O(N__71296),
            .I(N__71271));
    LocalMux I__16040 (
            .O(N__71291),
            .I(N__71268));
    LocalMux I__16039 (
            .O(N__71288),
            .I(\pid_side.error_10 ));
    Odrv4 I__16038 (
            .O(N__71285),
            .I(\pid_side.error_10 ));
    LocalMux I__16037 (
            .O(N__71282),
            .I(\pid_side.error_10 ));
    LocalMux I__16036 (
            .O(N__71277),
            .I(\pid_side.error_10 ));
    Odrv4 I__16035 (
            .O(N__71274),
            .I(\pid_side.error_10 ));
    Odrv4 I__16034 (
            .O(N__71271),
            .I(\pid_side.error_10 ));
    Odrv4 I__16033 (
            .O(N__71268),
            .I(\pid_side.error_10 ));
    CascadeMux I__16032 (
            .O(N__71253),
            .I(\pid_side.m87_0_ns_1_0_cascade_ ));
    InMux I__16031 (
            .O(N__71250),
            .I(N__71247));
    LocalMux I__16030 (
            .O(N__71247),
            .I(N__71244));
    Odrv4 I__16029 (
            .O(N__71244),
            .I(\pid_side.N_88_0_0 ));
    InMux I__16028 (
            .O(N__71241),
            .I(N__71237));
    InMux I__16027 (
            .O(N__71240),
            .I(N__71233));
    LocalMux I__16026 (
            .O(N__71237),
            .I(N__71230));
    InMux I__16025 (
            .O(N__71236),
            .I(N__71227));
    LocalMux I__16024 (
            .O(N__71233),
            .I(N__71224));
    Span4Mux_s3_h I__16023 (
            .O(N__71230),
            .I(N__71220));
    LocalMux I__16022 (
            .O(N__71227),
            .I(N__71217));
    Span4Mux_s2_h I__16021 (
            .O(N__71224),
            .I(N__71213));
    InMux I__16020 (
            .O(N__71223),
            .I(N__71209));
    Span4Mux_v I__16019 (
            .O(N__71220),
            .I(N__71206));
    Span4Mux_v I__16018 (
            .O(N__71217),
            .I(N__71203));
    CascadeMux I__16017 (
            .O(N__71216),
            .I(N__71200));
    Span4Mux_h I__16016 (
            .O(N__71213),
            .I(N__71195));
    InMux I__16015 (
            .O(N__71212),
            .I(N__71192));
    LocalMux I__16014 (
            .O(N__71209),
            .I(N__71189));
    Span4Mux_v I__16013 (
            .O(N__71206),
            .I(N__71184));
    Span4Mux_h I__16012 (
            .O(N__71203),
            .I(N__71184));
    InMux I__16011 (
            .O(N__71200),
            .I(N__71177));
    InMux I__16010 (
            .O(N__71199),
            .I(N__71177));
    InMux I__16009 (
            .O(N__71198),
            .I(N__71177));
    Odrv4 I__16008 (
            .O(N__71195),
            .I(\pid_side.error_11 ));
    LocalMux I__16007 (
            .O(N__71192),
            .I(\pid_side.error_11 ));
    Odrv4 I__16006 (
            .O(N__71189),
            .I(\pid_side.error_11 ));
    Odrv4 I__16005 (
            .O(N__71184),
            .I(\pid_side.error_11 ));
    LocalMux I__16004 (
            .O(N__71177),
            .I(\pid_side.error_11 ));
    InMux I__16003 (
            .O(N__71166),
            .I(N__71162));
    CascadeMux I__16002 (
            .O(N__71165),
            .I(N__71157));
    LocalMux I__16001 (
            .O(N__71162),
            .I(N__71151));
    CascadeMux I__16000 (
            .O(N__71161),
            .I(N__71143));
    InMux I__15999 (
            .O(N__71160),
            .I(N__71140));
    InMux I__15998 (
            .O(N__71157),
            .I(N__71137));
    InMux I__15997 (
            .O(N__71156),
            .I(N__71134));
    InMux I__15996 (
            .O(N__71155),
            .I(N__71131));
    InMux I__15995 (
            .O(N__71154),
            .I(N__71128));
    Span4Mux_h I__15994 (
            .O(N__71151),
            .I(N__71124));
    CascadeMux I__15993 (
            .O(N__71150),
            .I(N__71121));
    InMux I__15992 (
            .O(N__71149),
            .I(N__71118));
    CascadeMux I__15991 (
            .O(N__71148),
            .I(N__71113));
    InMux I__15990 (
            .O(N__71147),
            .I(N__71110));
    InMux I__15989 (
            .O(N__71146),
            .I(N__71104));
    InMux I__15988 (
            .O(N__71143),
            .I(N__71104));
    LocalMux I__15987 (
            .O(N__71140),
            .I(N__71101));
    LocalMux I__15986 (
            .O(N__71137),
            .I(N__71098));
    LocalMux I__15985 (
            .O(N__71134),
            .I(N__71093));
    LocalMux I__15984 (
            .O(N__71131),
            .I(N__71093));
    LocalMux I__15983 (
            .O(N__71128),
            .I(N__71090));
    InMux I__15982 (
            .O(N__71127),
            .I(N__71086));
    Span4Mux_v I__15981 (
            .O(N__71124),
            .I(N__71083));
    InMux I__15980 (
            .O(N__71121),
            .I(N__71080));
    LocalMux I__15979 (
            .O(N__71118),
            .I(N__71077));
    InMux I__15978 (
            .O(N__71117),
            .I(N__71071));
    InMux I__15977 (
            .O(N__71116),
            .I(N__71071));
    InMux I__15976 (
            .O(N__71113),
            .I(N__71068));
    LocalMux I__15975 (
            .O(N__71110),
            .I(N__71065));
    CascadeMux I__15974 (
            .O(N__71109),
            .I(N__71061));
    LocalMux I__15973 (
            .O(N__71104),
            .I(N__71056));
    Span4Mux_v I__15972 (
            .O(N__71101),
            .I(N__71047));
    Span4Mux_v I__15971 (
            .O(N__71098),
            .I(N__71047));
    Span4Mux_v I__15970 (
            .O(N__71093),
            .I(N__71047));
    Span4Mux_v I__15969 (
            .O(N__71090),
            .I(N__71047));
    InMux I__15968 (
            .O(N__71089),
            .I(N__71044));
    LocalMux I__15967 (
            .O(N__71086),
            .I(N__71035));
    Span4Mux_v I__15966 (
            .O(N__71083),
            .I(N__71035));
    LocalMux I__15965 (
            .O(N__71080),
            .I(N__71035));
    Span4Mux_v I__15964 (
            .O(N__71077),
            .I(N__71035));
    InMux I__15963 (
            .O(N__71076),
            .I(N__71032));
    LocalMux I__15962 (
            .O(N__71071),
            .I(N__71029));
    LocalMux I__15961 (
            .O(N__71068),
            .I(N__71024));
    Span4Mux_h I__15960 (
            .O(N__71065),
            .I(N__71024));
    InMux I__15959 (
            .O(N__71064),
            .I(N__71019));
    InMux I__15958 (
            .O(N__71061),
            .I(N__71019));
    InMux I__15957 (
            .O(N__71060),
            .I(N__71014));
    InMux I__15956 (
            .O(N__71059),
            .I(N__71014));
    Span4Mux_v I__15955 (
            .O(N__71056),
            .I(N__71009));
    Span4Mux_h I__15954 (
            .O(N__71047),
            .I(N__71009));
    LocalMux I__15953 (
            .O(N__71044),
            .I(xy_ki_0));
    Odrv4 I__15952 (
            .O(N__71035),
            .I(xy_ki_0));
    LocalMux I__15951 (
            .O(N__71032),
            .I(xy_ki_0));
    Odrv12 I__15950 (
            .O(N__71029),
            .I(xy_ki_0));
    Odrv4 I__15949 (
            .O(N__71024),
            .I(xy_ki_0));
    LocalMux I__15948 (
            .O(N__71019),
            .I(xy_ki_0));
    LocalMux I__15947 (
            .O(N__71014),
            .I(xy_ki_0));
    Odrv4 I__15946 (
            .O(N__71009),
            .I(xy_ki_0));
    InMux I__15945 (
            .O(N__70992),
            .I(N__70989));
    LocalMux I__15944 (
            .O(N__70989),
            .I(N__70985));
    InMux I__15943 (
            .O(N__70988),
            .I(N__70981));
    Span4Mux_v I__15942 (
            .O(N__70985),
            .I(N__70978));
    InMux I__15941 (
            .O(N__70984),
            .I(N__70974));
    LocalMux I__15940 (
            .O(N__70981),
            .I(N__70971));
    Span4Mux_s0_h I__15939 (
            .O(N__70978),
            .I(N__70968));
    InMux I__15938 (
            .O(N__70977),
            .I(N__70963));
    LocalMux I__15937 (
            .O(N__70974),
            .I(N__70958));
    Span12Mux_s7_h I__15936 (
            .O(N__70971),
            .I(N__70955));
    Sp12to4 I__15935 (
            .O(N__70968),
            .I(N__70952));
    InMux I__15934 (
            .O(N__70967),
            .I(N__70949));
    InMux I__15933 (
            .O(N__70966),
            .I(N__70946));
    LocalMux I__15932 (
            .O(N__70963),
            .I(N__70943));
    InMux I__15931 (
            .O(N__70962),
            .I(N__70938));
    InMux I__15930 (
            .O(N__70961),
            .I(N__70938));
    Span4Mux_h I__15929 (
            .O(N__70958),
            .I(N__70935));
    Odrv12 I__15928 (
            .O(N__70955),
            .I(\pid_side.error_12 ));
    Odrv12 I__15927 (
            .O(N__70952),
            .I(\pid_side.error_12 ));
    LocalMux I__15926 (
            .O(N__70949),
            .I(\pid_side.error_12 ));
    LocalMux I__15925 (
            .O(N__70946),
            .I(\pid_side.error_12 ));
    Odrv4 I__15924 (
            .O(N__70943),
            .I(\pid_side.error_12 ));
    LocalMux I__15923 (
            .O(N__70938),
            .I(\pid_side.error_12 ));
    Odrv4 I__15922 (
            .O(N__70935),
            .I(\pid_side.error_12 ));
    InMux I__15921 (
            .O(N__70920),
            .I(N__70916));
    InMux I__15920 (
            .O(N__70919),
            .I(N__70911));
    LocalMux I__15919 (
            .O(N__70916),
            .I(N__70908));
    InMux I__15918 (
            .O(N__70915),
            .I(N__70904));
    CascadeMux I__15917 (
            .O(N__70914),
            .I(N__70901));
    LocalMux I__15916 (
            .O(N__70911),
            .I(N__70898));
    Span4Mux_s2_h I__15915 (
            .O(N__70908),
            .I(N__70895));
    InMux I__15914 (
            .O(N__70907),
            .I(N__70889));
    LocalMux I__15913 (
            .O(N__70904),
            .I(N__70886));
    InMux I__15912 (
            .O(N__70901),
            .I(N__70883));
    Span4Mux_v I__15911 (
            .O(N__70898),
            .I(N__70880));
    Span4Mux_v I__15910 (
            .O(N__70895),
            .I(N__70877));
    InMux I__15909 (
            .O(N__70894),
            .I(N__70874));
    InMux I__15908 (
            .O(N__70893),
            .I(N__70869));
    InMux I__15907 (
            .O(N__70892),
            .I(N__70869));
    LocalMux I__15906 (
            .O(N__70889),
            .I(N__70866));
    Span4Mux_v I__15905 (
            .O(N__70886),
            .I(N__70863));
    LocalMux I__15904 (
            .O(N__70883),
            .I(N__70858));
    Sp12to4 I__15903 (
            .O(N__70880),
            .I(N__70858));
    Span4Mux_h I__15902 (
            .O(N__70877),
            .I(N__70855));
    LocalMux I__15901 (
            .O(N__70874),
            .I(\pid_side.error_13 ));
    LocalMux I__15900 (
            .O(N__70869),
            .I(\pid_side.error_13 ));
    Odrv4 I__15899 (
            .O(N__70866),
            .I(\pid_side.error_13 ));
    Odrv4 I__15898 (
            .O(N__70863),
            .I(\pid_side.error_13 ));
    Odrv12 I__15897 (
            .O(N__70858),
            .I(\pid_side.error_13 ));
    Odrv4 I__15896 (
            .O(N__70855),
            .I(\pid_side.error_13 ));
    CascadeMux I__15895 (
            .O(N__70842),
            .I(\pid_side.m36_1_ns_1_cascade_ ));
    InMux I__15894 (
            .O(N__70839),
            .I(N__70836));
    LocalMux I__15893 (
            .O(N__70836),
            .I(N__70833));
    Span4Mux_s0_h I__15892 (
            .O(N__70833),
            .I(N__70829));
    InMux I__15891 (
            .O(N__70832),
            .I(N__70826));
    Span4Mux_v I__15890 (
            .O(N__70829),
            .I(N__70818));
    LocalMux I__15889 (
            .O(N__70826),
            .I(N__70818));
    InMux I__15888 (
            .O(N__70825),
            .I(N__70815));
    InMux I__15887 (
            .O(N__70824),
            .I(N__70810));
    InMux I__15886 (
            .O(N__70823),
            .I(N__70810));
    Span4Mux_v I__15885 (
            .O(N__70818),
            .I(N__70804));
    LocalMux I__15884 (
            .O(N__70815),
            .I(N__70801));
    LocalMux I__15883 (
            .O(N__70810),
            .I(N__70798));
    InMux I__15882 (
            .O(N__70809),
            .I(N__70795));
    InMux I__15881 (
            .O(N__70808),
            .I(N__70792));
    InMux I__15880 (
            .O(N__70807),
            .I(N__70789));
    Span4Mux_h I__15879 (
            .O(N__70804),
            .I(N__70782));
    Span4Mux_h I__15878 (
            .O(N__70801),
            .I(N__70782));
    Span4Mux_v I__15877 (
            .O(N__70798),
            .I(N__70782));
    LocalMux I__15876 (
            .O(N__70795),
            .I(\pid_side.error_14 ));
    LocalMux I__15875 (
            .O(N__70792),
            .I(\pid_side.error_14 ));
    LocalMux I__15874 (
            .O(N__70789),
            .I(\pid_side.error_14 ));
    Odrv4 I__15873 (
            .O(N__70782),
            .I(\pid_side.error_14 ));
    InMux I__15872 (
            .O(N__70773),
            .I(N__70770));
    LocalMux I__15871 (
            .O(N__70770),
            .I(N__70766));
    InMux I__15870 (
            .O(N__70769),
            .I(N__70763));
    Span4Mux_v I__15869 (
            .O(N__70766),
            .I(N__70758));
    LocalMux I__15868 (
            .O(N__70763),
            .I(N__70758));
    Odrv4 I__15867 (
            .O(N__70758),
            .I(\pid_side.N_37_1 ));
    CascadeMux I__15866 (
            .O(N__70755),
            .I(N__70752));
    InMux I__15865 (
            .O(N__70752),
            .I(N__70749));
    LocalMux I__15864 (
            .O(N__70749),
            .I(N__70743));
    InMux I__15863 (
            .O(N__70748),
            .I(N__70738));
    InMux I__15862 (
            .O(N__70747),
            .I(N__70734));
    CascadeMux I__15861 (
            .O(N__70746),
            .I(N__70728));
    Span4Mux_v I__15860 (
            .O(N__70743),
            .I(N__70725));
    InMux I__15859 (
            .O(N__70742),
            .I(N__70722));
    InMux I__15858 (
            .O(N__70741),
            .I(N__70719));
    LocalMux I__15857 (
            .O(N__70738),
            .I(N__70716));
    InMux I__15856 (
            .O(N__70737),
            .I(N__70713));
    LocalMux I__15855 (
            .O(N__70734),
            .I(N__70710));
    InMux I__15854 (
            .O(N__70733),
            .I(N__70707));
    CascadeMux I__15853 (
            .O(N__70732),
            .I(N__70699));
    InMux I__15852 (
            .O(N__70731),
            .I(N__70693));
    InMux I__15851 (
            .O(N__70728),
            .I(N__70690));
    Span4Mux_v I__15850 (
            .O(N__70725),
            .I(N__70687));
    LocalMux I__15849 (
            .O(N__70722),
            .I(N__70684));
    LocalMux I__15848 (
            .O(N__70719),
            .I(N__70673));
    Span4Mux_h I__15847 (
            .O(N__70716),
            .I(N__70673));
    LocalMux I__15846 (
            .O(N__70713),
            .I(N__70673));
    Span4Mux_v I__15845 (
            .O(N__70710),
            .I(N__70673));
    LocalMux I__15844 (
            .O(N__70707),
            .I(N__70673));
    InMux I__15843 (
            .O(N__70706),
            .I(N__70670));
    InMux I__15842 (
            .O(N__70705),
            .I(N__70667));
    InMux I__15841 (
            .O(N__70704),
            .I(N__70664));
    InMux I__15840 (
            .O(N__70703),
            .I(N__70661));
    InMux I__15839 (
            .O(N__70702),
            .I(N__70657));
    InMux I__15838 (
            .O(N__70699),
            .I(N__70651));
    InMux I__15837 (
            .O(N__70698),
            .I(N__70651));
    InMux I__15836 (
            .O(N__70697),
            .I(N__70648));
    CascadeMux I__15835 (
            .O(N__70696),
            .I(N__70640));
    LocalMux I__15834 (
            .O(N__70693),
            .I(N__70629));
    LocalMux I__15833 (
            .O(N__70690),
            .I(N__70629));
    Span4Mux_v I__15832 (
            .O(N__70687),
            .I(N__70629));
    Span4Mux_h I__15831 (
            .O(N__70684),
            .I(N__70629));
    Span4Mux_v I__15830 (
            .O(N__70673),
            .I(N__70626));
    LocalMux I__15829 (
            .O(N__70670),
            .I(N__70617));
    LocalMux I__15828 (
            .O(N__70667),
            .I(N__70617));
    LocalMux I__15827 (
            .O(N__70664),
            .I(N__70617));
    LocalMux I__15826 (
            .O(N__70661),
            .I(N__70617));
    InMux I__15825 (
            .O(N__70660),
            .I(N__70611));
    LocalMux I__15824 (
            .O(N__70657),
            .I(N__70608));
    InMux I__15823 (
            .O(N__70656),
            .I(N__70605));
    LocalMux I__15822 (
            .O(N__70651),
            .I(N__70600));
    LocalMux I__15821 (
            .O(N__70648),
            .I(N__70600));
    InMux I__15820 (
            .O(N__70647),
            .I(N__70595));
    InMux I__15819 (
            .O(N__70646),
            .I(N__70595));
    InMux I__15818 (
            .O(N__70645),
            .I(N__70586));
    InMux I__15817 (
            .O(N__70644),
            .I(N__70586));
    InMux I__15816 (
            .O(N__70643),
            .I(N__70586));
    InMux I__15815 (
            .O(N__70640),
            .I(N__70586));
    InMux I__15814 (
            .O(N__70639),
            .I(N__70583));
    InMux I__15813 (
            .O(N__70638),
            .I(N__70580));
    Span4Mux_v I__15812 (
            .O(N__70629),
            .I(N__70577));
    Span4Mux_h I__15811 (
            .O(N__70626),
            .I(N__70572));
    Span4Mux_v I__15810 (
            .O(N__70617),
            .I(N__70572));
    InMux I__15809 (
            .O(N__70616),
            .I(N__70569));
    InMux I__15808 (
            .O(N__70615),
            .I(N__70566));
    InMux I__15807 (
            .O(N__70614),
            .I(N__70563));
    LocalMux I__15806 (
            .O(N__70611),
            .I(N__70556));
    Span4Mux_h I__15805 (
            .O(N__70608),
            .I(N__70556));
    LocalMux I__15804 (
            .O(N__70605),
            .I(N__70556));
    Span4Mux_h I__15803 (
            .O(N__70600),
            .I(N__70551));
    LocalMux I__15802 (
            .O(N__70595),
            .I(N__70551));
    LocalMux I__15801 (
            .O(N__70586),
            .I(xy_ki_2));
    LocalMux I__15800 (
            .O(N__70583),
            .I(xy_ki_2));
    LocalMux I__15799 (
            .O(N__70580),
            .I(xy_ki_2));
    Odrv4 I__15798 (
            .O(N__70577),
            .I(xy_ki_2));
    Odrv4 I__15797 (
            .O(N__70572),
            .I(xy_ki_2));
    LocalMux I__15796 (
            .O(N__70569),
            .I(xy_ki_2));
    LocalMux I__15795 (
            .O(N__70566),
            .I(xy_ki_2));
    LocalMux I__15794 (
            .O(N__70563),
            .I(xy_ki_2));
    Odrv4 I__15793 (
            .O(N__70556),
            .I(xy_ki_2));
    Odrv4 I__15792 (
            .O(N__70551),
            .I(xy_ki_2));
    CascadeMux I__15791 (
            .O(N__70530),
            .I(N__70522));
    CascadeMux I__15790 (
            .O(N__70529),
            .I(N__70518));
    InMux I__15789 (
            .O(N__70528),
            .I(N__70506));
    InMux I__15788 (
            .O(N__70527),
            .I(N__70503));
    InMux I__15787 (
            .O(N__70526),
            .I(N__70486));
    InMux I__15786 (
            .O(N__70525),
            .I(N__70486));
    InMux I__15785 (
            .O(N__70522),
            .I(N__70481));
    InMux I__15784 (
            .O(N__70521),
            .I(N__70481));
    InMux I__15783 (
            .O(N__70518),
            .I(N__70478));
    InMux I__15782 (
            .O(N__70517),
            .I(N__70475));
    CascadeMux I__15781 (
            .O(N__70516),
            .I(N__70472));
    CascadeMux I__15780 (
            .O(N__70515),
            .I(N__70463));
    CascadeMux I__15779 (
            .O(N__70514),
            .I(N__70460));
    InMux I__15778 (
            .O(N__70513),
            .I(N__70454));
    InMux I__15777 (
            .O(N__70512),
            .I(N__70446));
    InMux I__15776 (
            .O(N__70511),
            .I(N__70446));
    InMux I__15775 (
            .O(N__70510),
            .I(N__70446));
    InMux I__15774 (
            .O(N__70509),
            .I(N__70443));
    LocalMux I__15773 (
            .O(N__70506),
            .I(N__70438));
    LocalMux I__15772 (
            .O(N__70503),
            .I(N__70438));
    InMux I__15771 (
            .O(N__70502),
            .I(N__70435));
    CascadeMux I__15770 (
            .O(N__70501),
            .I(N__70428));
    InMux I__15769 (
            .O(N__70500),
            .I(N__70422));
    InMux I__15768 (
            .O(N__70499),
            .I(N__70422));
    InMux I__15767 (
            .O(N__70498),
            .I(N__70417));
    InMux I__15766 (
            .O(N__70497),
            .I(N__70417));
    CascadeMux I__15765 (
            .O(N__70496),
            .I(N__70412));
    CascadeMux I__15764 (
            .O(N__70495),
            .I(N__70404));
    CascadeMux I__15763 (
            .O(N__70494),
            .I(N__70400));
    InMux I__15762 (
            .O(N__70493),
            .I(N__70393));
    InMux I__15761 (
            .O(N__70492),
            .I(N__70393));
    InMux I__15760 (
            .O(N__70491),
            .I(N__70393));
    LocalMux I__15759 (
            .O(N__70486),
            .I(N__70384));
    LocalMux I__15758 (
            .O(N__70481),
            .I(N__70384));
    LocalMux I__15757 (
            .O(N__70478),
            .I(N__70384));
    LocalMux I__15756 (
            .O(N__70475),
            .I(N__70384));
    InMux I__15755 (
            .O(N__70472),
            .I(N__70381));
    InMux I__15754 (
            .O(N__70471),
            .I(N__70376));
    InMux I__15753 (
            .O(N__70470),
            .I(N__70371));
    InMux I__15752 (
            .O(N__70469),
            .I(N__70371));
    InMux I__15751 (
            .O(N__70468),
            .I(N__70366));
    InMux I__15750 (
            .O(N__70467),
            .I(N__70366));
    InMux I__15749 (
            .O(N__70466),
            .I(N__70361));
    InMux I__15748 (
            .O(N__70463),
            .I(N__70361));
    InMux I__15747 (
            .O(N__70460),
            .I(N__70355));
    InMux I__15746 (
            .O(N__70459),
            .I(N__70352));
    InMux I__15745 (
            .O(N__70458),
            .I(N__70347));
    InMux I__15744 (
            .O(N__70457),
            .I(N__70347));
    LocalMux I__15743 (
            .O(N__70454),
            .I(N__70344));
    InMux I__15742 (
            .O(N__70453),
            .I(N__70341));
    LocalMux I__15741 (
            .O(N__70446),
            .I(N__70332));
    LocalMux I__15740 (
            .O(N__70443),
            .I(N__70332));
    Span4Mux_v I__15739 (
            .O(N__70438),
            .I(N__70332));
    LocalMux I__15738 (
            .O(N__70435),
            .I(N__70332));
    InMux I__15737 (
            .O(N__70434),
            .I(N__70327));
    InMux I__15736 (
            .O(N__70433),
            .I(N__70327));
    InMux I__15735 (
            .O(N__70432),
            .I(N__70318));
    InMux I__15734 (
            .O(N__70431),
            .I(N__70318));
    InMux I__15733 (
            .O(N__70428),
            .I(N__70318));
    InMux I__15732 (
            .O(N__70427),
            .I(N__70318));
    LocalMux I__15731 (
            .O(N__70422),
            .I(N__70313));
    LocalMux I__15730 (
            .O(N__70417),
            .I(N__70313));
    CascadeMux I__15729 (
            .O(N__70416),
            .I(N__70309));
    CascadeMux I__15728 (
            .O(N__70415),
            .I(N__70305));
    InMux I__15727 (
            .O(N__70412),
            .I(N__70300));
    InMux I__15726 (
            .O(N__70411),
            .I(N__70300));
    CascadeMux I__15725 (
            .O(N__70410),
            .I(N__70297));
    InMux I__15724 (
            .O(N__70409),
            .I(N__70292));
    InMux I__15723 (
            .O(N__70408),
            .I(N__70283));
    InMux I__15722 (
            .O(N__70407),
            .I(N__70283));
    InMux I__15721 (
            .O(N__70404),
            .I(N__70283));
    InMux I__15720 (
            .O(N__70403),
            .I(N__70283));
    InMux I__15719 (
            .O(N__70400),
            .I(N__70280));
    LocalMux I__15718 (
            .O(N__70393),
            .I(N__70273));
    Span4Mux_v I__15717 (
            .O(N__70384),
            .I(N__70273));
    LocalMux I__15716 (
            .O(N__70381),
            .I(N__70273));
    InMux I__15715 (
            .O(N__70380),
            .I(N__70268));
    InMux I__15714 (
            .O(N__70379),
            .I(N__70268));
    LocalMux I__15713 (
            .O(N__70376),
            .I(N__70265));
    LocalMux I__15712 (
            .O(N__70371),
            .I(N__70260));
    LocalMux I__15711 (
            .O(N__70366),
            .I(N__70260));
    LocalMux I__15710 (
            .O(N__70361),
            .I(N__70257));
    InMux I__15709 (
            .O(N__70360),
            .I(N__70254));
    InMux I__15708 (
            .O(N__70359),
            .I(N__70247));
    InMux I__15707 (
            .O(N__70358),
            .I(N__70241));
    LocalMux I__15706 (
            .O(N__70355),
            .I(N__70236));
    LocalMux I__15705 (
            .O(N__70352),
            .I(N__70236));
    LocalMux I__15704 (
            .O(N__70347),
            .I(N__70233));
    Span4Mux_v I__15703 (
            .O(N__70344),
            .I(N__70228));
    LocalMux I__15702 (
            .O(N__70341),
            .I(N__70228));
    Span4Mux_h I__15701 (
            .O(N__70332),
            .I(N__70219));
    LocalMux I__15700 (
            .O(N__70327),
            .I(N__70219));
    LocalMux I__15699 (
            .O(N__70318),
            .I(N__70219));
    Span4Mux_v I__15698 (
            .O(N__70313),
            .I(N__70219));
    InMux I__15697 (
            .O(N__70312),
            .I(N__70216));
    InMux I__15696 (
            .O(N__70309),
            .I(N__70209));
    InMux I__15695 (
            .O(N__70308),
            .I(N__70209));
    InMux I__15694 (
            .O(N__70305),
            .I(N__70209));
    LocalMux I__15693 (
            .O(N__70300),
            .I(N__70206));
    InMux I__15692 (
            .O(N__70297),
            .I(N__70199));
    InMux I__15691 (
            .O(N__70296),
            .I(N__70199));
    InMux I__15690 (
            .O(N__70295),
            .I(N__70199));
    LocalMux I__15689 (
            .O(N__70292),
            .I(N__70188));
    LocalMux I__15688 (
            .O(N__70283),
            .I(N__70188));
    LocalMux I__15687 (
            .O(N__70280),
            .I(N__70188));
    Span4Mux_h I__15686 (
            .O(N__70273),
            .I(N__70188));
    LocalMux I__15685 (
            .O(N__70268),
            .I(N__70188));
    Span4Mux_v I__15684 (
            .O(N__70265),
            .I(N__70179));
    Span4Mux_v I__15683 (
            .O(N__70260),
            .I(N__70179));
    Span4Mux_h I__15682 (
            .O(N__70257),
            .I(N__70179));
    LocalMux I__15681 (
            .O(N__70254),
            .I(N__70179));
    InMux I__15680 (
            .O(N__70253),
            .I(N__70174));
    InMux I__15679 (
            .O(N__70252),
            .I(N__70174));
    InMux I__15678 (
            .O(N__70251),
            .I(N__70169));
    InMux I__15677 (
            .O(N__70250),
            .I(N__70169));
    LocalMux I__15676 (
            .O(N__70247),
            .I(N__70166));
    InMux I__15675 (
            .O(N__70246),
            .I(N__70161));
    InMux I__15674 (
            .O(N__70245),
            .I(N__70161));
    InMux I__15673 (
            .O(N__70244),
            .I(N__70158));
    LocalMux I__15672 (
            .O(N__70241),
            .I(N__70147));
    Span4Mux_h I__15671 (
            .O(N__70236),
            .I(N__70147));
    Span4Mux_v I__15670 (
            .O(N__70233),
            .I(N__70147));
    Span4Mux_h I__15669 (
            .O(N__70228),
            .I(N__70147));
    Span4Mux_v I__15668 (
            .O(N__70219),
            .I(N__70147));
    LocalMux I__15667 (
            .O(N__70216),
            .I(N__70142));
    LocalMux I__15666 (
            .O(N__70209),
            .I(N__70142));
    Span4Mux_h I__15665 (
            .O(N__70206),
            .I(N__70137));
    LocalMux I__15664 (
            .O(N__70199),
            .I(N__70137));
    Span4Mux_h I__15663 (
            .O(N__70188),
            .I(N__70130));
    Span4Mux_h I__15662 (
            .O(N__70179),
            .I(N__70130));
    LocalMux I__15661 (
            .O(N__70174),
            .I(N__70130));
    LocalMux I__15660 (
            .O(N__70169),
            .I(N__70125));
    Span12Mux_v I__15659 (
            .O(N__70166),
            .I(N__70125));
    LocalMux I__15658 (
            .O(N__70161),
            .I(xy_ki_3));
    LocalMux I__15657 (
            .O(N__70158),
            .I(xy_ki_3));
    Odrv4 I__15656 (
            .O(N__70147),
            .I(xy_ki_3));
    Odrv12 I__15655 (
            .O(N__70142),
            .I(xy_ki_3));
    Odrv4 I__15654 (
            .O(N__70137),
            .I(xy_ki_3));
    Odrv4 I__15653 (
            .O(N__70130),
            .I(xy_ki_3));
    Odrv12 I__15652 (
            .O(N__70125),
            .I(xy_ki_3));
    CascadeMux I__15651 (
            .O(N__70110),
            .I(\pid_side.N_37_1_cascade_ ));
    InMux I__15650 (
            .O(N__70107),
            .I(N__70104));
    LocalMux I__15649 (
            .O(N__70104),
            .I(N__70101));
    Span4Mux_s0_h I__15648 (
            .O(N__70101),
            .I(N__70096));
    InMux I__15647 (
            .O(N__70100),
            .I(N__70093));
    InMux I__15646 (
            .O(N__70099),
            .I(N__70084));
    Span4Mux_v I__15645 (
            .O(N__70096),
            .I(N__70074));
    LocalMux I__15644 (
            .O(N__70093),
            .I(N__70074));
    InMux I__15643 (
            .O(N__70092),
            .I(N__70069));
    InMux I__15642 (
            .O(N__70091),
            .I(N__70069));
    InMux I__15641 (
            .O(N__70090),
            .I(N__70060));
    InMux I__15640 (
            .O(N__70089),
            .I(N__70060));
    InMux I__15639 (
            .O(N__70088),
            .I(N__70060));
    InMux I__15638 (
            .O(N__70087),
            .I(N__70060));
    LocalMux I__15637 (
            .O(N__70084),
            .I(N__70057));
    InMux I__15636 (
            .O(N__70083),
            .I(N__70054));
    InMux I__15635 (
            .O(N__70082),
            .I(N__70051));
    InMux I__15634 (
            .O(N__70081),
            .I(N__70046));
    InMux I__15633 (
            .O(N__70080),
            .I(N__70046));
    InMux I__15632 (
            .O(N__70079),
            .I(N__70043));
    Span4Mux_v I__15631 (
            .O(N__70074),
            .I(N__70035));
    LocalMux I__15630 (
            .O(N__70069),
            .I(N__70030));
    LocalMux I__15629 (
            .O(N__70060),
            .I(N__70030));
    Span4Mux_v I__15628 (
            .O(N__70057),
            .I(N__70019));
    LocalMux I__15627 (
            .O(N__70054),
            .I(N__70019));
    LocalMux I__15626 (
            .O(N__70051),
            .I(N__70019));
    LocalMux I__15625 (
            .O(N__70046),
            .I(N__70019));
    LocalMux I__15624 (
            .O(N__70043),
            .I(N__70019));
    InMux I__15623 (
            .O(N__70042),
            .I(N__70014));
    InMux I__15622 (
            .O(N__70041),
            .I(N__70014));
    InMux I__15621 (
            .O(N__70040),
            .I(N__70009));
    InMux I__15620 (
            .O(N__70039),
            .I(N__70004));
    InMux I__15619 (
            .O(N__70038),
            .I(N__70004));
    Span4Mux_h I__15618 (
            .O(N__70035),
            .I(N__69999));
    Span4Mux_v I__15617 (
            .O(N__70030),
            .I(N__69999));
    Span4Mux_v I__15616 (
            .O(N__70019),
            .I(N__69994));
    LocalMux I__15615 (
            .O(N__70014),
            .I(N__69994));
    InMux I__15614 (
            .O(N__70013),
            .I(N__69989));
    InMux I__15613 (
            .O(N__70012),
            .I(N__69989));
    LocalMux I__15612 (
            .O(N__70009),
            .I(\pid_side.error_15 ));
    LocalMux I__15611 (
            .O(N__70004),
            .I(\pid_side.error_15 ));
    Odrv4 I__15610 (
            .O(N__69999),
            .I(\pid_side.error_15 ));
    Odrv4 I__15609 (
            .O(N__69994),
            .I(\pid_side.error_15 ));
    LocalMux I__15608 (
            .O(N__69989),
            .I(\pid_side.error_15 ));
    CascadeMux I__15607 (
            .O(N__69978),
            .I(N__69974));
    CascadeMux I__15606 (
            .O(N__69977),
            .I(N__69971));
    InMux I__15605 (
            .O(N__69974),
            .I(N__69966));
    InMux I__15604 (
            .O(N__69971),
            .I(N__69961));
    InMux I__15603 (
            .O(N__69970),
            .I(N__69961));
    CascadeMux I__15602 (
            .O(N__69969),
            .I(N__69958));
    LocalMux I__15601 (
            .O(N__69966),
            .I(N__69946));
    LocalMux I__15600 (
            .O(N__69961),
            .I(N__69943));
    InMux I__15599 (
            .O(N__69958),
            .I(N__69940));
    InMux I__15598 (
            .O(N__69957),
            .I(N__69937));
    InMux I__15597 (
            .O(N__69956),
            .I(N__69934));
    CascadeMux I__15596 (
            .O(N__69955),
            .I(N__69930));
    CascadeMux I__15595 (
            .O(N__69954),
            .I(N__69925));
    InMux I__15594 (
            .O(N__69953),
            .I(N__69922));
    InMux I__15593 (
            .O(N__69952),
            .I(N__69919));
    CascadeMux I__15592 (
            .O(N__69951),
            .I(N__69916));
    InMux I__15591 (
            .O(N__69950),
            .I(N__69909));
    InMux I__15590 (
            .O(N__69949),
            .I(N__69909));
    Span4Mux_h I__15589 (
            .O(N__69946),
            .I(N__69898));
    Span4Mux_h I__15588 (
            .O(N__69943),
            .I(N__69898));
    LocalMux I__15587 (
            .O(N__69940),
            .I(N__69898));
    LocalMux I__15586 (
            .O(N__69937),
            .I(N__69898));
    LocalMux I__15585 (
            .O(N__69934),
            .I(N__69898));
    InMux I__15584 (
            .O(N__69933),
            .I(N__69893));
    InMux I__15583 (
            .O(N__69930),
            .I(N__69893));
    InMux I__15582 (
            .O(N__69929),
            .I(N__69890));
    InMux I__15581 (
            .O(N__69928),
            .I(N__69887));
    InMux I__15580 (
            .O(N__69925),
            .I(N__69883));
    LocalMux I__15579 (
            .O(N__69922),
            .I(N__69880));
    LocalMux I__15578 (
            .O(N__69919),
            .I(N__69877));
    InMux I__15577 (
            .O(N__69916),
            .I(N__69874));
    InMux I__15576 (
            .O(N__69915),
            .I(N__69869));
    CascadeMux I__15575 (
            .O(N__69914),
            .I(N__69862));
    LocalMux I__15574 (
            .O(N__69909),
            .I(N__69854));
    Span4Mux_v I__15573 (
            .O(N__69898),
            .I(N__69854));
    LocalMux I__15572 (
            .O(N__69893),
            .I(N__69854));
    LocalMux I__15571 (
            .O(N__69890),
            .I(N__69848));
    LocalMux I__15570 (
            .O(N__69887),
            .I(N__69844));
    InMux I__15569 (
            .O(N__69886),
            .I(N__69841));
    LocalMux I__15568 (
            .O(N__69883),
            .I(N__69832));
    Span4Mux_h I__15567 (
            .O(N__69880),
            .I(N__69832));
    Span4Mux_h I__15566 (
            .O(N__69877),
            .I(N__69832));
    LocalMux I__15565 (
            .O(N__69874),
            .I(N__69832));
    InMux I__15564 (
            .O(N__69873),
            .I(N__69829));
    InMux I__15563 (
            .O(N__69872),
            .I(N__69826));
    LocalMux I__15562 (
            .O(N__69869),
            .I(N__69823));
    InMux I__15561 (
            .O(N__69868),
            .I(N__69820));
    CascadeMux I__15560 (
            .O(N__69867),
            .I(N__69817));
    InMux I__15559 (
            .O(N__69866),
            .I(N__69813));
    InMux I__15558 (
            .O(N__69865),
            .I(N__69810));
    InMux I__15557 (
            .O(N__69862),
            .I(N__69805));
    InMux I__15556 (
            .O(N__69861),
            .I(N__69805));
    Span4Mux_h I__15555 (
            .O(N__69854),
            .I(N__69802));
    InMux I__15554 (
            .O(N__69853),
            .I(N__69799));
    InMux I__15553 (
            .O(N__69852),
            .I(N__69796));
    InMux I__15552 (
            .O(N__69851),
            .I(N__69793));
    Span4Mux_v I__15551 (
            .O(N__69848),
            .I(N__69790));
    InMux I__15550 (
            .O(N__69847),
            .I(N__69787));
    Span4Mux_h I__15549 (
            .O(N__69844),
            .I(N__69781));
    LocalMux I__15548 (
            .O(N__69841),
            .I(N__69781));
    Span4Mux_v I__15547 (
            .O(N__69832),
            .I(N__69778));
    LocalMux I__15546 (
            .O(N__69829),
            .I(N__69775));
    LocalMux I__15545 (
            .O(N__69826),
            .I(N__69770));
    Span4Mux_h I__15544 (
            .O(N__69823),
            .I(N__69770));
    LocalMux I__15543 (
            .O(N__69820),
            .I(N__69767));
    InMux I__15542 (
            .O(N__69817),
            .I(N__69762));
    InMux I__15541 (
            .O(N__69816),
            .I(N__69759));
    LocalMux I__15540 (
            .O(N__69813),
            .I(N__69748));
    LocalMux I__15539 (
            .O(N__69810),
            .I(N__69748));
    LocalMux I__15538 (
            .O(N__69805),
            .I(N__69748));
    Span4Mux_h I__15537 (
            .O(N__69802),
            .I(N__69748));
    LocalMux I__15536 (
            .O(N__69799),
            .I(N__69748));
    LocalMux I__15535 (
            .O(N__69796),
            .I(N__69745));
    LocalMux I__15534 (
            .O(N__69793),
            .I(N__69740));
    Span4Mux_h I__15533 (
            .O(N__69790),
            .I(N__69740));
    LocalMux I__15532 (
            .O(N__69787),
            .I(N__69737));
    InMux I__15531 (
            .O(N__69786),
            .I(N__69734));
    Span4Mux_v I__15530 (
            .O(N__69781),
            .I(N__69723));
    Span4Mux_h I__15529 (
            .O(N__69778),
            .I(N__69723));
    Span4Mux_h I__15528 (
            .O(N__69775),
            .I(N__69723));
    Span4Mux_v I__15527 (
            .O(N__69770),
            .I(N__69723));
    Span4Mux_v I__15526 (
            .O(N__69767),
            .I(N__69723));
    InMux I__15525 (
            .O(N__69766),
            .I(N__69718));
    InMux I__15524 (
            .O(N__69765),
            .I(N__69718));
    LocalMux I__15523 (
            .O(N__69762),
            .I(N__69711));
    LocalMux I__15522 (
            .O(N__69759),
            .I(N__69711));
    Span4Mux_v I__15521 (
            .O(N__69748),
            .I(N__69711));
    Odrv4 I__15520 (
            .O(N__69745),
            .I(pid_front_N_331));
    Odrv4 I__15519 (
            .O(N__69740),
            .I(pid_front_N_331));
    Odrv12 I__15518 (
            .O(N__69737),
            .I(pid_front_N_331));
    LocalMux I__15517 (
            .O(N__69734),
            .I(pid_front_N_331));
    Odrv4 I__15516 (
            .O(N__69723),
            .I(pid_front_N_331));
    LocalMux I__15515 (
            .O(N__69718),
            .I(pid_front_N_331));
    Odrv4 I__15514 (
            .O(N__69711),
            .I(pid_front_N_331));
    InMux I__15513 (
            .O(N__69696),
            .I(N__69692));
    InMux I__15512 (
            .O(N__69695),
            .I(N__69689));
    LocalMux I__15511 (
            .O(N__69692),
            .I(N__69683));
    LocalMux I__15510 (
            .O(N__69689),
            .I(N__69683));
    InMux I__15509 (
            .O(N__69688),
            .I(N__69676));
    Span4Mux_v I__15508 (
            .O(N__69683),
            .I(N__69673));
    InMux I__15507 (
            .O(N__69682),
            .I(N__69668));
    InMux I__15506 (
            .O(N__69681),
            .I(N__69668));
    CascadeMux I__15505 (
            .O(N__69680),
            .I(N__69663));
    InMux I__15504 (
            .O(N__69679),
            .I(N__69648));
    LocalMux I__15503 (
            .O(N__69676),
            .I(N__69645));
    Span4Mux_h I__15502 (
            .O(N__69673),
            .I(N__69640));
    LocalMux I__15501 (
            .O(N__69668),
            .I(N__69640));
    InMux I__15500 (
            .O(N__69667),
            .I(N__69637));
    InMux I__15499 (
            .O(N__69666),
            .I(N__69627));
    InMux I__15498 (
            .O(N__69663),
            .I(N__69627));
    InMux I__15497 (
            .O(N__69662),
            .I(N__69620));
    InMux I__15496 (
            .O(N__69661),
            .I(N__69620));
    InMux I__15495 (
            .O(N__69660),
            .I(N__69617));
    InMux I__15494 (
            .O(N__69659),
            .I(N__69614));
    InMux I__15493 (
            .O(N__69658),
            .I(N__69611));
    InMux I__15492 (
            .O(N__69657),
            .I(N__69608));
    InMux I__15491 (
            .O(N__69656),
            .I(N__69603));
    InMux I__15490 (
            .O(N__69655),
            .I(N__69603));
    InMux I__15489 (
            .O(N__69654),
            .I(N__69596));
    InMux I__15488 (
            .O(N__69653),
            .I(N__69591));
    InMux I__15487 (
            .O(N__69652),
            .I(N__69591));
    InMux I__15486 (
            .O(N__69651),
            .I(N__69588));
    LocalMux I__15485 (
            .O(N__69648),
            .I(N__69577));
    Span4Mux_h I__15484 (
            .O(N__69645),
            .I(N__69577));
    Span4Mux_h I__15483 (
            .O(N__69640),
            .I(N__69577));
    LocalMux I__15482 (
            .O(N__69637),
            .I(N__69577));
    InMux I__15481 (
            .O(N__69636),
            .I(N__69573));
    InMux I__15480 (
            .O(N__69635),
            .I(N__69570));
    InMux I__15479 (
            .O(N__69634),
            .I(N__69567));
    InMux I__15478 (
            .O(N__69633),
            .I(N__69560));
    InMux I__15477 (
            .O(N__69632),
            .I(N__69560));
    LocalMux I__15476 (
            .O(N__69627),
            .I(N__69557));
    InMux I__15475 (
            .O(N__69626),
            .I(N__69554));
    InMux I__15474 (
            .O(N__69625),
            .I(N__69551));
    LocalMux I__15473 (
            .O(N__69620),
            .I(N__69545));
    LocalMux I__15472 (
            .O(N__69617),
            .I(N__69545));
    LocalMux I__15471 (
            .O(N__69614),
            .I(N__69538));
    LocalMux I__15470 (
            .O(N__69611),
            .I(N__69538));
    LocalMux I__15469 (
            .O(N__69608),
            .I(N__69538));
    LocalMux I__15468 (
            .O(N__69603),
            .I(N__69531));
    CascadeMux I__15467 (
            .O(N__69602),
            .I(N__69528));
    InMux I__15466 (
            .O(N__69601),
            .I(N__69523));
    InMux I__15465 (
            .O(N__69600),
            .I(N__69523));
    InMux I__15464 (
            .O(N__69599),
            .I(N__69520));
    LocalMux I__15463 (
            .O(N__69596),
            .I(N__69513));
    LocalMux I__15462 (
            .O(N__69591),
            .I(N__69513));
    LocalMux I__15461 (
            .O(N__69588),
            .I(N__69513));
    InMux I__15460 (
            .O(N__69587),
            .I(N__69508));
    InMux I__15459 (
            .O(N__69586),
            .I(N__69508));
    Span4Mux_v I__15458 (
            .O(N__69577),
            .I(N__69505));
    InMux I__15457 (
            .O(N__69576),
            .I(N__69502));
    LocalMux I__15456 (
            .O(N__69573),
            .I(N__69497));
    LocalMux I__15455 (
            .O(N__69570),
            .I(N__69494));
    LocalMux I__15454 (
            .O(N__69567),
            .I(N__69491));
    InMux I__15453 (
            .O(N__69566),
            .I(N__69486));
    InMux I__15452 (
            .O(N__69565),
            .I(N__69486));
    LocalMux I__15451 (
            .O(N__69560),
            .I(N__69481));
    Span4Mux_h I__15450 (
            .O(N__69557),
            .I(N__69481));
    LocalMux I__15449 (
            .O(N__69554),
            .I(N__69477));
    LocalMux I__15448 (
            .O(N__69551),
            .I(N__69474));
    InMux I__15447 (
            .O(N__69550),
            .I(N__69471));
    Span4Mux_v I__15446 (
            .O(N__69545),
            .I(N__69466));
    Span4Mux_v I__15445 (
            .O(N__69538),
            .I(N__69466));
    InMux I__15444 (
            .O(N__69537),
            .I(N__69459));
    InMux I__15443 (
            .O(N__69536),
            .I(N__69459));
    InMux I__15442 (
            .O(N__69535),
            .I(N__69459));
    CascadeMux I__15441 (
            .O(N__69534),
            .I(N__69456));
    Span4Mux_h I__15440 (
            .O(N__69531),
            .I(N__69453));
    InMux I__15439 (
            .O(N__69528),
            .I(N__69450));
    LocalMux I__15438 (
            .O(N__69523),
            .I(N__69447));
    LocalMux I__15437 (
            .O(N__69520),
            .I(N__69444));
    Span4Mux_v I__15436 (
            .O(N__69513),
            .I(N__69435));
    LocalMux I__15435 (
            .O(N__69508),
            .I(N__69435));
    Span4Mux_h I__15434 (
            .O(N__69505),
            .I(N__69435));
    LocalMux I__15433 (
            .O(N__69502),
            .I(N__69435));
    InMux I__15432 (
            .O(N__69501),
            .I(N__69430));
    InMux I__15431 (
            .O(N__69500),
            .I(N__69430));
    Span4Mux_h I__15430 (
            .O(N__69497),
            .I(N__69425));
    Span4Mux_v I__15429 (
            .O(N__69494),
            .I(N__69425));
    Span4Mux_v I__15428 (
            .O(N__69491),
            .I(N__69418));
    LocalMux I__15427 (
            .O(N__69486),
            .I(N__69418));
    Span4Mux_h I__15426 (
            .O(N__69481),
            .I(N__69418));
    InMux I__15425 (
            .O(N__69480),
            .I(N__69415));
    Span4Mux_h I__15424 (
            .O(N__69477),
            .I(N__69410));
    Span4Mux_v I__15423 (
            .O(N__69474),
            .I(N__69410));
    LocalMux I__15422 (
            .O(N__69471),
            .I(N__69403));
    Span4Mux_h I__15421 (
            .O(N__69466),
            .I(N__69403));
    LocalMux I__15420 (
            .O(N__69459),
            .I(N__69403));
    InMux I__15419 (
            .O(N__69456),
            .I(N__69400));
    Span4Mux_v I__15418 (
            .O(N__69453),
            .I(N__69395));
    LocalMux I__15417 (
            .O(N__69450),
            .I(N__69395));
    Span4Mux_v I__15416 (
            .O(N__69447),
            .I(N__69388));
    Span4Mux_v I__15415 (
            .O(N__69444),
            .I(N__69388));
    Span4Mux_v I__15414 (
            .O(N__69435),
            .I(N__69388));
    LocalMux I__15413 (
            .O(N__69430),
            .I(N__69379));
    Sp12to4 I__15412 (
            .O(N__69425),
            .I(N__69379));
    Sp12to4 I__15411 (
            .O(N__69418),
            .I(N__69379));
    LocalMux I__15410 (
            .O(N__69415),
            .I(N__69379));
    Span4Mux_v I__15409 (
            .O(N__69410),
            .I(N__69374));
    Span4Mux_v I__15408 (
            .O(N__69403),
            .I(N__69374));
    LocalMux I__15407 (
            .O(N__69400),
            .I(N__69367));
    Span4Mux_v I__15406 (
            .O(N__69395),
            .I(N__69367));
    Span4Mux_v I__15405 (
            .O(N__69388),
            .I(N__69367));
    Span12Mux_s11_v I__15404 (
            .O(N__69379),
            .I(N__69364));
    Odrv4 I__15403 (
            .O(N__69374),
            .I(xy_ki_4));
    Odrv4 I__15402 (
            .O(N__69367),
            .I(xy_ki_4));
    Odrv12 I__15401 (
            .O(N__69364),
            .I(xy_ki_4));
    CascadeMux I__15400 (
            .O(N__69357),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ));
    InMux I__15399 (
            .O(N__69354),
            .I(N__69351));
    LocalMux I__15398 (
            .O(N__69351),
            .I(N__69348));
    Span4Mux_h I__15397 (
            .O(N__69348),
            .I(N__69345));
    Odrv4 I__15396 (
            .O(N__69345),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_22 ));
    CascadeMux I__15395 (
            .O(N__69342),
            .I(N__69339));
    InMux I__15394 (
            .O(N__69339),
            .I(N__69336));
    LocalMux I__15393 (
            .O(N__69336),
            .I(N__69333));
    Span4Mux_h I__15392 (
            .O(N__69333),
            .I(N__69330));
    Span4Mux_v I__15391 (
            .O(N__69330),
            .I(N__69327));
    Odrv4 I__15390 (
            .O(N__69327),
            .I(\pid_side.error_i_regZ0Z_22 ));
    CEMux I__15389 (
            .O(N__69324),
            .I(N__69318));
    CEMux I__15388 (
            .O(N__69323),
            .I(N__69313));
    CEMux I__15387 (
            .O(N__69322),
            .I(N__69310));
    CEMux I__15386 (
            .O(N__69321),
            .I(N__69307));
    LocalMux I__15385 (
            .O(N__69318),
            .I(N__69300));
    CEMux I__15384 (
            .O(N__69317),
            .I(N__69296));
    CEMux I__15383 (
            .O(N__69316),
            .I(N__69293));
    LocalMux I__15382 (
            .O(N__69313),
            .I(N__69290));
    LocalMux I__15381 (
            .O(N__69310),
            .I(N__69287));
    LocalMux I__15380 (
            .O(N__69307),
            .I(N__69284));
    CEMux I__15379 (
            .O(N__69306),
            .I(N__69281));
    CEMux I__15378 (
            .O(N__69305),
            .I(N__69278));
    CEMux I__15377 (
            .O(N__69304),
            .I(N__69275));
    CEMux I__15376 (
            .O(N__69303),
            .I(N__69272));
    Span4Mux_h I__15375 (
            .O(N__69300),
            .I(N__69269));
    CEMux I__15374 (
            .O(N__69299),
            .I(N__69266));
    LocalMux I__15373 (
            .O(N__69296),
            .I(N__69261));
    LocalMux I__15372 (
            .O(N__69293),
            .I(N__69261));
    Span4Mux_h I__15371 (
            .O(N__69290),
            .I(N__69257));
    Span4Mux_v I__15370 (
            .O(N__69287),
            .I(N__69254));
    Span4Mux_h I__15369 (
            .O(N__69284),
            .I(N__69249));
    LocalMux I__15368 (
            .O(N__69281),
            .I(N__69249));
    LocalMux I__15367 (
            .O(N__69278),
            .I(N__69246));
    LocalMux I__15366 (
            .O(N__69275),
            .I(N__69243));
    LocalMux I__15365 (
            .O(N__69272),
            .I(N__69236));
    Span4Mux_h I__15364 (
            .O(N__69269),
            .I(N__69236));
    LocalMux I__15363 (
            .O(N__69266),
            .I(N__69236));
    Span4Mux_h I__15362 (
            .O(N__69261),
            .I(N__69233));
    CEMux I__15361 (
            .O(N__69260),
            .I(N__69230));
    Span4Mux_h I__15360 (
            .O(N__69257),
            .I(N__69225));
    Span4Mux_h I__15359 (
            .O(N__69254),
            .I(N__69225));
    Span4Mux_h I__15358 (
            .O(N__69249),
            .I(N__69222));
    Span4Mux_h I__15357 (
            .O(N__69246),
            .I(N__69219));
    Span4Mux_h I__15356 (
            .O(N__69243),
            .I(N__69216));
    Span4Mux_v I__15355 (
            .O(N__69236),
            .I(N__69213));
    Span4Mux_h I__15354 (
            .O(N__69233),
            .I(N__69210));
    LocalMux I__15353 (
            .O(N__69230),
            .I(N__69207));
    Span4Mux_v I__15352 (
            .O(N__69225),
            .I(N__69202));
    Span4Mux_v I__15351 (
            .O(N__69222),
            .I(N__69202));
    Span4Mux_h I__15350 (
            .O(N__69219),
            .I(N__69199));
    Span4Mux_v I__15349 (
            .O(N__69216),
            .I(N__69194));
    Span4Mux_h I__15348 (
            .O(N__69213),
            .I(N__69194));
    Span4Mux_v I__15347 (
            .O(N__69210),
            .I(N__69191));
    Sp12to4 I__15346 (
            .O(N__69207),
            .I(N__69188));
    Span4Mux_v I__15345 (
            .O(N__69202),
            .I(N__69185));
    Span4Mux_v I__15344 (
            .O(N__69199),
            .I(N__69182));
    Span4Mux_h I__15343 (
            .O(N__69194),
            .I(N__69177));
    Span4Mux_v I__15342 (
            .O(N__69191),
            .I(N__69177));
    Span12Mux_v I__15341 (
            .O(N__69188),
            .I(N__69172));
    Sp12to4 I__15340 (
            .O(N__69185),
            .I(N__69172));
    Odrv4 I__15339 (
            .O(N__69182),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__15338 (
            .O(N__69177),
            .I(\pid_side.state_ns_0_0 ));
    Odrv12 I__15337 (
            .O(N__69172),
            .I(\pid_side.state_ns_0_0 ));
    InMux I__15336 (
            .O(N__69165),
            .I(N__69159));
    InMux I__15335 (
            .O(N__69164),
            .I(N__69153));
    InMux I__15334 (
            .O(N__69163),
            .I(N__69150));
    InMux I__15333 (
            .O(N__69162),
            .I(N__69147));
    LocalMux I__15332 (
            .O(N__69159),
            .I(N__69143));
    InMux I__15331 (
            .O(N__69158),
            .I(N__69137));
    InMux I__15330 (
            .O(N__69157),
            .I(N__69137));
    InMux I__15329 (
            .O(N__69156),
            .I(N__69134));
    LocalMux I__15328 (
            .O(N__69153),
            .I(N__69130));
    LocalMux I__15327 (
            .O(N__69150),
            .I(N__69125));
    LocalMux I__15326 (
            .O(N__69147),
            .I(N__69125));
    InMux I__15325 (
            .O(N__69146),
            .I(N__69122));
    Span4Mux_v I__15324 (
            .O(N__69143),
            .I(N__69119));
    InMux I__15323 (
            .O(N__69142),
            .I(N__69116));
    LocalMux I__15322 (
            .O(N__69137),
            .I(N__69111));
    LocalMux I__15321 (
            .O(N__69134),
            .I(N__69111));
    InMux I__15320 (
            .O(N__69133),
            .I(N__69108));
    Sp12to4 I__15319 (
            .O(N__69130),
            .I(N__69105));
    Span12Mux_v I__15318 (
            .O(N__69125),
            .I(N__69102));
    LocalMux I__15317 (
            .O(N__69122),
            .I(N__69099));
    Span4Mux_h I__15316 (
            .O(N__69119),
            .I(N__69094));
    LocalMux I__15315 (
            .O(N__69116),
            .I(N__69094));
    Span4Mux_h I__15314 (
            .O(N__69111),
            .I(N__69091));
    LocalMux I__15313 (
            .O(N__69108),
            .I(drone_H_disp_side_0));
    Odrv12 I__15312 (
            .O(N__69105),
            .I(drone_H_disp_side_0));
    Odrv12 I__15311 (
            .O(N__69102),
            .I(drone_H_disp_side_0));
    Odrv4 I__15310 (
            .O(N__69099),
            .I(drone_H_disp_side_0));
    Odrv4 I__15309 (
            .O(N__69094),
            .I(drone_H_disp_side_0));
    Odrv4 I__15308 (
            .O(N__69091),
            .I(drone_H_disp_side_0));
    CascadeMux I__15307 (
            .O(N__69078),
            .I(N__69075));
    InMux I__15306 (
            .O(N__69075),
            .I(N__69072));
    LocalMux I__15305 (
            .O(N__69072),
            .I(N__69069));
    Odrv12 I__15304 (
            .O(N__69069),
            .I(side_command_4));
    InMux I__15303 (
            .O(N__69066),
            .I(bfn_18_20_0_));
    InMux I__15302 (
            .O(N__69063),
            .I(N__69060));
    LocalMux I__15301 (
            .O(N__69060),
            .I(N__69057));
    Odrv4 I__15300 (
            .O(N__69057),
            .I(drone_H_disp_side_i_9));
    CascadeMux I__15299 (
            .O(N__69054),
            .I(N__69051));
    InMux I__15298 (
            .O(N__69051),
            .I(N__69048));
    LocalMux I__15297 (
            .O(N__69048),
            .I(N__69045));
    Odrv4 I__15296 (
            .O(N__69045),
            .I(side_command_5));
    InMux I__15295 (
            .O(N__69042),
            .I(N__69033));
    InMux I__15294 (
            .O(N__69041),
            .I(N__69029));
    InMux I__15293 (
            .O(N__69040),
            .I(N__69020));
    InMux I__15292 (
            .O(N__69039),
            .I(N__69020));
    InMux I__15291 (
            .O(N__69038),
            .I(N__69020));
    InMux I__15290 (
            .O(N__69037),
            .I(N__69020));
    CascadeMux I__15289 (
            .O(N__69036),
            .I(N__69017));
    LocalMux I__15288 (
            .O(N__69033),
            .I(N__69013));
    InMux I__15287 (
            .O(N__69032),
            .I(N__69010));
    LocalMux I__15286 (
            .O(N__69029),
            .I(N__69007));
    LocalMux I__15285 (
            .O(N__69020),
            .I(N__69004));
    InMux I__15284 (
            .O(N__69017),
            .I(N__68999));
    InMux I__15283 (
            .O(N__69016),
            .I(N__68999));
    Span12Mux_s7_h I__15282 (
            .O(N__69013),
            .I(N__68996));
    LocalMux I__15281 (
            .O(N__69010),
            .I(N__68991));
    Span12Mux_v I__15280 (
            .O(N__69007),
            .I(N__68991));
    Span4Mux_h I__15279 (
            .O(N__69004),
            .I(N__68988));
    LocalMux I__15278 (
            .O(N__68999),
            .I(\pid_side.error_9 ));
    Odrv12 I__15277 (
            .O(N__68996),
            .I(\pid_side.error_9 ));
    Odrv12 I__15276 (
            .O(N__68991),
            .I(\pid_side.error_9 ));
    Odrv4 I__15275 (
            .O(N__68988),
            .I(\pid_side.error_9 ));
    InMux I__15274 (
            .O(N__68979),
            .I(\pid_side.error_cry_4 ));
    CascadeMux I__15273 (
            .O(N__68976),
            .I(N__68973));
    InMux I__15272 (
            .O(N__68973),
            .I(N__68970));
    LocalMux I__15271 (
            .O(N__68970),
            .I(N__68967));
    Odrv4 I__15270 (
            .O(N__68967),
            .I(side_command_6));
    InMux I__15269 (
            .O(N__68964),
            .I(\pid_side.error_cry_5 ));
    InMux I__15268 (
            .O(N__68961),
            .I(N__68958));
    LocalMux I__15267 (
            .O(N__68958),
            .I(\pid_side.error_axbZ0Z_7 ));
    InMux I__15266 (
            .O(N__68955),
            .I(\pid_side.error_cry_6 ));
    InMux I__15265 (
            .O(N__68952),
            .I(N__68949));
    LocalMux I__15264 (
            .O(N__68949),
            .I(\pid_side.error_axb_8_l_ofxZ0 ));
    CascadeMux I__15263 (
            .O(N__68946),
            .I(N__68943));
    InMux I__15262 (
            .O(N__68943),
            .I(N__68937));
    InMux I__15261 (
            .O(N__68942),
            .I(N__68930));
    InMux I__15260 (
            .O(N__68941),
            .I(N__68930));
    InMux I__15259 (
            .O(N__68940),
            .I(N__68930));
    LocalMux I__15258 (
            .O(N__68937),
            .I(drone_H_disp_side_12));
    LocalMux I__15257 (
            .O(N__68930),
            .I(drone_H_disp_side_12));
    InMux I__15256 (
            .O(N__68925),
            .I(\pid_side.error_cry_7 ));
    InMux I__15255 (
            .O(N__68922),
            .I(N__68919));
    LocalMux I__15254 (
            .O(N__68919),
            .I(drone_H_disp_side_i_12));
    CascadeMux I__15253 (
            .O(N__68916),
            .I(N__68913));
    InMux I__15252 (
            .O(N__68913),
            .I(N__68910));
    LocalMux I__15251 (
            .O(N__68910),
            .I(N__68905));
    InMux I__15250 (
            .O(N__68909),
            .I(N__68900));
    InMux I__15249 (
            .O(N__68908),
            .I(N__68900));
    Odrv4 I__15248 (
            .O(N__68905),
            .I(drone_H_disp_side_13));
    LocalMux I__15247 (
            .O(N__68900),
            .I(drone_H_disp_side_13));
    InMux I__15246 (
            .O(N__68895),
            .I(\pid_side.error_cry_8 ));
    InMux I__15245 (
            .O(N__68892),
            .I(N__68889));
    LocalMux I__15244 (
            .O(N__68889),
            .I(N__68886));
    Odrv4 I__15243 (
            .O(N__68886),
            .I(drone_H_disp_side_i_13));
    InMux I__15242 (
            .O(N__68883),
            .I(\pid_side.error_cry_9 ));
    CascadeMux I__15241 (
            .O(N__68880),
            .I(N__68877));
    InMux I__15240 (
            .O(N__68877),
            .I(N__68873));
    InMux I__15239 (
            .O(N__68876),
            .I(N__68870));
    LocalMux I__15238 (
            .O(N__68873),
            .I(drone_H_disp_side_15));
    LocalMux I__15237 (
            .O(N__68870),
            .I(drone_H_disp_side_15));
    CascadeMux I__15236 (
            .O(N__68865),
            .I(N__68861));
    InMux I__15235 (
            .O(N__68864),
            .I(N__68855));
    InMux I__15234 (
            .O(N__68861),
            .I(N__68855));
    InMux I__15233 (
            .O(N__68860),
            .I(N__68852));
    LocalMux I__15232 (
            .O(N__68855),
            .I(N__68849));
    LocalMux I__15231 (
            .O(N__68852),
            .I(N__68844));
    Span4Mux_v I__15230 (
            .O(N__68849),
            .I(N__68844));
    Odrv4 I__15229 (
            .O(N__68844),
            .I(drone_H_disp_side_14));
    InMux I__15228 (
            .O(N__68841),
            .I(\pid_side.error_cry_10 ));
    CascadeMux I__15227 (
            .O(N__68838),
            .I(N__68835));
    InMux I__15226 (
            .O(N__68835),
            .I(N__68832));
    LocalMux I__15225 (
            .O(N__68832),
            .I(\pid_side.error_axb_0 ));
    CascadeMux I__15224 (
            .O(N__68829),
            .I(N__68826));
    InMux I__15223 (
            .O(N__68826),
            .I(N__68823));
    LocalMux I__15222 (
            .O(N__68823),
            .I(N__68820));
    Span4Mux_h I__15221 (
            .O(N__68820),
            .I(N__68817));
    Span4Mux_h I__15220 (
            .O(N__68817),
            .I(N__68814));
    Span4Mux_h I__15219 (
            .O(N__68814),
            .I(N__68811));
    Odrv4 I__15218 (
            .O(N__68811),
            .I(\pid_side.error_axbZ0Z_1 ));
    InMux I__15217 (
            .O(N__68808),
            .I(\pid_side.error_cry_0 ));
    InMux I__15216 (
            .O(N__68805),
            .I(N__68802));
    LocalMux I__15215 (
            .O(N__68802),
            .I(\pid_side.error_axbZ0Z_2 ));
    InMux I__15214 (
            .O(N__68799),
            .I(\pid_side.error_cry_1 ));
    InMux I__15213 (
            .O(N__68796),
            .I(N__68793));
    LocalMux I__15212 (
            .O(N__68793),
            .I(N__68790));
    Span4Mux_h I__15211 (
            .O(N__68790),
            .I(N__68787));
    Span4Mux_v I__15210 (
            .O(N__68787),
            .I(N__68784));
    Span4Mux_h I__15209 (
            .O(N__68784),
            .I(N__68781));
    Span4Mux_h I__15208 (
            .O(N__68781),
            .I(N__68778));
    Odrv4 I__15207 (
            .O(N__68778),
            .I(\pid_side.error_axbZ0Z_3 ));
    InMux I__15206 (
            .O(N__68775),
            .I(\pid_side.error_cry_2 ));
    InMux I__15205 (
            .O(N__68772),
            .I(N__68769));
    LocalMux I__15204 (
            .O(N__68769),
            .I(side_command_0));
    CascadeMux I__15203 (
            .O(N__68766),
            .I(N__68763));
    InMux I__15202 (
            .O(N__68763),
            .I(N__68760));
    LocalMux I__15201 (
            .O(N__68760),
            .I(N__68757));
    Odrv4 I__15200 (
            .O(N__68757),
            .I(drone_H_disp_side_i_4));
    InMux I__15199 (
            .O(N__68754),
            .I(\pid_side.error_cry_3 ));
    InMux I__15198 (
            .O(N__68751),
            .I(N__68748));
    LocalMux I__15197 (
            .O(N__68748),
            .I(side_command_1));
    CascadeMux I__15196 (
            .O(N__68745),
            .I(N__68742));
    InMux I__15195 (
            .O(N__68742),
            .I(N__68739));
    LocalMux I__15194 (
            .O(N__68739),
            .I(drone_H_disp_side_i_5));
    InMux I__15193 (
            .O(N__68736),
            .I(\pid_side.error_cry_0_0 ));
    InMux I__15192 (
            .O(N__68733),
            .I(N__68730));
    LocalMux I__15191 (
            .O(N__68730),
            .I(drone_H_disp_side_i_6));
    CascadeMux I__15190 (
            .O(N__68727),
            .I(N__68724));
    InMux I__15189 (
            .O(N__68724),
            .I(N__68721));
    LocalMux I__15188 (
            .O(N__68721),
            .I(side_command_2));
    InMux I__15187 (
            .O(N__68718),
            .I(\pid_side.error_cry_1_0 ));
    InMux I__15186 (
            .O(N__68715),
            .I(N__68712));
    LocalMux I__15185 (
            .O(N__68712),
            .I(drone_H_disp_side_i_7));
    CascadeMux I__15184 (
            .O(N__68709),
            .I(N__68706));
    InMux I__15183 (
            .O(N__68706),
            .I(N__68703));
    LocalMux I__15182 (
            .O(N__68703),
            .I(side_command_3));
    InMux I__15181 (
            .O(N__68700),
            .I(\pid_side.error_cry_2_0 ));
    InMux I__15180 (
            .O(N__68697),
            .I(N__68694));
    LocalMux I__15179 (
            .O(N__68694),
            .I(N__68689));
    InMux I__15178 (
            .O(N__68693),
            .I(N__68686));
    InMux I__15177 (
            .O(N__68692),
            .I(N__68683));
    Span4Mux_h I__15176 (
            .O(N__68689),
            .I(N__68678));
    LocalMux I__15175 (
            .O(N__68686),
            .I(N__68678));
    LocalMux I__15174 (
            .O(N__68683),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    Odrv4 I__15173 (
            .O(N__68678),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    InMux I__15172 (
            .O(N__68673),
            .I(N__68670));
    LocalMux I__15171 (
            .O(N__68670),
            .I(N__68667));
    Span4Mux_h I__15170 (
            .O(N__68667),
            .I(N__68663));
    InMux I__15169 (
            .O(N__68666),
            .I(N__68660));
    Odrv4 I__15168 (
            .O(N__68663),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    LocalMux I__15167 (
            .O(N__68660),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    CascadeMux I__15166 (
            .O(N__68655),
            .I(N__68651));
    CascadeMux I__15165 (
            .O(N__68654),
            .I(N__68648));
    InMux I__15164 (
            .O(N__68651),
            .I(N__68643));
    InMux I__15163 (
            .O(N__68648),
            .I(N__68643));
    LocalMux I__15162 (
            .O(N__68643),
            .I(N__68640));
    Span4Mux_v I__15161 (
            .O(N__68640),
            .I(N__68633));
    InMux I__15160 (
            .O(N__68639),
            .I(N__68627));
    InMux I__15159 (
            .O(N__68638),
            .I(N__68627));
    InMux I__15158 (
            .O(N__68637),
            .I(N__68622));
    InMux I__15157 (
            .O(N__68636),
            .I(N__68622));
    Span4Mux_h I__15156 (
            .O(N__68633),
            .I(N__68619));
    InMux I__15155 (
            .O(N__68632),
            .I(N__68616));
    LocalMux I__15154 (
            .O(N__68627),
            .I(N__68613));
    LocalMux I__15153 (
            .O(N__68622),
            .I(N__68610));
    Span4Mux_h I__15152 (
            .O(N__68619),
            .I(N__68605));
    LocalMux I__15151 (
            .O(N__68616),
            .I(N__68605));
    Span12Mux_v I__15150 (
            .O(N__68613),
            .I(N__68600));
    Span12Mux_v I__15149 (
            .O(N__68610),
            .I(N__68600));
    Span4Mux_h I__15148 (
            .O(N__68605),
            .I(N__68597));
    Odrv12 I__15147 (
            .O(N__68600),
            .I(uart_drone_data_5));
    Odrv4 I__15146 (
            .O(N__68597),
            .I(uart_drone_data_5));
    InMux I__15145 (
            .O(N__68592),
            .I(N__68586));
    InMux I__15144 (
            .O(N__68591),
            .I(N__68586));
    LocalMux I__15143 (
            .O(N__68586),
            .I(\dron_frame_decoder_1.drone_H_disp_side_5 ));
    InMux I__15142 (
            .O(N__68583),
            .I(N__68577));
    InMux I__15141 (
            .O(N__68582),
            .I(N__68577));
    LocalMux I__15140 (
            .O(N__68577),
            .I(drone_H_disp_side_2));
    CascadeMux I__15139 (
            .O(N__68574),
            .I(N__68570));
    InMux I__15138 (
            .O(N__68573),
            .I(N__68565));
    InMux I__15137 (
            .O(N__68570),
            .I(N__68565));
    LocalMux I__15136 (
            .O(N__68565),
            .I(N__68558));
    CascadeMux I__15135 (
            .O(N__68564),
            .I(N__68555));
    InMux I__15134 (
            .O(N__68563),
            .I(N__68552));
    InMux I__15133 (
            .O(N__68562),
            .I(N__68547));
    InMux I__15132 (
            .O(N__68561),
            .I(N__68547));
    Span4Mux_v I__15131 (
            .O(N__68558),
            .I(N__68544));
    InMux I__15130 (
            .O(N__68555),
            .I(N__68539));
    LocalMux I__15129 (
            .O(N__68552),
            .I(N__68536));
    LocalMux I__15128 (
            .O(N__68547),
            .I(N__68533));
    Span4Mux_h I__15127 (
            .O(N__68544),
            .I(N__68530));
    InMux I__15126 (
            .O(N__68543),
            .I(N__68525));
    InMux I__15125 (
            .O(N__68542),
            .I(N__68525));
    LocalMux I__15124 (
            .O(N__68539),
            .I(N__68522));
    Span4Mux_v I__15123 (
            .O(N__68536),
            .I(N__68519));
    Span12Mux_h I__15122 (
            .O(N__68533),
            .I(N__68516));
    Span4Mux_v I__15121 (
            .O(N__68530),
            .I(N__68511));
    LocalMux I__15120 (
            .O(N__68525),
            .I(N__68511));
    Span12Mux_h I__15119 (
            .O(N__68522),
            .I(N__68508));
    Span4Mux_h I__15118 (
            .O(N__68519),
            .I(N__68505));
    Span12Mux_v I__15117 (
            .O(N__68516),
            .I(N__68502));
    Span4Mux_h I__15116 (
            .O(N__68511),
            .I(N__68499));
    Odrv12 I__15115 (
            .O(N__68508),
            .I(uart_drone_data_6));
    Odrv4 I__15114 (
            .O(N__68505),
            .I(uart_drone_data_6));
    Odrv12 I__15113 (
            .O(N__68502),
            .I(uart_drone_data_6));
    Odrv4 I__15112 (
            .O(N__68499),
            .I(uart_drone_data_6));
    InMux I__15111 (
            .O(N__68490),
            .I(N__68484));
    InMux I__15110 (
            .O(N__68489),
            .I(N__68484));
    LocalMux I__15109 (
            .O(N__68484),
            .I(\dron_frame_decoder_1.drone_H_disp_side_6 ));
    CascadeMux I__15108 (
            .O(N__68481),
            .I(\pid_side.un1_pid_prereg_0_9_cascade_ ));
    InMux I__15107 (
            .O(N__68478),
            .I(N__68475));
    LocalMux I__15106 (
            .O(N__68475),
            .I(N__68472));
    Span4Mux_h I__15105 (
            .O(N__68472),
            .I(N__68468));
    InMux I__15104 (
            .O(N__68471),
            .I(N__68465));
    Odrv4 I__15103 (
            .O(N__68468),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    LocalMux I__15102 (
            .O(N__68465),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    CascadeMux I__15101 (
            .O(N__68460),
            .I(N__68457));
    InMux I__15100 (
            .O(N__68457),
            .I(N__68454));
    LocalMux I__15099 (
            .O(N__68454),
            .I(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ));
    InMux I__15098 (
            .O(N__68451),
            .I(N__68447));
    CascadeMux I__15097 (
            .O(N__68450),
            .I(N__68444));
    LocalMux I__15096 (
            .O(N__68447),
            .I(N__68441));
    InMux I__15095 (
            .O(N__68444),
            .I(N__68438));
    Span4Mux_v I__15094 (
            .O(N__68441),
            .I(N__68433));
    LocalMux I__15093 (
            .O(N__68438),
            .I(N__68433));
    Span4Mux_v I__15092 (
            .O(N__68433),
            .I(N__68430));
    Odrv4 I__15091 (
            .O(N__68430),
            .I(\pid_side.un1_pid_prereg_0 ));
    InMux I__15090 (
            .O(N__68427),
            .I(N__68424));
    LocalMux I__15089 (
            .O(N__68424),
            .I(N__68421));
    Span4Mux_h I__15088 (
            .O(N__68421),
            .I(N__68418));
    Odrv4 I__15087 (
            .O(N__68418),
            .I(\pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ));
    InMux I__15086 (
            .O(N__68415),
            .I(N__68411));
    CascadeMux I__15085 (
            .O(N__68414),
            .I(N__68408));
    LocalMux I__15084 (
            .O(N__68411),
            .I(N__68405));
    InMux I__15083 (
            .O(N__68408),
            .I(N__68402));
    Span4Mux_h I__15082 (
            .O(N__68405),
            .I(N__68399));
    LocalMux I__15081 (
            .O(N__68402),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    Odrv4 I__15080 (
            .O(N__68399),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    CascadeMux I__15079 (
            .O(N__68394),
            .I(N__68391));
    InMux I__15078 (
            .O(N__68391),
            .I(N__68387));
    InMux I__15077 (
            .O(N__68390),
            .I(N__68384));
    LocalMux I__15076 (
            .O(N__68387),
            .I(N__68381));
    LocalMux I__15075 (
            .O(N__68384),
            .I(N__68376));
    Span4Mux_h I__15074 (
            .O(N__68381),
            .I(N__68376));
    Span4Mux_h I__15073 (
            .O(N__68376),
            .I(N__68373));
    Odrv4 I__15072 (
            .O(N__68373),
            .I(\pid_side.error_i_acumm_preregZ0Z_17 ));
    CascadeMux I__15071 (
            .O(N__68370),
            .I(\pid_side.un10lto27_10_cascade_ ));
    InMux I__15070 (
            .O(N__68367),
            .I(N__68364));
    LocalMux I__15069 (
            .O(N__68364),
            .I(N__68361));
    Odrv12 I__15068 (
            .O(N__68361),
            .I(\pid_side.un10lto27_11 ));
    InMux I__15067 (
            .O(N__68358),
            .I(N__68355));
    LocalMux I__15066 (
            .O(N__68355),
            .I(N__68352));
    Span4Mux_h I__15065 (
            .O(N__68352),
            .I(N__68349));
    Odrv4 I__15064 (
            .O(N__68349),
            .I(\pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ));
    CascadeMux I__15063 (
            .O(N__68346),
            .I(N__68343));
    InMux I__15062 (
            .O(N__68343),
            .I(N__68339));
    CascadeMux I__15061 (
            .O(N__68342),
            .I(N__68336));
    LocalMux I__15060 (
            .O(N__68339),
            .I(N__68333));
    InMux I__15059 (
            .O(N__68336),
            .I(N__68330));
    Span4Mux_h I__15058 (
            .O(N__68333),
            .I(N__68327));
    LocalMux I__15057 (
            .O(N__68330),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__15056 (
            .O(N__68327),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    InMux I__15055 (
            .O(N__68322),
            .I(N__68319));
    LocalMux I__15054 (
            .O(N__68319),
            .I(\pid_side.un10lto27_9 ));
    InMux I__15053 (
            .O(N__68316),
            .I(N__68309));
    InMux I__15052 (
            .O(N__68315),
            .I(N__68309));
    InMux I__15051 (
            .O(N__68314),
            .I(N__68306));
    LocalMux I__15050 (
            .O(N__68309),
            .I(N__68303));
    LocalMux I__15049 (
            .O(N__68306),
            .I(N__68300));
    Span4Mux_h I__15048 (
            .O(N__68303),
            .I(N__68297));
    Odrv4 I__15047 (
            .O(N__68300),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    Odrv4 I__15046 (
            .O(N__68297),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    InMux I__15045 (
            .O(N__68292),
            .I(N__68289));
    LocalMux I__15044 (
            .O(N__68289),
            .I(N__68285));
    InMux I__15043 (
            .O(N__68288),
            .I(N__68282));
    Odrv12 I__15042 (
            .O(N__68285),
            .I(\pid_side.error_i_acumm_preregZ0Z_18 ));
    LocalMux I__15041 (
            .O(N__68282),
            .I(\pid_side.error_i_acumm_preregZ0Z_18 ));
    InMux I__15040 (
            .O(N__68277),
            .I(N__68273));
    InMux I__15039 (
            .O(N__68276),
            .I(N__68270));
    LocalMux I__15038 (
            .O(N__68273),
            .I(N__68264));
    LocalMux I__15037 (
            .O(N__68270),
            .I(N__68264));
    InMux I__15036 (
            .O(N__68269),
            .I(N__68261));
    Span4Mux_v I__15035 (
            .O(N__68264),
            .I(N__68256));
    LocalMux I__15034 (
            .O(N__68261),
            .I(N__68256));
    Span4Mux_h I__15033 (
            .O(N__68256),
            .I(N__68253));
    Odrv4 I__15032 (
            .O(N__68253),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    InMux I__15031 (
            .O(N__68250),
            .I(N__68247));
    LocalMux I__15030 (
            .O(N__68247),
            .I(N__68243));
    InMux I__15029 (
            .O(N__68246),
            .I(N__68240));
    Odrv12 I__15028 (
            .O(N__68243),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__15027 (
            .O(N__68240),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    InMux I__15026 (
            .O(N__68235),
            .I(N__68232));
    LocalMux I__15025 (
            .O(N__68232),
            .I(N__68228));
    InMux I__15024 (
            .O(N__68231),
            .I(N__68225));
    Odrv12 I__15023 (
            .O(N__68228),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__15022 (
            .O(N__68225),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    InMux I__15021 (
            .O(N__68220),
            .I(N__68216));
    InMux I__15020 (
            .O(N__68219),
            .I(N__68213));
    LocalMux I__15019 (
            .O(N__68216),
            .I(N__68209));
    LocalMux I__15018 (
            .O(N__68213),
            .I(N__68206));
    InMux I__15017 (
            .O(N__68212),
            .I(N__68203));
    Span4Mux_h I__15016 (
            .O(N__68209),
            .I(N__68200));
    Odrv4 I__15015 (
            .O(N__68206),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    LocalMux I__15014 (
            .O(N__68203),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    Odrv4 I__15013 (
            .O(N__68200),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    InMux I__15012 (
            .O(N__68193),
            .I(N__68190));
    LocalMux I__15011 (
            .O(N__68190),
            .I(N__68186));
    InMux I__15010 (
            .O(N__68189),
            .I(N__68183));
    Odrv12 I__15009 (
            .O(N__68186),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__15008 (
            .O(N__68183),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    CascadeMux I__15007 (
            .O(N__68178),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10_cascade_ ));
    CascadeMux I__15006 (
            .O(N__68175),
            .I(N__68172));
    InMux I__15005 (
            .O(N__68172),
            .I(N__68169));
    LocalMux I__15004 (
            .O(N__68169),
            .I(N__68166));
    Span4Mux_h I__15003 (
            .O(N__68166),
            .I(N__68162));
    InMux I__15002 (
            .O(N__68165),
            .I(N__68159));
    Odrv4 I__15001 (
            .O(N__68162),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    LocalMux I__15000 (
            .O(N__68159),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    InMux I__14999 (
            .O(N__68154),
            .I(N__68144));
    InMux I__14998 (
            .O(N__68153),
            .I(N__68144));
    InMux I__14997 (
            .O(N__68152),
            .I(N__68144));
    InMux I__14996 (
            .O(N__68151),
            .I(N__68141));
    LocalMux I__14995 (
            .O(N__68144),
            .I(N__68138));
    LocalMux I__14994 (
            .O(N__68141),
            .I(N__68133));
    Span4Mux_h I__14993 (
            .O(N__68138),
            .I(N__68133));
    Odrv4 I__14992 (
            .O(N__68133),
            .I(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ));
    InMux I__14991 (
            .O(N__68130),
            .I(N__68124));
    InMux I__14990 (
            .O(N__68129),
            .I(N__68124));
    LocalMux I__14989 (
            .O(N__68124),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    InMux I__14988 (
            .O(N__68121),
            .I(N__68118));
    LocalMux I__14987 (
            .O(N__68118),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ));
    InMux I__14986 (
            .O(N__68115),
            .I(N__68110));
    InMux I__14985 (
            .O(N__68114),
            .I(N__68107));
    InMux I__14984 (
            .O(N__68113),
            .I(N__68104));
    LocalMux I__14983 (
            .O(N__68110),
            .I(N__68101));
    LocalMux I__14982 (
            .O(N__68107),
            .I(N__68098));
    LocalMux I__14981 (
            .O(N__68104),
            .I(N__68095));
    Span4Mux_v I__14980 (
            .O(N__68101),
            .I(N__68092));
    Span4Mux_h I__14979 (
            .O(N__68098),
            .I(N__68087));
    Span4Mux_v I__14978 (
            .O(N__68095),
            .I(N__68087));
    Odrv4 I__14977 (
            .O(N__68092),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    Odrv4 I__14976 (
            .O(N__68087),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    CascadeMux I__14975 (
            .O(N__68082),
            .I(\pid_side.un1_pid_prereg_9_0_cascade_ ));
    CascadeMux I__14974 (
            .O(N__68079),
            .I(N__68076));
    InMux I__14973 (
            .O(N__68076),
            .I(N__68073));
    LocalMux I__14972 (
            .O(N__68073),
            .I(N__68070));
    Odrv4 I__14971 (
            .O(N__68070),
            .I(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ));
    InMux I__14970 (
            .O(N__68067),
            .I(N__68064));
    LocalMux I__14969 (
            .O(N__68064),
            .I(N__68060));
    InMux I__14968 (
            .O(N__68063),
            .I(N__68057));
    Odrv4 I__14967 (
            .O(N__68060),
            .I(\pid_side.un1_pid_prereg_0_7 ));
    LocalMux I__14966 (
            .O(N__68057),
            .I(\pid_side.un1_pid_prereg_0_7 ));
    InMux I__14965 (
            .O(N__68052),
            .I(N__68049));
    LocalMux I__14964 (
            .O(N__68049),
            .I(N__68045));
    InMux I__14963 (
            .O(N__68048),
            .I(N__68042));
    Odrv4 I__14962 (
            .O(N__68045),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    LocalMux I__14961 (
            .O(N__68042),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    CascadeMux I__14960 (
            .O(N__68037),
            .I(\pid_side.un1_pid_prereg_0_8_cascade_ ));
    CascadeMux I__14959 (
            .O(N__68034),
            .I(N__68031));
    InMux I__14958 (
            .O(N__68031),
            .I(N__68028));
    LocalMux I__14957 (
            .O(N__68028),
            .I(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ));
    InMux I__14956 (
            .O(N__68025),
            .I(N__68022));
    LocalMux I__14955 (
            .O(N__68022),
            .I(N__68019));
    Span4Mux_v I__14954 (
            .O(N__68019),
            .I(N__68015));
    InMux I__14953 (
            .O(N__68018),
            .I(N__68012));
    Odrv4 I__14952 (
            .O(N__68015),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    LocalMux I__14951 (
            .O(N__68012),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    CascadeMux I__14950 (
            .O(N__68007),
            .I(\pid_side.un1_pid_prereg_0_7_cascade_ ));
    InMux I__14949 (
            .O(N__68004),
            .I(N__68001));
    LocalMux I__14948 (
            .O(N__68001),
            .I(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ));
    InMux I__14947 (
            .O(N__67998),
            .I(N__67993));
    InMux I__14946 (
            .O(N__67997),
            .I(N__67990));
    InMux I__14945 (
            .O(N__67996),
            .I(N__67987));
    LocalMux I__14944 (
            .O(N__67993),
            .I(N__67984));
    LocalMux I__14943 (
            .O(N__67990),
            .I(N__67979));
    LocalMux I__14942 (
            .O(N__67987),
            .I(N__67979));
    Span4Mux_h I__14941 (
            .O(N__67984),
            .I(N__67976));
    Span4Mux_h I__14940 (
            .O(N__67979),
            .I(N__67973));
    Odrv4 I__14939 (
            .O(N__67976),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    Odrv4 I__14938 (
            .O(N__67973),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    InMux I__14937 (
            .O(N__67968),
            .I(N__67959));
    InMux I__14936 (
            .O(N__67967),
            .I(N__67959));
    InMux I__14935 (
            .O(N__67966),
            .I(N__67959));
    LocalMux I__14934 (
            .O(N__67959),
            .I(\pid_side.un1_pid_prereg_0_4 ));
    InMux I__14933 (
            .O(N__67956),
            .I(N__67953));
    LocalMux I__14932 (
            .O(N__67953),
            .I(N__67949));
    InMux I__14931 (
            .O(N__67952),
            .I(N__67946));
    Odrv4 I__14930 (
            .O(N__67949),
            .I(\pid_side.error_d_reg_prev_esr_RNI83KO4Z0Z_12 ));
    LocalMux I__14929 (
            .O(N__67946),
            .I(\pid_side.error_d_reg_prev_esr_RNI83KO4Z0Z_12 ));
    CascadeMux I__14928 (
            .O(N__67941),
            .I(N__67938));
    InMux I__14927 (
            .O(N__67938),
            .I(N__67935));
    LocalMux I__14926 (
            .O(N__67935),
            .I(\pid_side.error_d_reg_prev_esr_RNI3AMCBZ0Z_10 ));
    InMux I__14925 (
            .O(N__67932),
            .I(N__67927));
    InMux I__14924 (
            .O(N__67931),
            .I(N__67922));
    InMux I__14923 (
            .O(N__67930),
            .I(N__67922));
    LocalMux I__14922 (
            .O(N__67927),
            .I(N__67919));
    LocalMux I__14921 (
            .O(N__67922),
            .I(N__67916));
    Span4Mux_h I__14920 (
            .O(N__67919),
            .I(N__67911));
    Span4Mux_h I__14919 (
            .O(N__67916),
            .I(N__67911));
    Odrv4 I__14918 (
            .O(N__67911),
            .I(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ));
    CascadeMux I__14917 (
            .O(N__67908),
            .I(\pid_side.un1_pid_prereg_153_0_cascade_ ));
    CascadeMux I__14916 (
            .O(N__67905),
            .I(N__67902));
    InMux I__14915 (
            .O(N__67902),
            .I(N__67899));
    LocalMux I__14914 (
            .O(N__67899),
            .I(\pid_side.error_d_reg_prev_esr_RNIO56DBZ0Z_10 ));
    CascadeMux I__14913 (
            .O(N__67896),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ));
    InMux I__14912 (
            .O(N__67893),
            .I(N__67887));
    InMux I__14911 (
            .O(N__67892),
            .I(N__67887));
    LocalMux I__14910 (
            .O(N__67887),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ));
    InMux I__14909 (
            .O(N__67884),
            .I(N__67881));
    LocalMux I__14908 (
            .O(N__67881),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ));
    InMux I__14907 (
            .O(N__67878),
            .I(N__67872));
    InMux I__14906 (
            .O(N__67877),
            .I(N__67872));
    LocalMux I__14905 (
            .O(N__67872),
            .I(N__67869));
    Odrv4 I__14904 (
            .O(N__67869),
            .I(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ));
    CascadeMux I__14903 (
            .O(N__67866),
            .I(N__67863));
    InMux I__14902 (
            .O(N__67863),
            .I(N__67858));
    InMux I__14901 (
            .O(N__67862),
            .I(N__67855));
    CascadeMux I__14900 (
            .O(N__67861),
            .I(N__67852));
    LocalMux I__14899 (
            .O(N__67858),
            .I(N__67849));
    LocalMux I__14898 (
            .O(N__67855),
            .I(N__67846));
    InMux I__14897 (
            .O(N__67852),
            .I(N__67843));
    Span4Mux_h I__14896 (
            .O(N__67849),
            .I(N__67836));
    Span4Mux_h I__14895 (
            .O(N__67846),
            .I(N__67836));
    LocalMux I__14894 (
            .O(N__67843),
            .I(N__67836));
    Span4Mux_v I__14893 (
            .O(N__67836),
            .I(N__67833));
    Odrv4 I__14892 (
            .O(N__67833),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    InMux I__14891 (
            .O(N__67830),
            .I(N__67827));
    LocalMux I__14890 (
            .O(N__67827),
            .I(N__67823));
    InMux I__14889 (
            .O(N__67826),
            .I(N__67820));
    Odrv4 I__14888 (
            .O(N__67823),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    LocalMux I__14887 (
            .O(N__67820),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    CascadeMux I__14886 (
            .O(N__67815),
            .I(N__67812));
    InMux I__14885 (
            .O(N__67812),
            .I(N__67809));
    LocalMux I__14884 (
            .O(N__67809),
            .I(N__67805));
    InMux I__14883 (
            .O(N__67808),
            .I(N__67802));
    Odrv4 I__14882 (
            .O(N__67805),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    LocalMux I__14881 (
            .O(N__67802),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    InMux I__14880 (
            .O(N__67797),
            .I(N__67794));
    LocalMux I__14879 (
            .O(N__67794),
            .I(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ));
    CascadeMux I__14878 (
            .O(N__67791),
            .I(\pid_side.un1_pid_prereg_0_5_cascade_ ));
    CascadeMux I__14877 (
            .O(N__67788),
            .I(N__67785));
    InMux I__14876 (
            .O(N__67785),
            .I(N__67782));
    LocalMux I__14875 (
            .O(N__67782),
            .I(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ));
    InMux I__14874 (
            .O(N__67779),
            .I(N__67773));
    InMux I__14873 (
            .O(N__67778),
            .I(N__67773));
    LocalMux I__14872 (
            .O(N__67773),
            .I(\pid_side.un1_pid_prereg_0_5 ));
    CascadeMux I__14871 (
            .O(N__67770),
            .I(\pid_side.un1_pid_prereg_0_6_cascade_ ));
    InMux I__14870 (
            .O(N__67767),
            .I(N__67764));
    LocalMux I__14869 (
            .O(N__67764),
            .I(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ));
    CascadeMux I__14868 (
            .O(N__67761),
            .I(N__67753));
    CascadeMux I__14867 (
            .O(N__67760),
            .I(N__67749));
    CascadeMux I__14866 (
            .O(N__67759),
            .I(N__67746));
    CascadeMux I__14865 (
            .O(N__67758),
            .I(N__67743));
    InMux I__14864 (
            .O(N__67757),
            .I(N__67732));
    InMux I__14863 (
            .O(N__67756),
            .I(N__67732));
    InMux I__14862 (
            .O(N__67753),
            .I(N__67732));
    InMux I__14861 (
            .O(N__67752),
            .I(N__67732));
    InMux I__14860 (
            .O(N__67749),
            .I(N__67718));
    InMux I__14859 (
            .O(N__67746),
            .I(N__67718));
    InMux I__14858 (
            .O(N__67743),
            .I(N__67718));
    InMux I__14857 (
            .O(N__67742),
            .I(N__67718));
    InMux I__14856 (
            .O(N__67741),
            .I(N__67718));
    LocalMux I__14855 (
            .O(N__67732),
            .I(N__67715));
    InMux I__14854 (
            .O(N__67731),
            .I(N__67708));
    InMux I__14853 (
            .O(N__67730),
            .I(N__67708));
    InMux I__14852 (
            .O(N__67729),
            .I(N__67708));
    LocalMux I__14851 (
            .O(N__67718),
            .I(N__67703));
    Span4Mux_h I__14850 (
            .O(N__67715),
            .I(N__67703));
    LocalMux I__14849 (
            .O(N__67708),
            .I(\pid_side.N_76 ));
    Odrv4 I__14848 (
            .O(N__67703),
            .I(\pid_side.N_76 ));
    InMux I__14847 (
            .O(N__67698),
            .I(N__67695));
    LocalMux I__14846 (
            .O(N__67695),
            .I(N__67690));
    InMux I__14845 (
            .O(N__67694),
            .I(N__67685));
    InMux I__14844 (
            .O(N__67693),
            .I(N__67685));
    Span4Mux_v I__14843 (
            .O(N__67690),
            .I(N__67682));
    LocalMux I__14842 (
            .O(N__67685),
            .I(N__67679));
    Odrv4 I__14841 (
            .O(N__67682),
            .I(\pid_side.pid_preregZ0Z_9 ));
    Odrv4 I__14840 (
            .O(N__67679),
            .I(\pid_side.pid_preregZ0Z_9 ));
    InMux I__14839 (
            .O(N__67674),
            .I(N__67670));
    InMux I__14838 (
            .O(N__67673),
            .I(N__67667));
    LocalMux I__14837 (
            .O(N__67670),
            .I(N__67662));
    LocalMux I__14836 (
            .O(N__67667),
            .I(N__67662));
    Span4Mux_h I__14835 (
            .O(N__67662),
            .I(N__67659));
    Odrv4 I__14834 (
            .O(N__67659),
            .I(side_order_9));
    CascadeMux I__14833 (
            .O(N__67656),
            .I(N__67652));
    InMux I__14832 (
            .O(N__67655),
            .I(N__67636));
    InMux I__14831 (
            .O(N__67652),
            .I(N__67636));
    InMux I__14830 (
            .O(N__67651),
            .I(N__67636));
    CascadeMux I__14829 (
            .O(N__67650),
            .I(N__67633));
    CascadeMux I__14828 (
            .O(N__67649),
            .I(N__67628));
    InMux I__14827 (
            .O(N__67648),
            .I(N__67620));
    InMux I__14826 (
            .O(N__67647),
            .I(N__67609));
    InMux I__14825 (
            .O(N__67646),
            .I(N__67609));
    InMux I__14824 (
            .O(N__67645),
            .I(N__67609));
    InMux I__14823 (
            .O(N__67644),
            .I(N__67609));
    InMux I__14822 (
            .O(N__67643),
            .I(N__67609));
    LocalMux I__14821 (
            .O(N__67636),
            .I(N__67606));
    InMux I__14820 (
            .O(N__67633),
            .I(N__67599));
    InMux I__14819 (
            .O(N__67632),
            .I(N__67599));
    InMux I__14818 (
            .O(N__67631),
            .I(N__67599));
    InMux I__14817 (
            .O(N__67628),
            .I(N__67586));
    InMux I__14816 (
            .O(N__67627),
            .I(N__67586));
    InMux I__14815 (
            .O(N__67626),
            .I(N__67586));
    InMux I__14814 (
            .O(N__67625),
            .I(N__67586));
    InMux I__14813 (
            .O(N__67624),
            .I(N__67586));
    InMux I__14812 (
            .O(N__67623),
            .I(N__67586));
    LocalMux I__14811 (
            .O(N__67620),
            .I(N__67583));
    LocalMux I__14810 (
            .O(N__67609),
            .I(N__67580));
    Span4Mux_v I__14809 (
            .O(N__67606),
            .I(N__67573));
    LocalMux I__14808 (
            .O(N__67599),
            .I(N__67573));
    LocalMux I__14807 (
            .O(N__67586),
            .I(N__67573));
    Span4Mux_v I__14806 (
            .O(N__67583),
            .I(N__67570));
    Span4Mux_v I__14805 (
            .O(N__67580),
            .I(N__67565));
    Span4Mux_h I__14804 (
            .O(N__67573),
            .I(N__67565));
    Odrv4 I__14803 (
            .O(N__67570),
            .I(\pid_side.pid_preregZ0Z_30 ));
    Odrv4 I__14802 (
            .O(N__67565),
            .I(\pid_side.pid_preregZ0Z_30 ));
    InMux I__14801 (
            .O(N__67560),
            .I(N__67556));
    CascadeMux I__14800 (
            .O(N__67559),
            .I(N__67553));
    LocalMux I__14799 (
            .O(N__67556),
            .I(N__67550));
    InMux I__14798 (
            .O(N__67553),
            .I(N__67547));
    Span4Mux_h I__14797 (
            .O(N__67550),
            .I(N__67542));
    LocalMux I__14796 (
            .O(N__67547),
            .I(N__67539));
    InMux I__14795 (
            .O(N__67546),
            .I(N__67534));
    InMux I__14794 (
            .O(N__67545),
            .I(N__67534));
    Odrv4 I__14793 (
            .O(N__67542),
            .I(\pid_side.N_98 ));
    Odrv4 I__14792 (
            .O(N__67539),
            .I(\pid_side.N_98 ));
    LocalMux I__14791 (
            .O(N__67534),
            .I(\pid_side.N_98 ));
    InMux I__14790 (
            .O(N__67527),
            .I(N__67520));
    InMux I__14789 (
            .O(N__67526),
            .I(N__67520));
    InMux I__14788 (
            .O(N__67525),
            .I(N__67514));
    LocalMux I__14787 (
            .O(N__67520),
            .I(N__67511));
    InMux I__14786 (
            .O(N__67519),
            .I(N__67506));
    InMux I__14785 (
            .O(N__67518),
            .I(N__67506));
    InMux I__14784 (
            .O(N__67517),
            .I(N__67503));
    LocalMux I__14783 (
            .O(N__67514),
            .I(N__67500));
    Span4Mux_h I__14782 (
            .O(N__67511),
            .I(N__67497));
    LocalMux I__14781 (
            .O(N__67506),
            .I(N__67492));
    LocalMux I__14780 (
            .O(N__67503),
            .I(N__67492));
    Odrv4 I__14779 (
            .O(N__67500),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__14778 (
            .O(N__67497),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__14777 (
            .O(N__67492),
            .I(\pid_side.pid_preregZ0Z_13 ));
    CascadeMux I__14776 (
            .O(N__67485),
            .I(N__67482));
    InMux I__14775 (
            .O(N__67482),
            .I(N__67479));
    LocalMux I__14774 (
            .O(N__67479),
            .I(N__67475));
    InMux I__14773 (
            .O(N__67478),
            .I(N__67472));
    Span4Mux_v I__14772 (
            .O(N__67475),
            .I(N__67467));
    LocalMux I__14771 (
            .O(N__67472),
            .I(N__67467));
    Span4Mux_h I__14770 (
            .O(N__67467),
            .I(N__67464));
    Odrv4 I__14769 (
            .O(N__67464),
            .I(side_order_13));
    CEMux I__14768 (
            .O(N__67461),
            .I(N__67458));
    LocalMux I__14767 (
            .O(N__67458),
            .I(N__67454));
    CEMux I__14766 (
            .O(N__67457),
            .I(N__67451));
    Span4Mux_h I__14765 (
            .O(N__67454),
            .I(N__67446));
    LocalMux I__14764 (
            .O(N__67451),
            .I(N__67446));
    Span4Mux_h I__14763 (
            .O(N__67446),
            .I(N__67441));
    CEMux I__14762 (
            .O(N__67445),
            .I(N__67438));
    CEMux I__14761 (
            .O(N__67444),
            .I(N__67435));
    Odrv4 I__14760 (
            .O(N__67441),
            .I(\pid_side.state_0_1 ));
    LocalMux I__14759 (
            .O(N__67438),
            .I(\pid_side.state_0_1 ));
    LocalMux I__14758 (
            .O(N__67435),
            .I(\pid_side.state_0_1 ));
    SRMux I__14757 (
            .O(N__67428),
            .I(N__67422));
    SRMux I__14756 (
            .O(N__67427),
            .I(N__67419));
    SRMux I__14755 (
            .O(N__67426),
            .I(N__67416));
    SRMux I__14754 (
            .O(N__67425),
            .I(N__67413));
    LocalMux I__14753 (
            .O(N__67422),
            .I(N__67410));
    LocalMux I__14752 (
            .O(N__67419),
            .I(N__67405));
    LocalMux I__14751 (
            .O(N__67416),
            .I(N__67405));
    LocalMux I__14750 (
            .O(N__67413),
            .I(N__67398));
    Span4Mux_v I__14749 (
            .O(N__67410),
            .I(N__67398));
    Span4Mux_h I__14748 (
            .O(N__67405),
            .I(N__67398));
    Span4Mux_h I__14747 (
            .O(N__67398),
            .I(N__67395));
    Odrv4 I__14746 (
            .O(N__67395),
            .I(\pid_side.un1_reset_0_i ));
    CascadeMux I__14745 (
            .O(N__67392),
            .I(\pid_side.state_RNINK4UZ0Z_0_cascade_ ));
    IoInMux I__14744 (
            .O(N__67389),
            .I(N__67386));
    LocalMux I__14743 (
            .O(N__67386),
            .I(N__67383));
    Span4Mux_s2_v I__14742 (
            .O(N__67383),
            .I(N__67380));
    Span4Mux_v I__14741 (
            .O(N__67380),
            .I(N__67374));
    InMux I__14740 (
            .O(N__67379),
            .I(N__67371));
    InMux I__14739 (
            .O(N__67378),
            .I(N__67364));
    InMux I__14738 (
            .O(N__67377),
            .I(N__67361));
    Span4Mux_v I__14737 (
            .O(N__67374),
            .I(N__67356));
    LocalMux I__14736 (
            .O(N__67371),
            .I(N__67356));
    InMux I__14735 (
            .O(N__67370),
            .I(N__67353));
    InMux I__14734 (
            .O(N__67369),
            .I(N__67348));
    InMux I__14733 (
            .O(N__67368),
            .I(N__67348));
    InMux I__14732 (
            .O(N__67367),
            .I(N__67345));
    LocalMux I__14731 (
            .O(N__67364),
            .I(N__67339));
    LocalMux I__14730 (
            .O(N__67361),
            .I(N__67334));
    Span4Mux_h I__14729 (
            .O(N__67356),
            .I(N__67334));
    LocalMux I__14728 (
            .O(N__67353),
            .I(N__67329));
    LocalMux I__14727 (
            .O(N__67348),
            .I(N__67329));
    LocalMux I__14726 (
            .O(N__67345),
            .I(N__67326));
    InMux I__14725 (
            .O(N__67344),
            .I(N__67319));
    InMux I__14724 (
            .O(N__67343),
            .I(N__67319));
    InMux I__14723 (
            .O(N__67342),
            .I(N__67319));
    Span4Mux_v I__14722 (
            .O(N__67339),
            .I(N__67316));
    Span4Mux_v I__14721 (
            .O(N__67334),
            .I(N__67313));
    Span4Mux_h I__14720 (
            .O(N__67329),
            .I(N__67309));
    Span4Mux_v I__14719 (
            .O(N__67326),
            .I(N__67304));
    LocalMux I__14718 (
            .O(N__67319),
            .I(N__67304));
    Span4Mux_h I__14717 (
            .O(N__67316),
            .I(N__67299));
    Span4Mux_v I__14716 (
            .O(N__67313),
            .I(N__67299));
    InMux I__14715 (
            .O(N__67312),
            .I(N__67296));
    Span4Mux_v I__14714 (
            .O(N__67309),
            .I(N__67293));
    Span4Mux_v I__14713 (
            .O(N__67304),
            .I(N__67288));
    Span4Mux_h I__14712 (
            .O(N__67299),
            .I(N__67288));
    LocalMux I__14711 (
            .O(N__67296),
            .I(debug_CH1_0A_c));
    Odrv4 I__14710 (
            .O(N__67293),
            .I(debug_CH1_0A_c));
    Odrv4 I__14709 (
            .O(N__67288),
            .I(debug_CH1_0A_c));
    InMux I__14708 (
            .O(N__67281),
            .I(N__67274));
    InMux I__14707 (
            .O(N__67280),
            .I(N__67274));
    CascadeMux I__14706 (
            .O(N__67279),
            .I(N__67269));
    LocalMux I__14705 (
            .O(N__67274),
            .I(N__67265));
    InMux I__14704 (
            .O(N__67273),
            .I(N__67262));
    CascadeMux I__14703 (
            .O(N__67272),
            .I(N__67257));
    InMux I__14702 (
            .O(N__67269),
            .I(N__67254));
    InMux I__14701 (
            .O(N__67268),
            .I(N__67251));
    Span4Mux_h I__14700 (
            .O(N__67265),
            .I(N__67248));
    LocalMux I__14699 (
            .O(N__67262),
            .I(N__67245));
    InMux I__14698 (
            .O(N__67261),
            .I(N__67242));
    InMux I__14697 (
            .O(N__67260),
            .I(N__67237));
    InMux I__14696 (
            .O(N__67257),
            .I(N__67237));
    LocalMux I__14695 (
            .O(N__67254),
            .I(N__67232));
    LocalMux I__14694 (
            .O(N__67251),
            .I(N__67232));
    Sp12to4 I__14693 (
            .O(N__67248),
            .I(N__67227));
    Span12Mux_s6_v I__14692 (
            .O(N__67245),
            .I(N__67227));
    LocalMux I__14691 (
            .O(N__67242),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__14690 (
            .O(N__67237),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__14689 (
            .O(N__67232),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv12 I__14688 (
            .O(N__67227),
            .I(\pid_side.stateZ0Z_0 ));
    InMux I__14687 (
            .O(N__67218),
            .I(N__67214));
    InMux I__14686 (
            .O(N__67217),
            .I(N__67211));
    LocalMux I__14685 (
            .O(N__67214),
            .I(N__67208));
    LocalMux I__14684 (
            .O(N__67211),
            .I(N__67205));
    Span4Mux_v I__14683 (
            .O(N__67208),
            .I(N__67202));
    Span4Mux_v I__14682 (
            .O(N__67205),
            .I(N__67199));
    Span4Mux_h I__14681 (
            .O(N__67202),
            .I(N__67196));
    Span4Mux_v I__14680 (
            .O(N__67199),
            .I(N__67191));
    Span4Mux_h I__14679 (
            .O(N__67196),
            .I(N__67191));
    Odrv4 I__14678 (
            .O(N__67191),
            .I(\pid_side.state_ns_0 ));
    InMux I__14677 (
            .O(N__67188),
            .I(N__67182));
    InMux I__14676 (
            .O(N__67187),
            .I(N__67182));
    LocalMux I__14675 (
            .O(N__67182),
            .I(N__67179));
    Span4Mux_h I__14674 (
            .O(N__67179),
            .I(N__67176));
    Span4Mux_v I__14673 (
            .O(N__67176),
            .I(N__67173));
    Odrv4 I__14672 (
            .O(N__67173),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ));
    InMux I__14671 (
            .O(N__67170),
            .I(N__67166));
    CascadeMux I__14670 (
            .O(N__67169),
            .I(N__67162));
    LocalMux I__14669 (
            .O(N__67166),
            .I(N__67159));
    InMux I__14668 (
            .O(N__67165),
            .I(N__67154));
    InMux I__14667 (
            .O(N__67162),
            .I(N__67154));
    Span4Mux_v I__14666 (
            .O(N__67159),
            .I(N__67151));
    LocalMux I__14665 (
            .O(N__67154),
            .I(N__67148));
    Span4Mux_h I__14664 (
            .O(N__67151),
            .I(N__67143));
    Span4Mux_h I__14663 (
            .O(N__67148),
            .I(N__67143));
    Odrv4 I__14662 (
            .O(N__67143),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    CascadeMux I__14661 (
            .O(N__67140),
            .I(N__67133));
    InMux I__14660 (
            .O(N__67139),
            .I(N__67130));
    CascadeMux I__14659 (
            .O(N__67138),
            .I(N__67125));
    CascadeMux I__14658 (
            .O(N__67137),
            .I(N__67122));
    CascadeMux I__14657 (
            .O(N__67136),
            .I(N__67118));
    InMux I__14656 (
            .O(N__67133),
            .I(N__67113));
    LocalMux I__14655 (
            .O(N__67130),
            .I(N__67110));
    InMux I__14654 (
            .O(N__67129),
            .I(N__67095));
    InMux I__14653 (
            .O(N__67128),
            .I(N__67095));
    InMux I__14652 (
            .O(N__67125),
            .I(N__67095));
    InMux I__14651 (
            .O(N__67122),
            .I(N__67095));
    InMux I__14650 (
            .O(N__67121),
            .I(N__67095));
    InMux I__14649 (
            .O(N__67118),
            .I(N__67095));
    InMux I__14648 (
            .O(N__67117),
            .I(N__67095));
    CascadeMux I__14647 (
            .O(N__67116),
            .I(N__67091));
    LocalMux I__14646 (
            .O(N__67113),
            .I(N__67088));
    Span4Mux_v I__14645 (
            .O(N__67110),
            .I(N__67083));
    LocalMux I__14644 (
            .O(N__67095),
            .I(N__67083));
    InMux I__14643 (
            .O(N__67094),
            .I(N__67078));
    InMux I__14642 (
            .O(N__67091),
            .I(N__67078));
    Span4Mux_v I__14641 (
            .O(N__67088),
            .I(N__67069));
    Span4Mux_v I__14640 (
            .O(N__67083),
            .I(N__67069));
    LocalMux I__14639 (
            .O(N__67078),
            .I(N__67069));
    InMux I__14638 (
            .O(N__67077),
            .I(N__67066));
    InMux I__14637 (
            .O(N__67076),
            .I(N__67063));
    Span4Mux_h I__14636 (
            .O(N__67069),
            .I(N__67060));
    LocalMux I__14635 (
            .O(N__67066),
            .I(N__67055));
    LocalMux I__14634 (
            .O(N__67063),
            .I(N__67050));
    Span4Mux_h I__14633 (
            .O(N__67060),
            .I(N__67050));
    InMux I__14632 (
            .O(N__67059),
            .I(N__67045));
    InMux I__14631 (
            .O(N__67058),
            .I(N__67045));
    Odrv4 I__14630 (
            .O(N__67055),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__14629 (
            .O(N__67050),
            .I(\pid_side.stateZ0Z_1 ));
    LocalMux I__14628 (
            .O(N__67045),
            .I(\pid_side.stateZ0Z_1 ));
    InMux I__14627 (
            .O(N__67038),
            .I(N__67026));
    InMux I__14626 (
            .O(N__67037),
            .I(N__67026));
    InMux I__14625 (
            .O(N__67036),
            .I(N__67026));
    InMux I__14624 (
            .O(N__67035),
            .I(N__67026));
    LocalMux I__14623 (
            .O(N__67026),
            .I(N__67023));
    Span4Mux_v I__14622 (
            .O(N__67023),
            .I(N__67020));
    Odrv4 I__14621 (
            .O(N__67020),
            .I(\pid_side.error_i_acumm_3_sqmuxa ));
    InMux I__14620 (
            .O(N__67017),
            .I(N__67014));
    LocalMux I__14619 (
            .O(N__67014),
            .I(\pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ));
    CascadeMux I__14618 (
            .O(N__67011),
            .I(N__67007));
    InMux I__14617 (
            .O(N__67010),
            .I(N__67004));
    InMux I__14616 (
            .O(N__67007),
            .I(N__67001));
    LocalMux I__14615 (
            .O(N__67004),
            .I(N__66996));
    LocalMux I__14614 (
            .O(N__67001),
            .I(N__66996));
    Odrv4 I__14613 (
            .O(N__66996),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    InMux I__14612 (
            .O(N__66993),
            .I(N__66990));
    LocalMux I__14611 (
            .O(N__66990),
            .I(N__66987));
    Odrv4 I__14610 (
            .O(N__66987),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__14609 (
            .O(N__66984),
            .I(N__66980));
    CascadeMux I__14608 (
            .O(N__66983),
            .I(N__66977));
    LocalMux I__14607 (
            .O(N__66980),
            .I(N__66974));
    InMux I__14606 (
            .O(N__66977),
            .I(N__66971));
    Span4Mux_v I__14605 (
            .O(N__66974),
            .I(N__66968));
    LocalMux I__14604 (
            .O(N__66971),
            .I(N__66965));
    Odrv4 I__14603 (
            .O(N__66968),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    Odrv4 I__14602 (
            .O(N__66965),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    InMux I__14601 (
            .O(N__66960),
            .I(N__66957));
    LocalMux I__14600 (
            .O(N__66957),
            .I(N__66954));
    Odrv4 I__14599 (
            .O(N__66954),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    CascadeMux I__14598 (
            .O(N__66951),
            .I(N__66947));
    InMux I__14597 (
            .O(N__66950),
            .I(N__66944));
    InMux I__14596 (
            .O(N__66947),
            .I(N__66941));
    LocalMux I__14595 (
            .O(N__66944),
            .I(N__66936));
    LocalMux I__14594 (
            .O(N__66941),
            .I(N__66936));
    Span4Mux_h I__14593 (
            .O(N__66936),
            .I(N__66933));
    Odrv4 I__14592 (
            .O(N__66933),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    CascadeMux I__14591 (
            .O(N__66930),
            .I(N__66927));
    InMux I__14590 (
            .O(N__66927),
            .I(N__66922));
    InMux I__14589 (
            .O(N__66926),
            .I(N__66917));
    InMux I__14588 (
            .O(N__66925),
            .I(N__66917));
    LocalMux I__14587 (
            .O(N__66922),
            .I(\pid_side.pid_preregZ0Z_1 ));
    LocalMux I__14586 (
            .O(N__66917),
            .I(\pid_side.pid_preregZ0Z_1 ));
    InMux I__14585 (
            .O(N__66912),
            .I(N__66909));
    LocalMux I__14584 (
            .O(N__66909),
            .I(N__66906));
    Span4Mux_h I__14583 (
            .O(N__66906),
            .I(N__66902));
    InMux I__14582 (
            .O(N__66905),
            .I(N__66899));
    Span4Mux_v I__14581 (
            .O(N__66902),
            .I(N__66894));
    LocalMux I__14580 (
            .O(N__66899),
            .I(N__66894));
    Span4Mux_h I__14579 (
            .O(N__66894),
            .I(N__66891));
    Odrv4 I__14578 (
            .O(N__66891),
            .I(side_order_1));
    InMux I__14577 (
            .O(N__66888),
            .I(N__66883));
    InMux I__14576 (
            .O(N__66887),
            .I(N__66878));
    InMux I__14575 (
            .O(N__66886),
            .I(N__66878));
    LocalMux I__14574 (
            .O(N__66883),
            .I(\pid_side.pid_preregZ0Z_2 ));
    LocalMux I__14573 (
            .O(N__66878),
            .I(\pid_side.pid_preregZ0Z_2 ));
    CascadeMux I__14572 (
            .O(N__66873),
            .I(N__66870));
    InMux I__14571 (
            .O(N__66870),
            .I(N__66866));
    InMux I__14570 (
            .O(N__66869),
            .I(N__66863));
    LocalMux I__14569 (
            .O(N__66866),
            .I(N__66860));
    LocalMux I__14568 (
            .O(N__66863),
            .I(N__66857));
    Span4Mux_v I__14567 (
            .O(N__66860),
            .I(N__66852));
    Span4Mux_h I__14566 (
            .O(N__66857),
            .I(N__66852));
    Odrv4 I__14565 (
            .O(N__66852),
            .I(side_order_2));
    InMux I__14564 (
            .O(N__66849),
            .I(N__66839));
    InMux I__14563 (
            .O(N__66848),
            .I(N__66839));
    InMux I__14562 (
            .O(N__66847),
            .I(N__66839));
    CascadeMux I__14561 (
            .O(N__66846),
            .I(N__66835));
    LocalMux I__14560 (
            .O(N__66839),
            .I(N__66832));
    InMux I__14559 (
            .O(N__66838),
            .I(N__66828));
    InMux I__14558 (
            .O(N__66835),
            .I(N__66825));
    Span4Mux_h I__14557 (
            .O(N__66832),
            .I(N__66822));
    InMux I__14556 (
            .O(N__66831),
            .I(N__66819));
    LocalMux I__14555 (
            .O(N__66828),
            .I(\pid_side.N_75 ));
    LocalMux I__14554 (
            .O(N__66825),
            .I(\pid_side.N_75 ));
    Odrv4 I__14553 (
            .O(N__66822),
            .I(\pid_side.N_75 ));
    LocalMux I__14552 (
            .O(N__66819),
            .I(\pid_side.N_75 ));
    CascadeMux I__14551 (
            .O(N__66810),
            .I(N__66806));
    CascadeMux I__14550 (
            .O(N__66809),
            .I(N__66802));
    InMux I__14549 (
            .O(N__66806),
            .I(N__66799));
    InMux I__14548 (
            .O(N__66805),
            .I(N__66794));
    InMux I__14547 (
            .O(N__66802),
            .I(N__66794));
    LocalMux I__14546 (
            .O(N__66799),
            .I(\pid_side.pid_preregZ0Z_3 ));
    LocalMux I__14545 (
            .O(N__66794),
            .I(\pid_side.pid_preregZ0Z_3 ));
    InMux I__14544 (
            .O(N__66789),
            .I(N__66786));
    LocalMux I__14543 (
            .O(N__66786),
            .I(N__66782));
    InMux I__14542 (
            .O(N__66785),
            .I(N__66779));
    Span4Mux_v I__14541 (
            .O(N__66782),
            .I(N__66774));
    LocalMux I__14540 (
            .O(N__66779),
            .I(N__66774));
    Span4Mux_v I__14539 (
            .O(N__66774),
            .I(N__66771));
    Odrv4 I__14538 (
            .O(N__66771),
            .I(side_order_3));
    InMux I__14537 (
            .O(N__66768),
            .I(N__66765));
    LocalMux I__14536 (
            .O(N__66765),
            .I(N__66762));
    Span4Mux_h I__14535 (
            .O(N__66762),
            .I(N__66758));
    CascadeMux I__14534 (
            .O(N__66761),
            .I(N__66755));
    Span4Mux_h I__14533 (
            .O(N__66758),
            .I(N__66752));
    InMux I__14532 (
            .O(N__66755),
            .I(N__66749));
    Odrv4 I__14531 (
            .O(N__66752),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    LocalMux I__14530 (
            .O(N__66749),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    InMux I__14529 (
            .O(N__66744),
            .I(N__66741));
    LocalMux I__14528 (
            .O(N__66741),
            .I(N__66738));
    Span4Mux_v I__14527 (
            .O(N__66738),
            .I(N__66735));
    Span4Mux_h I__14526 (
            .O(N__66735),
            .I(N__66730));
    InMux I__14525 (
            .O(N__66734),
            .I(N__66725));
    InMux I__14524 (
            .O(N__66733),
            .I(N__66725));
    Odrv4 I__14523 (
            .O(N__66730),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__14522 (
            .O(N__66725),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__14521 (
            .O(N__66720),
            .I(N__66717));
    LocalMux I__14520 (
            .O(N__66717),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__14519 (
            .O(N__66714),
            .I(N__66711));
    LocalMux I__14518 (
            .O(N__66711),
            .I(N__66707));
    CascadeMux I__14517 (
            .O(N__66710),
            .I(N__66704));
    Span4Mux_v I__14516 (
            .O(N__66707),
            .I(N__66701));
    InMux I__14515 (
            .O(N__66704),
            .I(N__66698));
    Span4Mux_h I__14514 (
            .O(N__66701),
            .I(N__66693));
    LocalMux I__14513 (
            .O(N__66698),
            .I(N__66693));
    Odrv4 I__14512 (
            .O(N__66693),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    InMux I__14511 (
            .O(N__66690),
            .I(N__66687));
    LocalMux I__14510 (
            .O(N__66687),
            .I(N__66684));
    Span4Mux_h I__14509 (
            .O(N__66684),
            .I(N__66681));
    Span4Mux_h I__14508 (
            .O(N__66681),
            .I(N__66676));
    InMux I__14507 (
            .O(N__66680),
            .I(N__66671));
    InMux I__14506 (
            .O(N__66679),
            .I(N__66671));
    Odrv4 I__14505 (
            .O(N__66676),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    LocalMux I__14504 (
            .O(N__66671),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__14503 (
            .O(N__66666),
            .I(N__66663));
    LocalMux I__14502 (
            .O(N__66663),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__14501 (
            .O(N__66660),
            .I(N__66657));
    LocalMux I__14500 (
            .O(N__66657),
            .I(N__66653));
    CascadeMux I__14499 (
            .O(N__66656),
            .I(N__66650));
    Span4Mux_v I__14498 (
            .O(N__66653),
            .I(N__66647));
    InMux I__14497 (
            .O(N__66650),
            .I(N__66644));
    Span4Mux_h I__14496 (
            .O(N__66647),
            .I(N__66641));
    LocalMux I__14495 (
            .O(N__66644),
            .I(N__66638));
    Odrv4 I__14494 (
            .O(N__66641),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    Odrv4 I__14493 (
            .O(N__66638),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    InMux I__14492 (
            .O(N__66633),
            .I(N__66630));
    LocalMux I__14491 (
            .O(N__66630),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__14490 (
            .O(N__66627),
            .I(N__66624));
    LocalMux I__14489 (
            .O(N__66624),
            .I(N__66621));
    Odrv4 I__14488 (
            .O(N__66621),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    CascadeMux I__14487 (
            .O(N__66618),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0_cascade_ ));
    InMux I__14486 (
            .O(N__66615),
            .I(N__66612));
    LocalMux I__14485 (
            .O(N__66612),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__14484 (
            .O(N__66609),
            .I(N__66606));
    LocalMux I__14483 (
            .O(N__66606),
            .I(N__66601));
    InMux I__14482 (
            .O(N__66605),
            .I(N__66596));
    InMux I__14481 (
            .O(N__66604),
            .I(N__66596));
    Span12Mux_h I__14480 (
            .O(N__66601),
            .I(N__66593));
    LocalMux I__14479 (
            .O(N__66596),
            .I(N__66590));
    Odrv12 I__14478 (
            .O(N__66593),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__14477 (
            .O(N__66590),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__14476 (
            .O(N__66585),
            .I(N__66582));
    LocalMux I__14475 (
            .O(N__66582),
            .I(N__66578));
    CascadeMux I__14474 (
            .O(N__66581),
            .I(N__66575));
    Span4Mux_h I__14473 (
            .O(N__66578),
            .I(N__66572));
    InMux I__14472 (
            .O(N__66575),
            .I(N__66569));
    Odrv4 I__14471 (
            .O(N__66572),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    LocalMux I__14470 (
            .O(N__66569),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    InMux I__14469 (
            .O(N__66564),
            .I(N__66560));
    CascadeMux I__14468 (
            .O(N__66563),
            .I(N__66557));
    LocalMux I__14467 (
            .O(N__66560),
            .I(N__66554));
    InMux I__14466 (
            .O(N__66557),
            .I(N__66548));
    Span4Mux_h I__14465 (
            .O(N__66554),
            .I(N__66545));
    InMux I__14464 (
            .O(N__66553),
            .I(N__66540));
    InMux I__14463 (
            .O(N__66552),
            .I(N__66540));
    InMux I__14462 (
            .O(N__66551),
            .I(N__66537));
    LocalMux I__14461 (
            .O(N__66548),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__14460 (
            .O(N__66545),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__14459 (
            .O(N__66540),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__14458 (
            .O(N__66537),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    InMux I__14457 (
            .O(N__66528),
            .I(N__66525));
    LocalMux I__14456 (
            .O(N__66525),
            .I(N__66520));
    CascadeMux I__14455 (
            .O(N__66524),
            .I(N__66516));
    InMux I__14454 (
            .O(N__66523),
            .I(N__66511));
    Span4Mux_h I__14453 (
            .O(N__66520),
            .I(N__66508));
    InMux I__14452 (
            .O(N__66519),
            .I(N__66505));
    InMux I__14451 (
            .O(N__66516),
            .I(N__66502));
    InMux I__14450 (
            .O(N__66515),
            .I(N__66497));
    InMux I__14449 (
            .O(N__66514),
            .I(N__66497));
    LocalMux I__14448 (
            .O(N__66511),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__14447 (
            .O(N__66508),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__14446 (
            .O(N__66505),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__14445 (
            .O(N__66502),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__14444 (
            .O(N__66497),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    CascadeMux I__14443 (
            .O(N__66486),
            .I(N__66483));
    InMux I__14442 (
            .O(N__66483),
            .I(N__66477));
    InMux I__14441 (
            .O(N__66482),
            .I(N__66474));
    InMux I__14440 (
            .O(N__66481),
            .I(N__66471));
    CascadeMux I__14439 (
            .O(N__66480),
            .I(N__66465));
    LocalMux I__14438 (
            .O(N__66477),
            .I(N__66462));
    LocalMux I__14437 (
            .O(N__66474),
            .I(N__66457));
    LocalMux I__14436 (
            .O(N__66471),
            .I(N__66457));
    InMux I__14435 (
            .O(N__66470),
            .I(N__66454));
    InMux I__14434 (
            .O(N__66469),
            .I(N__66447));
    InMux I__14433 (
            .O(N__66468),
            .I(N__66447));
    InMux I__14432 (
            .O(N__66465),
            .I(N__66447));
    Odrv12 I__14431 (
            .O(N__66462),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__14430 (
            .O(N__66457),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__14429 (
            .O(N__66454),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__14428 (
            .O(N__66447),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__14427 (
            .O(N__66438),
            .I(N__66434));
    InMux I__14426 (
            .O(N__66437),
            .I(N__66429));
    InMux I__14425 (
            .O(N__66434),
            .I(N__66424));
    InMux I__14424 (
            .O(N__66433),
            .I(N__66424));
    CascadeMux I__14423 (
            .O(N__66432),
            .I(N__66421));
    LocalMux I__14422 (
            .O(N__66429),
            .I(N__66415));
    LocalMux I__14421 (
            .O(N__66424),
            .I(N__66412));
    InMux I__14420 (
            .O(N__66421),
            .I(N__66407));
    InMux I__14419 (
            .O(N__66420),
            .I(N__66407));
    InMux I__14418 (
            .O(N__66419),
            .I(N__66402));
    InMux I__14417 (
            .O(N__66418),
            .I(N__66402));
    Span4Mux_v I__14416 (
            .O(N__66415),
            .I(N__66397));
    Span4Mux_v I__14415 (
            .O(N__66412),
            .I(N__66397));
    LocalMux I__14414 (
            .O(N__66407),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__14413 (
            .O(N__66402),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__14412 (
            .O(N__66397),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__14411 (
            .O(N__66390),
            .I(N__66386));
    InMux I__14410 (
            .O(N__66389),
            .I(N__66378));
    InMux I__14409 (
            .O(N__66386),
            .I(N__66378));
    InMux I__14408 (
            .O(N__66385),
            .I(N__66378));
    LocalMux I__14407 (
            .O(N__66378),
            .I(N__66374));
    InMux I__14406 (
            .O(N__66377),
            .I(N__66371));
    Odrv4 I__14405 (
            .O(N__66374),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ));
    LocalMux I__14404 (
            .O(N__66371),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ));
    CascadeMux I__14403 (
            .O(N__66366),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ));
    InMux I__14402 (
            .O(N__66363),
            .I(N__66360));
    LocalMux I__14401 (
            .O(N__66360),
            .I(N__66357));
    Odrv4 I__14400 (
            .O(N__66357),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    InMux I__14399 (
            .O(N__66354),
            .I(N__66351));
    LocalMux I__14398 (
            .O(N__66351),
            .I(N__66348));
    Span4Mux_v I__14397 (
            .O(N__66348),
            .I(N__66343));
    InMux I__14396 (
            .O(N__66347),
            .I(N__66340));
    InMux I__14395 (
            .O(N__66346),
            .I(N__66337));
    Span4Mux_h I__14394 (
            .O(N__66343),
            .I(N__66334));
    LocalMux I__14393 (
            .O(N__66340),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__14392 (
            .O(N__66337),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    Odrv4 I__14391 (
            .O(N__66334),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    CascadeMux I__14390 (
            .O(N__66327),
            .I(N__66323));
    InMux I__14389 (
            .O(N__66326),
            .I(N__66318));
    InMux I__14388 (
            .O(N__66323),
            .I(N__66318));
    LocalMux I__14387 (
            .O(N__66318),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__14386 (
            .O(N__66315),
            .I(N__66312));
    LocalMux I__14385 (
            .O(N__66312),
            .I(N__66309));
    Span4Mux_v I__14384 (
            .O(N__66309),
            .I(N__66304));
    InMux I__14383 (
            .O(N__66308),
            .I(N__66301));
    InMux I__14382 (
            .O(N__66307),
            .I(N__66298));
    Span4Mux_h I__14381 (
            .O(N__66304),
            .I(N__66295));
    LocalMux I__14380 (
            .O(N__66301),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__14379 (
            .O(N__66298),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__14378 (
            .O(N__66295),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__14377 (
            .O(N__66288),
            .I(N__66285));
    LocalMux I__14376 (
            .O(N__66285),
            .I(N__66282));
    Span4Mux_h I__14375 (
            .O(N__66282),
            .I(N__66279));
    Span4Mux_v I__14374 (
            .O(N__66279),
            .I(N__66276));
    Odrv4 I__14373 (
            .O(N__66276),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    CascadeMux I__14372 (
            .O(N__66273),
            .I(N__66270));
    InMux I__14371 (
            .O(N__66270),
            .I(N__66267));
    LocalMux I__14370 (
            .O(N__66267),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__14369 (
            .O(N__66264),
            .I(N__66261));
    LocalMux I__14368 (
            .O(N__66261),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__14367 (
            .O(N__66258),
            .I(N__66255));
    LocalMux I__14366 (
            .O(N__66255),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    CascadeMux I__14365 (
            .O(N__66252),
            .I(N__66248));
    InMux I__14364 (
            .O(N__66251),
            .I(N__66245));
    InMux I__14363 (
            .O(N__66248),
            .I(N__66242));
    LocalMux I__14362 (
            .O(N__66245),
            .I(N__66239));
    LocalMux I__14361 (
            .O(N__66242),
            .I(N__66236));
    Span4Mux_h I__14360 (
            .O(N__66239),
            .I(N__66231));
    Span4Mux_h I__14359 (
            .O(N__66236),
            .I(N__66231));
    Odrv4 I__14358 (
            .O(N__66231),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__14357 (
            .O(N__66228),
            .I(N__66219));
    InMux I__14356 (
            .O(N__66227),
            .I(N__66219));
    InMux I__14355 (
            .O(N__66226),
            .I(N__66219));
    LocalMux I__14354 (
            .O(N__66219),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__14353 (
            .O(N__66216),
            .I(N__66213));
    LocalMux I__14352 (
            .O(N__66213),
            .I(N__66209));
    InMux I__14351 (
            .O(N__66212),
            .I(N__66206));
    Sp12to4 I__14350 (
            .O(N__66209),
            .I(N__66203));
    LocalMux I__14349 (
            .O(N__66206),
            .I(N__66200));
    Span12Mux_s11_v I__14348 (
            .O(N__66203),
            .I(N__66197));
    Span4Mux_h I__14347 (
            .O(N__66200),
            .I(N__66194));
    Odrv12 I__14346 (
            .O(N__66197),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    Odrv4 I__14345 (
            .O(N__66194),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__14344 (
            .O(N__66189),
            .I(N__66186));
    LocalMux I__14343 (
            .O(N__66186),
            .I(N__66183));
    Span4Mux_v I__14342 (
            .O(N__66183),
            .I(N__66180));
    Span4Mux_h I__14341 (
            .O(N__66180),
            .I(N__66177));
    Odrv4 I__14340 (
            .O(N__66177),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__14339 (
            .O(N__66174),
            .I(N__66171));
    LocalMux I__14338 (
            .O(N__66171),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__14337 (
            .O(N__66168),
            .I(N__66164));
    CascadeMux I__14336 (
            .O(N__66167),
            .I(N__66161));
    LocalMux I__14335 (
            .O(N__66164),
            .I(N__66158));
    InMux I__14334 (
            .O(N__66161),
            .I(N__66155));
    Odrv12 I__14333 (
            .O(N__66158),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    LocalMux I__14332 (
            .O(N__66155),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    CascadeMux I__14331 (
            .O(N__66150),
            .I(N__66146));
    InMux I__14330 (
            .O(N__66149),
            .I(N__66143));
    InMux I__14329 (
            .O(N__66146),
            .I(N__66139));
    LocalMux I__14328 (
            .O(N__66143),
            .I(N__66136));
    InMux I__14327 (
            .O(N__66142),
            .I(N__66133));
    LocalMux I__14326 (
            .O(N__66139),
            .I(N__66128));
    Span4Mux_h I__14325 (
            .O(N__66136),
            .I(N__66128));
    LocalMux I__14324 (
            .O(N__66133),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__14323 (
            .O(N__66128),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__14322 (
            .O(N__66123),
            .I(N__66120));
    LocalMux I__14321 (
            .O(N__66120),
            .I(N__66117));
    Span4Mux_h I__14320 (
            .O(N__66117),
            .I(N__66114));
    Odrv4 I__14319 (
            .O(N__66114),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__14318 (
            .O(N__66111),
            .I(N__66108));
    LocalMux I__14317 (
            .O(N__66108),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    CascadeMux I__14316 (
            .O(N__66105),
            .I(\pid_side.N_116_0_0_cascade_ ));
    InMux I__14315 (
            .O(N__66102),
            .I(N__66099));
    LocalMux I__14314 (
            .O(N__66099),
            .I(\pid_side.un4_error_i_reg_31_ns_1_0 ));
    CascadeMux I__14313 (
            .O(N__66096),
            .I(\pid_side.g2_cascade_ ));
    InMux I__14312 (
            .O(N__66093),
            .I(N__66090));
    LocalMux I__14311 (
            .O(N__66090),
            .I(\pid_side.N_117_0 ));
    InMux I__14310 (
            .O(N__66087),
            .I(N__66084));
    LocalMux I__14309 (
            .O(N__66084),
            .I(N__66081));
    Span4Mux_h I__14308 (
            .O(N__66081),
            .I(N__66078));
    Odrv4 I__14307 (
            .O(N__66078),
            .I(\pid_side.g0_i_m4_0_1 ));
    InMux I__14306 (
            .O(N__66075),
            .I(N__66072));
    LocalMux I__14305 (
            .O(N__66072),
            .I(\pid_side.N_10 ));
    InMux I__14304 (
            .O(N__66069),
            .I(N__66056));
    InMux I__14303 (
            .O(N__66068),
            .I(N__66056));
    InMux I__14302 (
            .O(N__66067),
            .I(N__66049));
    InMux I__14301 (
            .O(N__66066),
            .I(N__66049));
    InMux I__14300 (
            .O(N__66065),
            .I(N__66049));
    CascadeMux I__14299 (
            .O(N__66064),
            .I(N__66046));
    CascadeMux I__14298 (
            .O(N__66063),
            .I(N__66035));
    CascadeMux I__14297 (
            .O(N__66062),
            .I(N__66031));
    InMux I__14296 (
            .O(N__66061),
            .I(N__66024));
    LocalMux I__14295 (
            .O(N__66056),
            .I(N__66019));
    LocalMux I__14294 (
            .O(N__66049),
            .I(N__66019));
    InMux I__14293 (
            .O(N__66046),
            .I(N__66016));
    InMux I__14292 (
            .O(N__66045),
            .I(N__66013));
    InMux I__14291 (
            .O(N__66044),
            .I(N__66008));
    InMux I__14290 (
            .O(N__66043),
            .I(N__66008));
    InMux I__14289 (
            .O(N__66042),
            .I(N__66005));
    InMux I__14288 (
            .O(N__66041),
            .I(N__66000));
    InMux I__14287 (
            .O(N__66040),
            .I(N__66000));
    InMux I__14286 (
            .O(N__66039),
            .I(N__65994));
    InMux I__14285 (
            .O(N__66038),
            .I(N__65994));
    InMux I__14284 (
            .O(N__66035),
            .I(N__65991));
    InMux I__14283 (
            .O(N__66034),
            .I(N__65986));
    InMux I__14282 (
            .O(N__66031),
            .I(N__65986));
    InMux I__14281 (
            .O(N__66030),
            .I(N__65982));
    InMux I__14280 (
            .O(N__66029),
            .I(N__65979));
    InMux I__14279 (
            .O(N__66028),
            .I(N__65974));
    InMux I__14278 (
            .O(N__66027),
            .I(N__65974));
    LocalMux I__14277 (
            .O(N__66024),
            .I(N__65971));
    Span4Mux_v I__14276 (
            .O(N__66019),
            .I(N__65966));
    LocalMux I__14275 (
            .O(N__66016),
            .I(N__65966));
    LocalMux I__14274 (
            .O(N__66013),
            .I(N__65963));
    LocalMux I__14273 (
            .O(N__66008),
            .I(N__65960));
    LocalMux I__14272 (
            .O(N__66005),
            .I(N__65957));
    LocalMux I__14271 (
            .O(N__66000),
            .I(N__65954));
    InMux I__14270 (
            .O(N__65999),
            .I(N__65951));
    LocalMux I__14269 (
            .O(N__65994),
            .I(N__65944));
    LocalMux I__14268 (
            .O(N__65991),
            .I(N__65944));
    LocalMux I__14267 (
            .O(N__65986),
            .I(N__65944));
    InMux I__14266 (
            .O(N__65985),
            .I(N__65941));
    LocalMux I__14265 (
            .O(N__65982),
            .I(N__65938));
    LocalMux I__14264 (
            .O(N__65979),
            .I(N__65933));
    LocalMux I__14263 (
            .O(N__65974),
            .I(N__65933));
    Span4Mux_h I__14262 (
            .O(N__65971),
            .I(N__65924));
    Span4Mux_h I__14261 (
            .O(N__65966),
            .I(N__65924));
    Span4Mux_v I__14260 (
            .O(N__65963),
            .I(N__65924));
    Span4Mux_h I__14259 (
            .O(N__65960),
            .I(N__65924));
    Span4Mux_h I__14258 (
            .O(N__65957),
            .I(N__65919));
    Span4Mux_h I__14257 (
            .O(N__65954),
            .I(N__65919));
    LocalMux I__14256 (
            .O(N__65951),
            .I(xy_ki_2_rep1));
    Odrv12 I__14255 (
            .O(N__65944),
            .I(xy_ki_2_rep1));
    LocalMux I__14254 (
            .O(N__65941),
            .I(xy_ki_2_rep1));
    Odrv4 I__14253 (
            .O(N__65938),
            .I(xy_ki_2_rep1));
    Odrv4 I__14252 (
            .O(N__65933),
            .I(xy_ki_2_rep1));
    Odrv4 I__14251 (
            .O(N__65924),
            .I(xy_ki_2_rep1));
    Odrv4 I__14250 (
            .O(N__65919),
            .I(xy_ki_2_rep1));
    InMux I__14249 (
            .O(N__65904),
            .I(N__65901));
    LocalMux I__14248 (
            .O(N__65901),
            .I(\pid_side.N_61_0_0 ));
    CascadeMux I__14247 (
            .O(N__65898),
            .I(\pid_side.N_60_0_0_cascade_ ));
    InMux I__14246 (
            .O(N__65895),
            .I(N__65892));
    LocalMux I__14245 (
            .O(N__65892),
            .I(N__65889));
    Odrv4 I__14244 (
            .O(N__65889),
            .I(\pid_side.un4_error_i_reg_30_ns_1_0 ));
    InMux I__14243 (
            .O(N__65886),
            .I(N__65883));
    LocalMux I__14242 (
            .O(N__65883),
            .I(N__65880));
    Span12Mux_s8_v I__14241 (
            .O(N__65880),
            .I(N__65877));
    Odrv12 I__14240 (
            .O(N__65877),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    CEMux I__14239 (
            .O(N__65874),
            .I(N__65870));
    CEMux I__14238 (
            .O(N__65873),
            .I(N__65867));
    LocalMux I__14237 (
            .O(N__65870),
            .I(N__65862));
    LocalMux I__14236 (
            .O(N__65867),
            .I(N__65859));
    CEMux I__14235 (
            .O(N__65866),
            .I(N__65856));
    CEMux I__14234 (
            .O(N__65865),
            .I(N__65852));
    Span4Mux_v I__14233 (
            .O(N__65862),
            .I(N__65847));
    Span4Mux_v I__14232 (
            .O(N__65859),
            .I(N__65847));
    LocalMux I__14231 (
            .O(N__65856),
            .I(N__65844));
    CEMux I__14230 (
            .O(N__65855),
            .I(N__65841));
    LocalMux I__14229 (
            .O(N__65852),
            .I(N__65838));
    Span4Mux_h I__14228 (
            .O(N__65847),
            .I(N__65835));
    Span4Mux_h I__14227 (
            .O(N__65844),
            .I(N__65832));
    LocalMux I__14226 (
            .O(N__65841),
            .I(N__65827));
    Span4Mux_h I__14225 (
            .O(N__65838),
            .I(N__65827));
    Odrv4 I__14224 (
            .O(N__65835),
            .I(\ppm_encoder_1.N_2569_0 ));
    Odrv4 I__14223 (
            .O(N__65832),
            .I(\ppm_encoder_1.N_2569_0 ));
    Odrv4 I__14222 (
            .O(N__65827),
            .I(\ppm_encoder_1.N_2569_0 ));
    CascadeMux I__14221 (
            .O(N__65820),
            .I(\pid_side.m21_1_cascade_ ));
    InMux I__14220 (
            .O(N__65817),
            .I(N__65814));
    LocalMux I__14219 (
            .O(N__65814),
            .I(N__65809));
    InMux I__14218 (
            .O(N__65813),
            .I(N__65804));
    InMux I__14217 (
            .O(N__65812),
            .I(N__65804));
    Odrv4 I__14216 (
            .O(N__65809),
            .I(\pid_side.N_22_0 ));
    LocalMux I__14215 (
            .O(N__65804),
            .I(\pid_side.N_22_0 ));
    InMux I__14214 (
            .O(N__65799),
            .I(N__65796));
    LocalMux I__14213 (
            .O(N__65796),
            .I(\pid_side.m30_1_ns_1 ));
    InMux I__14212 (
            .O(N__65793),
            .I(N__65790));
    LocalMux I__14211 (
            .O(N__65790),
            .I(\pid_side.error_cry_4_c_RNINOGZ0Z52 ));
    InMux I__14210 (
            .O(N__65787),
            .I(N__65784));
    LocalMux I__14209 (
            .O(N__65784),
            .I(\pid_side.N_30_1 ));
    InMux I__14208 (
            .O(N__65781),
            .I(N__65773));
    InMux I__14207 (
            .O(N__65780),
            .I(N__65773));
    InMux I__14206 (
            .O(N__65779),
            .I(N__65770));
    InMux I__14205 (
            .O(N__65778),
            .I(N__65767));
    LocalMux I__14204 (
            .O(N__65773),
            .I(N__65764));
    LocalMux I__14203 (
            .O(N__65770),
            .I(N__65759));
    LocalMux I__14202 (
            .O(N__65767),
            .I(N__65759));
    Odrv4 I__14201 (
            .O(N__65764),
            .I(\pid_side.m1_0_03 ));
    Odrv4 I__14200 (
            .O(N__65759),
            .I(\pid_side.m1_0_03 ));
    CascadeMux I__14199 (
            .O(N__65754),
            .I(\pid_side.m1_0_03_cascade_ ));
    InMux I__14198 (
            .O(N__65751),
            .I(N__65748));
    LocalMux I__14197 (
            .O(N__65748),
            .I(N__65730));
    InMux I__14196 (
            .O(N__65747),
            .I(N__65727));
    InMux I__14195 (
            .O(N__65746),
            .I(N__65724));
    InMux I__14194 (
            .O(N__65745),
            .I(N__65719));
    InMux I__14193 (
            .O(N__65744),
            .I(N__65719));
    InMux I__14192 (
            .O(N__65743),
            .I(N__65716));
    InMux I__14191 (
            .O(N__65742),
            .I(N__65707));
    InMux I__14190 (
            .O(N__65741),
            .I(N__65707));
    InMux I__14189 (
            .O(N__65740),
            .I(N__65707));
    InMux I__14188 (
            .O(N__65739),
            .I(N__65707));
    InMux I__14187 (
            .O(N__65738),
            .I(N__65702));
    InMux I__14186 (
            .O(N__65737),
            .I(N__65702));
    InMux I__14185 (
            .O(N__65736),
            .I(N__65699));
    InMux I__14184 (
            .O(N__65735),
            .I(N__65689));
    InMux I__14183 (
            .O(N__65734),
            .I(N__65689));
    InMux I__14182 (
            .O(N__65733),
            .I(N__65689));
    Span4Mux_h I__14181 (
            .O(N__65730),
            .I(N__65686));
    LocalMux I__14180 (
            .O(N__65727),
            .I(N__65683));
    LocalMux I__14179 (
            .O(N__65724),
            .I(N__65673));
    LocalMux I__14178 (
            .O(N__65719),
            .I(N__65673));
    LocalMux I__14177 (
            .O(N__65716),
            .I(N__65670));
    LocalMux I__14176 (
            .O(N__65707),
            .I(N__65665));
    LocalMux I__14175 (
            .O(N__65702),
            .I(N__65665));
    LocalMux I__14174 (
            .O(N__65699),
            .I(N__65662));
    CascadeMux I__14173 (
            .O(N__65698),
            .I(N__65659));
    CascadeMux I__14172 (
            .O(N__65697),
            .I(N__65656));
    InMux I__14171 (
            .O(N__65696),
            .I(N__65653));
    LocalMux I__14170 (
            .O(N__65689),
            .I(N__65650));
    Span4Mux_h I__14169 (
            .O(N__65686),
            .I(N__65645));
    Span4Mux_h I__14168 (
            .O(N__65683),
            .I(N__65645));
    InMux I__14167 (
            .O(N__65682),
            .I(N__65638));
    InMux I__14166 (
            .O(N__65681),
            .I(N__65638));
    InMux I__14165 (
            .O(N__65680),
            .I(N__65638));
    InMux I__14164 (
            .O(N__65679),
            .I(N__65633));
    InMux I__14163 (
            .O(N__65678),
            .I(N__65633));
    Span4Mux_h I__14162 (
            .O(N__65673),
            .I(N__65630));
    Span4Mux_h I__14161 (
            .O(N__65670),
            .I(N__65623));
    Span4Mux_v I__14160 (
            .O(N__65665),
            .I(N__65623));
    Span4Mux_h I__14159 (
            .O(N__65662),
            .I(N__65623));
    InMux I__14158 (
            .O(N__65659),
            .I(N__65618));
    InMux I__14157 (
            .O(N__65656),
            .I(N__65618));
    LocalMux I__14156 (
            .O(N__65653),
            .I(xy_ki_2_rep2));
    Odrv12 I__14155 (
            .O(N__65650),
            .I(xy_ki_2_rep2));
    Odrv4 I__14154 (
            .O(N__65645),
            .I(xy_ki_2_rep2));
    LocalMux I__14153 (
            .O(N__65638),
            .I(xy_ki_2_rep2));
    LocalMux I__14152 (
            .O(N__65633),
            .I(xy_ki_2_rep2));
    Odrv4 I__14151 (
            .O(N__65630),
            .I(xy_ki_2_rep2));
    Odrv4 I__14150 (
            .O(N__65623),
            .I(xy_ki_2_rep2));
    LocalMux I__14149 (
            .O(N__65618),
            .I(xy_ki_2_rep2));
    InMux I__14148 (
            .O(N__65601),
            .I(N__65598));
    LocalMux I__14147 (
            .O(N__65598),
            .I(N__65595));
    Span4Mux_h I__14146 (
            .O(N__65595),
            .I(N__65592));
    Odrv4 I__14145 (
            .O(N__65592),
            .I(\pid_side.m1_2_03 ));
    InMux I__14144 (
            .O(N__65589),
            .I(N__65586));
    LocalMux I__14143 (
            .O(N__65586),
            .I(\pid_side.N_126_0 ));
    InMux I__14142 (
            .O(N__65583),
            .I(N__65580));
    LocalMux I__14141 (
            .O(N__65580),
            .I(N__65577));
    Odrv4 I__14140 (
            .O(N__65577),
            .I(\pid_side.g3_0 ));
    CascadeMux I__14139 (
            .O(N__65574),
            .I(\pid_side.g1_0_cascade_ ));
    InMux I__14138 (
            .O(N__65571),
            .I(N__65568));
    LocalMux I__14137 (
            .O(N__65568),
            .I(N__65565));
    Span4Mux_v I__14136 (
            .O(N__65565),
            .I(N__65562));
    Span4Mux_v I__14135 (
            .O(N__65562),
            .I(N__65559));
    Odrv4 I__14134 (
            .O(N__65559),
            .I(\pid_side.error_i_regZ0Z_21 ));
    InMux I__14133 (
            .O(N__65556),
            .I(N__65553));
    LocalMux I__14132 (
            .O(N__65553),
            .I(\pid_side.N_89_0_0 ));
    CascadeMux I__14131 (
            .O(N__65550),
            .I(\pid_side.g0_9_1_cascade_ ));
    CascadeMux I__14130 (
            .O(N__65547),
            .I(\pid_side.N_22_0_0_cascade_ ));
    InMux I__14129 (
            .O(N__65544),
            .I(N__65541));
    LocalMux I__14128 (
            .O(N__65541),
            .I(\pid_side.N_57_0_0 ));
    CascadeMux I__14127 (
            .O(N__65538),
            .I(\pid_side.g1_cascade_ ));
    CascadeMux I__14126 (
            .O(N__65535),
            .I(N__65532));
    InMux I__14125 (
            .O(N__65532),
            .I(N__65529));
    LocalMux I__14124 (
            .O(N__65529),
            .I(N__65526));
    Span4Mux_h I__14123 (
            .O(N__65526),
            .I(N__65523));
    Span4Mux_v I__14122 (
            .O(N__65523),
            .I(N__65520));
    Odrv4 I__14121 (
            .O(N__65520),
            .I(\pid_side.error_i_regZ0Z_20 ));
    InMux I__14120 (
            .O(N__65517),
            .I(N__65514));
    LocalMux I__14119 (
            .O(N__65514),
            .I(\pid_side.g3 ));
    CascadeMux I__14118 (
            .O(N__65511),
            .I(\pid_side.m88_0_ns_1_0_cascade_ ));
    InMux I__14117 (
            .O(N__65508),
            .I(N__65505));
    LocalMux I__14116 (
            .O(N__65505),
            .I(N__65502));
    Odrv4 I__14115 (
            .O(N__65502),
            .I(\pid_side.m48_ns_1 ));
    CascadeMux I__14114 (
            .O(N__65499),
            .I(\pid_side.N_126_cascade_ ));
    CascadeMux I__14113 (
            .O(N__65496),
            .I(\pid_side.m131_0_ns_1_cascade_ ));
    InMux I__14112 (
            .O(N__65493),
            .I(N__65490));
    LocalMux I__14111 (
            .O(N__65490),
            .I(N__65487));
    Span4Mux_h I__14110 (
            .O(N__65487),
            .I(N__65484));
    Odrv4 I__14109 (
            .O(N__65484),
            .I(\pid_side.m21_2_03_0 ));
    InMux I__14108 (
            .O(N__65481),
            .I(N__65475));
    InMux I__14107 (
            .O(N__65480),
            .I(N__65475));
    LocalMux I__14106 (
            .O(N__65475),
            .I(\pid_side.N_89_0 ));
    InMux I__14105 (
            .O(N__65472),
            .I(N__65469));
    LocalMux I__14104 (
            .O(N__65469),
            .I(\pid_side.m93_0_ns_1 ));
    InMux I__14103 (
            .O(N__65466),
            .I(N__65463));
    LocalMux I__14102 (
            .O(N__65463),
            .I(\pid_side.m13_2_03_4_i_0 ));
    CascadeMux I__14101 (
            .O(N__65460),
            .I(N__65453));
    InMux I__14100 (
            .O(N__65459),
            .I(N__65445));
    InMux I__14099 (
            .O(N__65458),
            .I(N__65442));
    CascadeMux I__14098 (
            .O(N__65457),
            .I(N__65438));
    InMux I__14097 (
            .O(N__65456),
            .I(N__65431));
    InMux I__14096 (
            .O(N__65453),
            .I(N__65431));
    InMux I__14095 (
            .O(N__65452),
            .I(N__65431));
    CascadeMux I__14094 (
            .O(N__65451),
            .I(N__65426));
    CascadeMux I__14093 (
            .O(N__65450),
            .I(N__65423));
    InMux I__14092 (
            .O(N__65449),
            .I(N__65420));
    InMux I__14091 (
            .O(N__65448),
            .I(N__65417));
    LocalMux I__14090 (
            .O(N__65445),
            .I(N__65414));
    LocalMux I__14089 (
            .O(N__65442),
            .I(N__65411));
    InMux I__14088 (
            .O(N__65441),
            .I(N__65408));
    InMux I__14087 (
            .O(N__65438),
            .I(N__65403));
    LocalMux I__14086 (
            .O(N__65431),
            .I(N__65400));
    InMux I__14085 (
            .O(N__65430),
            .I(N__65395));
    InMux I__14084 (
            .O(N__65429),
            .I(N__65395));
    InMux I__14083 (
            .O(N__65426),
            .I(N__65390));
    InMux I__14082 (
            .O(N__65423),
            .I(N__65390));
    LocalMux I__14081 (
            .O(N__65420),
            .I(N__65385));
    LocalMux I__14080 (
            .O(N__65417),
            .I(N__65385));
    Span4Mux_h I__14079 (
            .O(N__65414),
            .I(N__65381));
    Span4Mux_v I__14078 (
            .O(N__65411),
            .I(N__65376));
    LocalMux I__14077 (
            .O(N__65408),
            .I(N__65376));
    InMux I__14076 (
            .O(N__65407),
            .I(N__65371));
    InMux I__14075 (
            .O(N__65406),
            .I(N__65371));
    LocalMux I__14074 (
            .O(N__65403),
            .I(N__65360));
    Span4Mux_v I__14073 (
            .O(N__65400),
            .I(N__65360));
    LocalMux I__14072 (
            .O(N__65395),
            .I(N__65360));
    LocalMux I__14071 (
            .O(N__65390),
            .I(N__65360));
    Span4Mux_h I__14070 (
            .O(N__65385),
            .I(N__65360));
    InMux I__14069 (
            .O(N__65384),
            .I(N__65357));
    Span4Mux_v I__14068 (
            .O(N__65381),
            .I(N__65350));
    Span4Mux_h I__14067 (
            .O(N__65376),
            .I(N__65350));
    LocalMux I__14066 (
            .O(N__65371),
            .I(N__65350));
    Span4Mux_v I__14065 (
            .O(N__65360),
            .I(N__65345));
    LocalMux I__14064 (
            .O(N__65357),
            .I(N__65345));
    Span4Mux_v I__14063 (
            .O(N__65350),
            .I(N__65342));
    Span4Mux_h I__14062 (
            .O(N__65345),
            .I(N__65339));
    Span4Mux_v I__14061 (
            .O(N__65342),
            .I(N__65336));
    Span4Mux_v I__14060 (
            .O(N__65339),
            .I(N__65333));
    Odrv4 I__14059 (
            .O(N__65336),
            .I(pid_side_N_166));
    Odrv4 I__14058 (
            .O(N__65333),
            .I(pid_side_N_166));
    CascadeMux I__14057 (
            .O(N__65328),
            .I(\pid_side.m13_2_03_4_i_0_cascade_ ));
    CascadeMux I__14056 (
            .O(N__65325),
            .I(N__65322));
    InMux I__14055 (
            .O(N__65322),
            .I(N__65319));
    LocalMux I__14054 (
            .O(N__65319),
            .I(N__65315));
    InMux I__14053 (
            .O(N__65318),
            .I(N__65312));
    Span4Mux_h I__14052 (
            .O(N__65315),
            .I(N__65309));
    LocalMux I__14051 (
            .O(N__65312),
            .I(\pid_side.error_i_regZ0Z_9 ));
    Odrv4 I__14050 (
            .O(N__65309),
            .I(\pid_side.error_i_regZ0Z_9 ));
    InMux I__14049 (
            .O(N__65304),
            .I(N__65298));
    InMux I__14048 (
            .O(N__65303),
            .I(N__65298));
    LocalMux I__14047 (
            .O(N__65298),
            .I(\pid_side.N_88_0 ));
    CascadeMux I__14046 (
            .O(N__65295),
            .I(\pid_side.N_88_0_cascade_ ));
    InMux I__14045 (
            .O(N__65292),
            .I(N__65288));
    InMux I__14044 (
            .O(N__65291),
            .I(N__65285));
    LocalMux I__14043 (
            .O(N__65288),
            .I(\pid_side.N_126 ));
    LocalMux I__14042 (
            .O(N__65285),
            .I(\pid_side.N_126 ));
    InMux I__14041 (
            .O(N__65280),
            .I(N__65277));
    LocalMux I__14040 (
            .O(N__65277),
            .I(N__65274));
    Odrv4 I__14039 (
            .O(N__65274),
            .I(\pid_side.N_127 ));
    InMux I__14038 (
            .O(N__65271),
            .I(N__65268));
    LocalMux I__14037 (
            .O(N__65268),
            .I(N__65265));
    Odrv4 I__14036 (
            .O(N__65265),
            .I(\pid_side.error_cry_4_c_RNINOG52Z0Z_1 ));
    CascadeMux I__14035 (
            .O(N__65262),
            .I(\pid_side.N_36_0_0_cascade_ ));
    InMux I__14034 (
            .O(N__65259),
            .I(N__65250));
    InMux I__14033 (
            .O(N__65258),
            .I(N__65250));
    InMux I__14032 (
            .O(N__65257),
            .I(N__65250));
    LocalMux I__14031 (
            .O(N__65250),
            .I(drone_H_disp_side_11));
    CascadeMux I__14030 (
            .O(N__65247),
            .I(N__65244));
    InMux I__14029 (
            .O(N__65244),
            .I(N__65238));
    InMux I__14028 (
            .O(N__65243),
            .I(N__65238));
    LocalMux I__14027 (
            .O(N__65238),
            .I(side_command_7));
    InMux I__14026 (
            .O(N__65235),
            .I(N__65232));
    LocalMux I__14025 (
            .O(N__65232),
            .I(N__65228));
    InMux I__14024 (
            .O(N__65231),
            .I(N__65225));
    Span4Mux_h I__14023 (
            .O(N__65228),
            .I(N__65222));
    LocalMux I__14022 (
            .O(N__65225),
            .I(N__65218));
    Span4Mux_v I__14021 (
            .O(N__65222),
            .I(N__65215));
    InMux I__14020 (
            .O(N__65221),
            .I(N__65212));
    Span4Mux_h I__14019 (
            .O(N__65218),
            .I(N__65202));
    Span4Mux_h I__14018 (
            .O(N__65215),
            .I(N__65202));
    LocalMux I__14017 (
            .O(N__65212),
            .I(N__65202));
    InMux I__14016 (
            .O(N__65211),
            .I(N__65197));
    InMux I__14015 (
            .O(N__65210),
            .I(N__65194));
    InMux I__14014 (
            .O(N__65209),
            .I(N__65191));
    Span4Mux_v I__14013 (
            .O(N__65202),
            .I(N__65188));
    InMux I__14012 (
            .O(N__65201),
            .I(N__65183));
    InMux I__14011 (
            .O(N__65200),
            .I(N__65183));
    LocalMux I__14010 (
            .O(N__65197),
            .I(N__65180));
    LocalMux I__14009 (
            .O(N__65194),
            .I(N__65175));
    LocalMux I__14008 (
            .O(N__65191),
            .I(N__65175));
    Span4Mux_h I__14007 (
            .O(N__65188),
            .I(N__65172));
    LocalMux I__14006 (
            .O(N__65183),
            .I(N__65169));
    Span4Mux_v I__14005 (
            .O(N__65180),
            .I(N__65166));
    Span12Mux_v I__14004 (
            .O(N__65175),
            .I(N__65163));
    Span4Mux_h I__14003 (
            .O(N__65172),
            .I(N__65160));
    Span4Mux_h I__14002 (
            .O(N__65169),
            .I(N__65157));
    Odrv4 I__14001 (
            .O(N__65166),
            .I(uart_drone_data_4));
    Odrv12 I__14000 (
            .O(N__65163),
            .I(uart_drone_data_4));
    Odrv4 I__13999 (
            .O(N__65160),
            .I(uart_drone_data_4));
    Odrv4 I__13998 (
            .O(N__65157),
            .I(uart_drone_data_4));
    CascadeMux I__13997 (
            .O(N__65148),
            .I(N__65143));
    InMux I__13996 (
            .O(N__65147),
            .I(N__65139));
    InMux I__13995 (
            .O(N__65146),
            .I(N__65132));
    InMux I__13994 (
            .O(N__65143),
            .I(N__65132));
    InMux I__13993 (
            .O(N__65142),
            .I(N__65132));
    LocalMux I__13992 (
            .O(N__65139),
            .I(N__65127));
    LocalMux I__13991 (
            .O(N__65132),
            .I(N__65127));
    Span4Mux_h I__13990 (
            .O(N__65127),
            .I(N__65121));
    CascadeMux I__13989 (
            .O(N__65126),
            .I(N__65118));
    InMux I__13988 (
            .O(N__65125),
            .I(N__65115));
    InMux I__13987 (
            .O(N__65124),
            .I(N__65112));
    Span4Mux_v I__13986 (
            .O(N__65121),
            .I(N__65109));
    InMux I__13985 (
            .O(N__65118),
            .I(N__65106));
    LocalMux I__13984 (
            .O(N__65115),
            .I(N__65101));
    LocalMux I__13983 (
            .O(N__65112),
            .I(N__65101));
    Span4Mux_v I__13982 (
            .O(N__65109),
            .I(N__65096));
    LocalMux I__13981 (
            .O(N__65106),
            .I(N__65096));
    Span12Mux_h I__13980 (
            .O(N__65101),
            .I(N__65093));
    Span4Mux_h I__13979 (
            .O(N__65096),
            .I(N__65090));
    Odrv12 I__13978 (
            .O(N__65093),
            .I(uart_drone_data_7));
    Odrv4 I__13977 (
            .O(N__65090),
            .I(uart_drone_data_7));
    InMux I__13976 (
            .O(N__65085),
            .I(N__65079));
    InMux I__13975 (
            .O(N__65084),
            .I(N__65079));
    LocalMux I__13974 (
            .O(N__65079),
            .I(\dron_frame_decoder_1.drone_H_disp_side_7 ));
    InMux I__13973 (
            .O(N__65076),
            .I(N__65070));
    InMux I__13972 (
            .O(N__65075),
            .I(N__65070));
    LocalMux I__13971 (
            .O(N__65070),
            .I(N__65067));
    Span4Mux_v I__13970 (
            .O(N__65067),
            .I(N__65062));
    InMux I__13969 (
            .O(N__65066),
            .I(N__65059));
    InMux I__13968 (
            .O(N__65065),
            .I(N__65056));
    Odrv4 I__13967 (
            .O(N__65062),
            .I(\pid_side.N_12_1 ));
    LocalMux I__13966 (
            .O(N__65059),
            .I(\pid_side.N_12_1 ));
    LocalMux I__13965 (
            .O(N__65056),
            .I(\pid_side.N_12_1 ));
    InMux I__13964 (
            .O(N__65049),
            .I(N__65043));
    InMux I__13963 (
            .O(N__65048),
            .I(N__65043));
    LocalMux I__13962 (
            .O(N__65043),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    InMux I__13961 (
            .O(N__65040),
            .I(N__65036));
    InMux I__13960 (
            .O(N__65039),
            .I(N__65033));
    LocalMux I__13959 (
            .O(N__65036),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ));
    LocalMux I__13958 (
            .O(N__65033),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ));
    CEMux I__13957 (
            .O(N__65028),
            .I(N__65024));
    CEMux I__13956 (
            .O(N__65027),
            .I(N__65021));
    LocalMux I__13955 (
            .O(N__65024),
            .I(N__65018));
    LocalMux I__13954 (
            .O(N__65021),
            .I(N__65015));
    Span4Mux_h I__13953 (
            .O(N__65018),
            .I(N__65012));
    Span4Mux_h I__13952 (
            .O(N__65015),
            .I(N__65009));
    Span4Mux_v I__13951 (
            .O(N__65012),
            .I(N__65006));
    Span4Mux_v I__13950 (
            .O(N__65009),
            .I(N__65003));
    Odrv4 I__13949 (
            .O(N__65006),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    Odrv4 I__13948 (
            .O(N__65003),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__13947 (
            .O(N__64998),
            .I(N__64989));
    InMux I__13946 (
            .O(N__64997),
            .I(N__64989));
    InMux I__13945 (
            .O(N__64996),
            .I(N__64986));
    InMux I__13944 (
            .O(N__64995),
            .I(N__64980));
    InMux I__13943 (
            .O(N__64994),
            .I(N__64980));
    LocalMux I__13942 (
            .O(N__64989),
            .I(N__64977));
    LocalMux I__13941 (
            .O(N__64986),
            .I(N__64974));
    InMux I__13940 (
            .O(N__64985),
            .I(N__64971));
    LocalMux I__13939 (
            .O(N__64980),
            .I(N__64968));
    Span4Mux_v I__13938 (
            .O(N__64977),
            .I(N__64963));
    Span4Mux_v I__13937 (
            .O(N__64974),
            .I(N__64960));
    LocalMux I__13936 (
            .O(N__64971),
            .I(N__64957));
    Span4Mux_v I__13935 (
            .O(N__64968),
            .I(N__64954));
    InMux I__13934 (
            .O(N__64967),
            .I(N__64951));
    InMux I__13933 (
            .O(N__64966),
            .I(N__64948));
    Span4Mux_h I__13932 (
            .O(N__64963),
            .I(N__64945));
    Span4Mux_h I__13931 (
            .O(N__64960),
            .I(N__64942));
    Span4Mux_h I__13930 (
            .O(N__64957),
            .I(N__64933));
    Span4Mux_v I__13929 (
            .O(N__64954),
            .I(N__64933));
    LocalMux I__13928 (
            .O(N__64951),
            .I(N__64933));
    LocalMux I__13927 (
            .O(N__64948),
            .I(N__64933));
    Span4Mux_h I__13926 (
            .O(N__64945),
            .I(N__64930));
    Span4Mux_v I__13925 (
            .O(N__64942),
            .I(N__64925));
    Span4Mux_v I__13924 (
            .O(N__64933),
            .I(N__64925));
    Odrv4 I__13923 (
            .O(N__64930),
            .I(uart_drone_data_3));
    Odrv4 I__13922 (
            .O(N__64925),
            .I(uart_drone_data_3));
    InMux I__13921 (
            .O(N__64920),
            .I(N__64917));
    LocalMux I__13920 (
            .O(N__64917),
            .I(N__64914));
    Odrv4 I__13919 (
            .O(N__64914),
            .I(\pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ));
    CascadeMux I__13918 (
            .O(N__64911),
            .I(N__64908));
    InMux I__13917 (
            .O(N__64908),
            .I(N__64905));
    LocalMux I__13916 (
            .O(N__64905),
            .I(N__64902));
    Span4Mux_h I__13915 (
            .O(N__64902),
            .I(N__64899));
    Odrv4 I__13914 (
            .O(N__64899),
            .I(\pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ));
    InMux I__13913 (
            .O(N__64896),
            .I(N__64893));
    LocalMux I__13912 (
            .O(N__64893),
            .I(N__64890));
    Span4Mux_h I__13911 (
            .O(N__64890),
            .I(N__64887));
    Odrv4 I__13910 (
            .O(N__64887),
            .I(\pid_side.pid_preregZ0Z_29 ));
    InMux I__13909 (
            .O(N__64884),
            .I(\pid_side.un1_pid_prereg_0_cry_28 ));
    InMux I__13908 (
            .O(N__64881),
            .I(N__64878));
    LocalMux I__13907 (
            .O(N__64878),
            .I(N__64875));
    Odrv4 I__13906 (
            .O(N__64875),
            .I(\pid_side.un1_pid_prereg_0_axb_30 ));
    InMux I__13905 (
            .O(N__64872),
            .I(\pid_side.un1_pid_prereg_0_cry_29 ));
    InMux I__13904 (
            .O(N__64869),
            .I(N__64866));
    LocalMux I__13903 (
            .O(N__64866),
            .I(N__64862));
    InMux I__13902 (
            .O(N__64865),
            .I(N__64858));
    Span4Mux_h I__13901 (
            .O(N__64862),
            .I(N__64855));
    InMux I__13900 (
            .O(N__64861),
            .I(N__64852));
    LocalMux I__13899 (
            .O(N__64858),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    Odrv4 I__13898 (
            .O(N__64855),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    LocalMux I__13897 (
            .O(N__64852),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    CascadeMux I__13896 (
            .O(N__64845),
            .I(\pid_side.un1_pid_prereg_0_21_cascade_ ));
    CascadeMux I__13895 (
            .O(N__64842),
            .I(N__64839));
    InMux I__13894 (
            .O(N__64839),
            .I(N__64836));
    LocalMux I__13893 (
            .O(N__64836),
            .I(\pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ));
    InMux I__13892 (
            .O(N__64833),
            .I(N__64829));
    InMux I__13891 (
            .O(N__64832),
            .I(N__64825));
    LocalMux I__13890 (
            .O(N__64829),
            .I(N__64822));
    InMux I__13889 (
            .O(N__64828),
            .I(N__64819));
    LocalMux I__13888 (
            .O(N__64825),
            .I(N__64814));
    Span4Mux_v I__13887 (
            .O(N__64822),
            .I(N__64814));
    LocalMux I__13886 (
            .O(N__64819),
            .I(N__64811));
    Odrv4 I__13885 (
            .O(N__64814),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    Odrv4 I__13884 (
            .O(N__64811),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    InMux I__13883 (
            .O(N__64806),
            .I(N__64803));
    LocalMux I__13882 (
            .O(N__64803),
            .I(N__64799));
    InMux I__13881 (
            .O(N__64802),
            .I(N__64796));
    Odrv4 I__13880 (
            .O(N__64799),
            .I(\pid_side.un1_pid_prereg_0_20 ));
    LocalMux I__13879 (
            .O(N__64796),
            .I(\pid_side.un1_pid_prereg_0_20 ));
    InMux I__13878 (
            .O(N__64791),
            .I(N__64787));
    InMux I__13877 (
            .O(N__64790),
            .I(N__64784));
    LocalMux I__13876 (
            .O(N__64787),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    LocalMux I__13875 (
            .O(N__64784),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    InMux I__13874 (
            .O(N__64779),
            .I(N__64775));
    InMux I__13873 (
            .O(N__64778),
            .I(N__64772));
    LocalMux I__13872 (
            .O(N__64775),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    LocalMux I__13871 (
            .O(N__64772),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    CascadeMux I__13870 (
            .O(N__64767),
            .I(\pid_side.un1_pid_prereg_0_20_cascade_ ));
    CascadeMux I__13869 (
            .O(N__64764),
            .I(N__64761));
    InMux I__13868 (
            .O(N__64761),
            .I(N__64758));
    LocalMux I__13867 (
            .O(N__64758),
            .I(N__64755));
    Span4Mux_v I__13866 (
            .O(N__64755),
            .I(N__64751));
    InMux I__13865 (
            .O(N__64754),
            .I(N__64748));
    Odrv4 I__13864 (
            .O(N__64751),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    LocalMux I__13863 (
            .O(N__64748),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    InMux I__13862 (
            .O(N__64743),
            .I(N__64740));
    LocalMux I__13861 (
            .O(N__64740),
            .I(\pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ));
    CascadeMux I__13860 (
            .O(N__64737),
            .I(N__64723));
    CascadeMux I__13859 (
            .O(N__64736),
            .I(N__64719));
    CascadeMux I__13858 (
            .O(N__64735),
            .I(N__64716));
    CascadeMux I__13857 (
            .O(N__64734),
            .I(N__64713));
    CascadeMux I__13856 (
            .O(N__64733),
            .I(N__64710));
    CascadeMux I__13855 (
            .O(N__64732),
            .I(N__64707));
    CascadeMux I__13854 (
            .O(N__64731),
            .I(N__64704));
    CascadeMux I__13853 (
            .O(N__64730),
            .I(N__64701));
    InMux I__13852 (
            .O(N__64729),
            .I(N__64698));
    InMux I__13851 (
            .O(N__64728),
            .I(N__64687));
    InMux I__13850 (
            .O(N__64727),
            .I(N__64687));
    InMux I__13849 (
            .O(N__64726),
            .I(N__64687));
    InMux I__13848 (
            .O(N__64723),
            .I(N__64687));
    InMux I__13847 (
            .O(N__64722),
            .I(N__64687));
    InMux I__13846 (
            .O(N__64719),
            .I(N__64682));
    InMux I__13845 (
            .O(N__64716),
            .I(N__64682));
    InMux I__13844 (
            .O(N__64713),
            .I(N__64679));
    InMux I__13843 (
            .O(N__64710),
            .I(N__64676));
    InMux I__13842 (
            .O(N__64707),
            .I(N__64673));
    InMux I__13841 (
            .O(N__64704),
            .I(N__64668));
    InMux I__13840 (
            .O(N__64701),
            .I(N__64668));
    LocalMux I__13839 (
            .O(N__64698),
            .I(N__64663));
    LocalMux I__13838 (
            .O(N__64687),
            .I(N__64663));
    LocalMux I__13837 (
            .O(N__64682),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    LocalMux I__13836 (
            .O(N__64679),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    LocalMux I__13835 (
            .O(N__64676),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    LocalMux I__13834 (
            .O(N__64673),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    LocalMux I__13833 (
            .O(N__64668),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__13832 (
            .O(N__64663),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    InMux I__13831 (
            .O(N__64650),
            .I(N__64644));
    InMux I__13830 (
            .O(N__64649),
            .I(N__64644));
    LocalMux I__13829 (
            .O(N__64644),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ));
    InMux I__13828 (
            .O(N__64641),
            .I(N__64638));
    LocalMux I__13827 (
            .O(N__64638),
            .I(N__64635));
    Span4Mux_h I__13826 (
            .O(N__64635),
            .I(N__64632));
    Odrv4 I__13825 (
            .O(N__64632),
            .I(\pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ));
    InMux I__13824 (
            .O(N__64629),
            .I(N__64626));
    LocalMux I__13823 (
            .O(N__64626),
            .I(N__64623));
    Span4Mux_h I__13822 (
            .O(N__64623),
            .I(N__64620));
    Odrv4 I__13821 (
            .O(N__64620),
            .I(\pid_side.pid_preregZ0Z_21 ));
    InMux I__13820 (
            .O(N__64617),
            .I(\pid_side.un1_pid_prereg_0_cry_20 ));
    InMux I__13819 (
            .O(N__64614),
            .I(N__64611));
    LocalMux I__13818 (
            .O(N__64611),
            .I(N__64608));
    Odrv4 I__13817 (
            .O(N__64608),
            .I(\pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ));
    CascadeMux I__13816 (
            .O(N__64605),
            .I(N__64602));
    InMux I__13815 (
            .O(N__64602),
            .I(N__64599));
    LocalMux I__13814 (
            .O(N__64599),
            .I(N__64596));
    Odrv4 I__13813 (
            .O(N__64596),
            .I(\pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ));
    InMux I__13812 (
            .O(N__64593),
            .I(N__64590));
    LocalMux I__13811 (
            .O(N__64590),
            .I(N__64587));
    Span4Mux_h I__13810 (
            .O(N__64587),
            .I(N__64584));
    Odrv4 I__13809 (
            .O(N__64584),
            .I(\pid_side.pid_preregZ0Z_22 ));
    InMux I__13808 (
            .O(N__64581),
            .I(\pid_side.un1_pid_prereg_0_cry_21 ));
    InMux I__13807 (
            .O(N__64578),
            .I(N__64575));
    LocalMux I__13806 (
            .O(N__64575),
            .I(\pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ));
    CascadeMux I__13805 (
            .O(N__64572),
            .I(N__64569));
    InMux I__13804 (
            .O(N__64569),
            .I(N__64566));
    LocalMux I__13803 (
            .O(N__64566),
            .I(\pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ));
    CascadeMux I__13802 (
            .O(N__64563),
            .I(N__64560));
    InMux I__13801 (
            .O(N__64560),
            .I(N__64557));
    LocalMux I__13800 (
            .O(N__64557),
            .I(N__64554));
    Span4Mux_v I__13799 (
            .O(N__64554),
            .I(N__64551));
    Odrv4 I__13798 (
            .O(N__64551),
            .I(\pid_side.pid_preregZ0Z_23 ));
    InMux I__13797 (
            .O(N__64548),
            .I(bfn_17_16_0_));
    InMux I__13796 (
            .O(N__64545),
            .I(N__64542));
    LocalMux I__13795 (
            .O(N__64542),
            .I(\pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ));
    CascadeMux I__13794 (
            .O(N__64539),
            .I(N__64536));
    InMux I__13793 (
            .O(N__64536),
            .I(N__64533));
    LocalMux I__13792 (
            .O(N__64533),
            .I(\pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ));
    InMux I__13791 (
            .O(N__64530),
            .I(N__64527));
    LocalMux I__13790 (
            .O(N__64527),
            .I(N__64524));
    Span4Mux_h I__13789 (
            .O(N__64524),
            .I(N__64521));
    Odrv4 I__13788 (
            .O(N__64521),
            .I(\pid_side.pid_preregZ0Z_24 ));
    InMux I__13787 (
            .O(N__64518),
            .I(\pid_side.un1_pid_prereg_0_cry_23 ));
    InMux I__13786 (
            .O(N__64515),
            .I(N__64512));
    LocalMux I__13785 (
            .O(N__64512),
            .I(\pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ));
    CascadeMux I__13784 (
            .O(N__64509),
            .I(N__64506));
    InMux I__13783 (
            .O(N__64506),
            .I(N__64503));
    LocalMux I__13782 (
            .O(N__64503),
            .I(\pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ));
    InMux I__13781 (
            .O(N__64500),
            .I(N__64497));
    LocalMux I__13780 (
            .O(N__64497),
            .I(N__64494));
    Span4Mux_v I__13779 (
            .O(N__64494),
            .I(N__64491));
    Odrv4 I__13778 (
            .O(N__64491),
            .I(\pid_side.pid_preregZ0Z_25 ));
    InMux I__13777 (
            .O(N__64488),
            .I(\pid_side.un1_pid_prereg_0_cry_24 ));
    CascadeMux I__13776 (
            .O(N__64485),
            .I(N__64482));
    InMux I__13775 (
            .O(N__64482),
            .I(N__64479));
    LocalMux I__13774 (
            .O(N__64479),
            .I(\pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ));
    InMux I__13773 (
            .O(N__64476),
            .I(N__64473));
    LocalMux I__13772 (
            .O(N__64473),
            .I(N__64470));
    Span4Mux_v I__13771 (
            .O(N__64470),
            .I(N__64467));
    Odrv4 I__13770 (
            .O(N__64467),
            .I(\pid_side.pid_preregZ0Z_26 ));
    InMux I__13769 (
            .O(N__64464),
            .I(\pid_side.un1_pid_prereg_0_cry_25 ));
    InMux I__13768 (
            .O(N__64461),
            .I(N__64458));
    LocalMux I__13767 (
            .O(N__64458),
            .I(N__64455));
    Odrv4 I__13766 (
            .O(N__64455),
            .I(\pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ));
    CascadeMux I__13765 (
            .O(N__64452),
            .I(N__64449));
    InMux I__13764 (
            .O(N__64449),
            .I(N__64446));
    LocalMux I__13763 (
            .O(N__64446),
            .I(N__64443));
    Span4Mux_h I__13762 (
            .O(N__64443),
            .I(N__64440));
    Odrv4 I__13761 (
            .O(N__64440),
            .I(\pid_side.pid_preregZ0Z_27 ));
    InMux I__13760 (
            .O(N__64437),
            .I(\pid_side.un1_pid_prereg_0_cry_26 ));
    InMux I__13759 (
            .O(N__64434),
            .I(N__64431));
    LocalMux I__13758 (
            .O(N__64431),
            .I(N__64428));
    Odrv4 I__13757 (
            .O(N__64428),
            .I(\pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ));
    CascadeMux I__13756 (
            .O(N__64425),
            .I(N__64422));
    InMux I__13755 (
            .O(N__64422),
            .I(N__64419));
    LocalMux I__13754 (
            .O(N__64419),
            .I(N__64416));
    Odrv4 I__13753 (
            .O(N__64416),
            .I(\pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ));
    InMux I__13752 (
            .O(N__64413),
            .I(N__64410));
    LocalMux I__13751 (
            .O(N__64410),
            .I(N__64407));
    Span4Mux_v I__13750 (
            .O(N__64407),
            .I(N__64404));
    Odrv4 I__13749 (
            .O(N__64404),
            .I(\pid_side.pid_preregZ0Z_28 ));
    InMux I__13748 (
            .O(N__64401),
            .I(\pid_side.un1_pid_prereg_0_cry_27 ));
    InMux I__13747 (
            .O(N__64398),
            .I(\pid_side.un1_pid_prereg_0_cry_12 ));
    InMux I__13746 (
            .O(N__64395),
            .I(N__64392));
    LocalMux I__13745 (
            .O(N__64392),
            .I(N__64389));
    Odrv4 I__13744 (
            .O(N__64389),
            .I(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__13743 (
            .O(N__64386),
            .I(\pid_side.un1_pid_prereg_0_cry_13 ));
    InMux I__13742 (
            .O(N__64383),
            .I(N__64380));
    LocalMux I__13741 (
            .O(N__64380),
            .I(\pid_side.error_d_reg_prev_esr_RNINPDOKZ0Z_12 ));
    InMux I__13740 (
            .O(N__64377),
            .I(N__64371));
    InMux I__13739 (
            .O(N__64376),
            .I(N__64371));
    LocalMux I__13738 (
            .O(N__64371),
            .I(N__64368));
    Odrv4 I__13737 (
            .O(N__64368),
            .I(\pid_side.pid_preregZ0Z_15 ));
    InMux I__13736 (
            .O(N__64365),
            .I(bfn_17_15_0_));
    InMux I__13735 (
            .O(N__64362),
            .I(N__64359));
    LocalMux I__13734 (
            .O(N__64359),
            .I(\pid_side.error_d_reg_prev_esr_RNITHHEAZ0Z_12 ));
    CascadeMux I__13733 (
            .O(N__64356),
            .I(N__64353));
    InMux I__13732 (
            .O(N__64353),
            .I(N__64350));
    LocalMux I__13731 (
            .O(N__64350),
            .I(\pid_side.error_d_reg_prev_esr_RNIJ1F8FZ0Z_12 ));
    InMux I__13730 (
            .O(N__64347),
            .I(N__64341));
    InMux I__13729 (
            .O(N__64346),
            .I(N__64341));
    LocalMux I__13728 (
            .O(N__64341),
            .I(N__64338));
    Odrv4 I__13727 (
            .O(N__64338),
            .I(\pid_side.pid_preregZ0Z_16 ));
    InMux I__13726 (
            .O(N__64335),
            .I(\pid_side.un1_pid_prereg_0_cry_15 ));
    InMux I__13725 (
            .O(N__64332),
            .I(N__64329));
    LocalMux I__13724 (
            .O(N__64329),
            .I(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ));
    CascadeMux I__13723 (
            .O(N__64326),
            .I(N__64323));
    InMux I__13722 (
            .O(N__64323),
            .I(N__64320));
    LocalMux I__13721 (
            .O(N__64320),
            .I(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ));
    InMux I__13720 (
            .O(N__64317),
            .I(N__64311));
    InMux I__13719 (
            .O(N__64316),
            .I(N__64311));
    LocalMux I__13718 (
            .O(N__64311),
            .I(N__64308));
    Odrv4 I__13717 (
            .O(N__64308),
            .I(\pid_side.pid_preregZ0Z_17 ));
    InMux I__13716 (
            .O(N__64305),
            .I(\pid_side.un1_pid_prereg_0_cry_16 ));
    CascadeMux I__13715 (
            .O(N__64302),
            .I(N__64299));
    InMux I__13714 (
            .O(N__64299),
            .I(N__64296));
    LocalMux I__13713 (
            .O(N__64296),
            .I(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ));
    InMux I__13712 (
            .O(N__64293),
            .I(N__64287));
    InMux I__13711 (
            .O(N__64292),
            .I(N__64287));
    LocalMux I__13710 (
            .O(N__64287),
            .I(N__64284));
    Odrv4 I__13709 (
            .O(N__64284),
            .I(\pid_side.pid_preregZ0Z_18 ));
    InMux I__13708 (
            .O(N__64281),
            .I(\pid_side.un1_pid_prereg_0_cry_17 ));
    CascadeMux I__13707 (
            .O(N__64278),
            .I(N__64274));
    InMux I__13706 (
            .O(N__64277),
            .I(N__64269));
    InMux I__13705 (
            .O(N__64274),
            .I(N__64269));
    LocalMux I__13704 (
            .O(N__64269),
            .I(N__64266));
    Odrv12 I__13703 (
            .O(N__64266),
            .I(\pid_side.pid_preregZ0Z_19 ));
    InMux I__13702 (
            .O(N__64263),
            .I(\pid_side.un1_pid_prereg_0_cry_18 ));
    InMux I__13701 (
            .O(N__64260),
            .I(N__64257));
    LocalMux I__13700 (
            .O(N__64257),
            .I(N__64254));
    Span4Mux_h I__13699 (
            .O(N__64254),
            .I(N__64251));
    Odrv4 I__13698 (
            .O(N__64251),
            .I(\pid_side.pid_preregZ0Z_20 ));
    InMux I__13697 (
            .O(N__64248),
            .I(\pid_side.un1_pid_prereg_0_cry_19 ));
    CascadeMux I__13696 (
            .O(N__64245),
            .I(N__64242));
    InMux I__13695 (
            .O(N__64242),
            .I(N__64239));
    LocalMux I__13694 (
            .O(N__64239),
            .I(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ));
    CascadeMux I__13693 (
            .O(N__64236),
            .I(N__64232));
    CascadeMux I__13692 (
            .O(N__64235),
            .I(N__64229));
    InMux I__13691 (
            .O(N__64232),
            .I(N__64226));
    InMux I__13690 (
            .O(N__64229),
            .I(N__64222));
    LocalMux I__13689 (
            .O(N__64226),
            .I(N__64219));
    CascadeMux I__13688 (
            .O(N__64225),
            .I(N__64216));
    LocalMux I__13687 (
            .O(N__64222),
            .I(N__64213));
    Span4Mux_h I__13686 (
            .O(N__64219),
            .I(N__64209));
    InMux I__13685 (
            .O(N__64216),
            .I(N__64206));
    Span4Mux_v I__13684 (
            .O(N__64213),
            .I(N__64203));
    InMux I__13683 (
            .O(N__64212),
            .I(N__64200));
    Odrv4 I__13682 (
            .O(N__64209),
            .I(\pid_side.pid_preregZ0Z_5 ));
    LocalMux I__13681 (
            .O(N__64206),
            .I(\pid_side.pid_preregZ0Z_5 ));
    Odrv4 I__13680 (
            .O(N__64203),
            .I(\pid_side.pid_preregZ0Z_5 ));
    LocalMux I__13679 (
            .O(N__64200),
            .I(\pid_side.pid_preregZ0Z_5 ));
    InMux I__13678 (
            .O(N__64191),
            .I(\pid_side.un1_pid_prereg_0_cry_4 ));
    InMux I__13677 (
            .O(N__64188),
            .I(N__64185));
    LocalMux I__13676 (
            .O(N__64185),
            .I(N__64180));
    InMux I__13675 (
            .O(N__64184),
            .I(N__64175));
    InMux I__13674 (
            .O(N__64183),
            .I(N__64175));
    Odrv4 I__13673 (
            .O(N__64180),
            .I(\pid_side.pid_preregZ0Z_6 ));
    LocalMux I__13672 (
            .O(N__64175),
            .I(\pid_side.pid_preregZ0Z_6 ));
    InMux I__13671 (
            .O(N__64170),
            .I(\pid_side.un1_pid_prereg_0_cry_5 ));
    InMux I__13670 (
            .O(N__64167),
            .I(N__64164));
    LocalMux I__13669 (
            .O(N__64164),
            .I(N__64160));
    CascadeMux I__13668 (
            .O(N__64163),
            .I(N__64156));
    Span4Mux_v I__13667 (
            .O(N__64160),
            .I(N__64153));
    InMux I__13666 (
            .O(N__64159),
            .I(N__64148));
    InMux I__13665 (
            .O(N__64156),
            .I(N__64148));
    Span4Mux_h I__13664 (
            .O(N__64153),
            .I(N__64145));
    LocalMux I__13663 (
            .O(N__64148),
            .I(N__64142));
    Odrv4 I__13662 (
            .O(N__64145),
            .I(\pid_side.pid_preregZ0Z_7 ));
    Odrv4 I__13661 (
            .O(N__64142),
            .I(\pid_side.pid_preregZ0Z_7 ));
    InMux I__13660 (
            .O(N__64137),
            .I(bfn_17_14_0_));
    InMux I__13659 (
            .O(N__64134),
            .I(N__64131));
    LocalMux I__13658 (
            .O(N__64131),
            .I(N__64128));
    Span4Mux_v I__13657 (
            .O(N__64128),
            .I(N__64123));
    InMux I__13656 (
            .O(N__64127),
            .I(N__64118));
    InMux I__13655 (
            .O(N__64126),
            .I(N__64118));
    Span4Mux_h I__13654 (
            .O(N__64123),
            .I(N__64115));
    LocalMux I__13653 (
            .O(N__64118),
            .I(N__64112));
    Odrv4 I__13652 (
            .O(N__64115),
            .I(\pid_side.pid_preregZ0Z_8 ));
    Odrv4 I__13651 (
            .O(N__64112),
            .I(\pid_side.pid_preregZ0Z_8 ));
    InMux I__13650 (
            .O(N__64107),
            .I(\pid_side.un1_pid_prereg_0_cry_7 ));
    InMux I__13649 (
            .O(N__64104),
            .I(\pid_side.un1_pid_prereg_0_cry_8 ));
    InMux I__13648 (
            .O(N__64101),
            .I(N__64096));
    InMux I__13647 (
            .O(N__64100),
            .I(N__64091));
    InMux I__13646 (
            .O(N__64099),
            .I(N__64091));
    LocalMux I__13645 (
            .O(N__64096),
            .I(N__64088));
    LocalMux I__13644 (
            .O(N__64091),
            .I(N__64085));
    Span4Mux_h I__13643 (
            .O(N__64088),
            .I(N__64082));
    Span4Mux_v I__13642 (
            .O(N__64085),
            .I(N__64079));
    Odrv4 I__13641 (
            .O(N__64082),
            .I(\pid_side.pid_preregZ0Z_10 ));
    Odrv4 I__13640 (
            .O(N__64079),
            .I(\pid_side.pid_preregZ0Z_10 ));
    InMux I__13639 (
            .O(N__64074),
            .I(\pid_side.un1_pid_prereg_0_cry_9 ));
    CascadeMux I__13638 (
            .O(N__64071),
            .I(N__64068));
    InMux I__13637 (
            .O(N__64068),
            .I(N__64065));
    LocalMux I__13636 (
            .O(N__64065),
            .I(N__64062));
    Span4Mux_h I__13635 (
            .O(N__64062),
            .I(N__64059));
    Odrv4 I__13634 (
            .O(N__64059),
            .I(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ));
    InMux I__13633 (
            .O(N__64056),
            .I(N__64051));
    CascadeMux I__13632 (
            .O(N__64055),
            .I(N__64048));
    CascadeMux I__13631 (
            .O(N__64054),
            .I(N__64045));
    LocalMux I__13630 (
            .O(N__64051),
            .I(N__64042));
    InMux I__13629 (
            .O(N__64048),
            .I(N__64037));
    InMux I__13628 (
            .O(N__64045),
            .I(N__64037));
    Span4Mux_h I__13627 (
            .O(N__64042),
            .I(N__64034));
    LocalMux I__13626 (
            .O(N__64037),
            .I(N__64031));
    Odrv4 I__13625 (
            .O(N__64034),
            .I(\pid_side.pid_preregZ0Z_11 ));
    Odrv4 I__13624 (
            .O(N__64031),
            .I(\pid_side.pid_preregZ0Z_11 ));
    InMux I__13623 (
            .O(N__64026),
            .I(\pid_side.un1_pid_prereg_0_cry_10 ));
    CascadeMux I__13622 (
            .O(N__64023),
            .I(N__64019));
    InMux I__13621 (
            .O(N__64022),
            .I(N__64015));
    InMux I__13620 (
            .O(N__64019),
            .I(N__64012));
    CascadeMux I__13619 (
            .O(N__64018),
            .I(N__64007));
    LocalMux I__13618 (
            .O(N__64015),
            .I(N__64002));
    LocalMux I__13617 (
            .O(N__64012),
            .I(N__64002));
    InMux I__13616 (
            .O(N__64011),
            .I(N__63997));
    InMux I__13615 (
            .O(N__64010),
            .I(N__63997));
    InMux I__13614 (
            .O(N__64007),
            .I(N__63994));
    Span4Mux_h I__13613 (
            .O(N__64002),
            .I(N__63991));
    LocalMux I__13612 (
            .O(N__63997),
            .I(N__63986));
    LocalMux I__13611 (
            .O(N__63994),
            .I(N__63986));
    Odrv4 I__13610 (
            .O(N__63991),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv4 I__13609 (
            .O(N__63986),
            .I(\pid_side.pid_preregZ0Z_12 ));
    InMux I__13608 (
            .O(N__63981),
            .I(\pid_side.un1_pid_prereg_0_cry_11 ));
    InMux I__13607 (
            .O(N__63978),
            .I(N__63973));
    InMux I__13606 (
            .O(N__63977),
            .I(N__63968));
    InMux I__13605 (
            .O(N__63976),
            .I(N__63968));
    LocalMux I__13604 (
            .O(N__63973),
            .I(\pid_side.pid_preregZ0Z_14 ));
    LocalMux I__13603 (
            .O(N__63968),
            .I(\pid_side.pid_preregZ0Z_14 ));
    CascadeMux I__13602 (
            .O(N__63963),
            .I(\pid_side.pid_prereg_esr_RNIE1A2Z0Z_17_cascade_ ));
    InMux I__13601 (
            .O(N__63960),
            .I(N__63956));
    InMux I__13600 (
            .O(N__63959),
            .I(N__63953));
    LocalMux I__13599 (
            .O(N__63956),
            .I(N__63950));
    LocalMux I__13598 (
            .O(N__63953),
            .I(N__63947));
    Span4Mux_v I__13597 (
            .O(N__63950),
            .I(N__63944));
    Span4Mux_h I__13596 (
            .O(N__63947),
            .I(N__63941));
    Odrv4 I__13595 (
            .O(N__63944),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ));
    Odrv4 I__13594 (
            .O(N__63941),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ));
    InMux I__13593 (
            .O(N__63936),
            .I(N__63933));
    LocalMux I__13592 (
            .O(N__63933),
            .I(N__63930));
    Span4Mux_v I__13591 (
            .O(N__63930),
            .I(N__63925));
    InMux I__13590 (
            .O(N__63929),
            .I(N__63920));
    InMux I__13589 (
            .O(N__63928),
            .I(N__63920));
    Odrv4 I__13588 (
            .O(N__63925),
            .I(\pid_side.pid_preregZ0Z_0 ));
    LocalMux I__13587 (
            .O(N__63920),
            .I(\pid_side.pid_preregZ0Z_0 ));
    InMux I__13586 (
            .O(N__63915),
            .I(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__13585 (
            .O(N__63912),
            .I(\pid_side.un1_pid_prereg_0_cry_0 ));
    InMux I__13584 (
            .O(N__63909),
            .I(\pid_side.un1_pid_prereg_0_cry_1 ));
    CascadeMux I__13583 (
            .O(N__63906),
            .I(N__63903));
    InMux I__13582 (
            .O(N__63903),
            .I(N__63900));
    LocalMux I__13581 (
            .O(N__63900),
            .I(N__63897));
    Odrv4 I__13580 (
            .O(N__63897),
            .I(\pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ));
    InMux I__13579 (
            .O(N__63894),
            .I(\pid_side.un1_pid_prereg_0_cry_2 ));
    InMux I__13578 (
            .O(N__63891),
            .I(N__63888));
    LocalMux I__13577 (
            .O(N__63888),
            .I(\pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ));
    CascadeMux I__13576 (
            .O(N__63885),
            .I(N__63881));
    InMux I__13575 (
            .O(N__63884),
            .I(N__63878));
    InMux I__13574 (
            .O(N__63881),
            .I(N__63875));
    LocalMux I__13573 (
            .O(N__63878),
            .I(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ));
    LocalMux I__13572 (
            .O(N__63875),
            .I(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ));
    InMux I__13571 (
            .O(N__63870),
            .I(N__63867));
    LocalMux I__13570 (
            .O(N__63867),
            .I(N__63862));
    InMux I__13569 (
            .O(N__63866),
            .I(N__63859));
    CascadeMux I__13568 (
            .O(N__63865),
            .I(N__63856));
    Span4Mux_v I__13567 (
            .O(N__63862),
            .I(N__63850));
    LocalMux I__13566 (
            .O(N__63859),
            .I(N__63850));
    InMux I__13565 (
            .O(N__63856),
            .I(N__63845));
    InMux I__13564 (
            .O(N__63855),
            .I(N__63845));
    Odrv4 I__13563 (
            .O(N__63850),
            .I(\pid_side.pid_preregZ0Z_4 ));
    LocalMux I__13562 (
            .O(N__63845),
            .I(\pid_side.pid_preregZ0Z_4 ));
    InMux I__13561 (
            .O(N__63840),
            .I(\pid_side.un1_pid_prereg_0_cry_3 ));
    InMux I__13560 (
            .O(N__63837),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__13559 (
            .O(N__63834),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    CascadeMux I__13558 (
            .O(N__63831),
            .I(N__63828));
    InMux I__13557 (
            .O(N__63828),
            .I(N__63825));
    LocalMux I__13556 (
            .O(N__63825),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ));
    InMux I__13555 (
            .O(N__63822),
            .I(N__63819));
    LocalMux I__13554 (
            .O(N__63819),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    IoInMux I__13553 (
            .O(N__63816),
            .I(N__63813));
    LocalMux I__13552 (
            .O(N__63813),
            .I(N__63810));
    Span4Mux_s3_v I__13551 (
            .O(N__63810),
            .I(N__63807));
    Sp12to4 I__13550 (
            .O(N__63807),
            .I(N__63804));
    Span12Mux_h I__13549 (
            .O(N__63804),
            .I(N__63801));
    Span12Mux_v I__13548 (
            .O(N__63801),
            .I(N__63798));
    Odrv12 I__13547 (
            .O(N__63798),
            .I(\pid_side.state_RNIIIOOZ0Z_0 ));
    InMux I__13546 (
            .O(N__63795),
            .I(N__63792));
    LocalMux I__13545 (
            .O(N__63792),
            .I(N__63789));
    Span4Mux_v I__13544 (
            .O(N__63789),
            .I(N__63786));
    Span4Mux_v I__13543 (
            .O(N__63786),
            .I(N__63783));
    Odrv4 I__13542 (
            .O(N__63783),
            .I(\pid_side.N_61_0 ));
    InMux I__13541 (
            .O(N__63780),
            .I(N__63777));
    LocalMux I__13540 (
            .O(N__63777),
            .I(N__63774));
    Odrv4 I__13539 (
            .O(N__63774),
            .I(\pid_side.un11lto30_i_a2_2_and ));
    InMux I__13538 (
            .O(N__63771),
            .I(N__63768));
    LocalMux I__13537 (
            .O(N__63768),
            .I(N__63765));
    Odrv4 I__13536 (
            .O(N__63765),
            .I(\pid_side.un11lto30_i_a2_3_and ));
    InMux I__13535 (
            .O(N__63762),
            .I(N__63759));
    LocalMux I__13534 (
            .O(N__63759),
            .I(N__63756));
    Odrv4 I__13533 (
            .O(N__63756),
            .I(\ppm_encoder_1.throttle_RNIB72M6Z0Z_8 ));
    InMux I__13532 (
            .O(N__63753),
            .I(bfn_17_9_0_));
    InMux I__13531 (
            .O(N__63750),
            .I(N__63747));
    LocalMux I__13530 (
            .O(N__63747),
            .I(N__63744));
    Odrv4 I__13529 (
            .O(N__63744),
            .I(\ppm_encoder_1.throttle_RNIGC2M6Z0Z_9 ));
    InMux I__13528 (
            .O(N__63741),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__13527 (
            .O(N__63738),
            .I(N__63735));
    LocalMux I__13526 (
            .O(N__63735),
            .I(\ppm_encoder_1.elevator_RNIOVAA6Z0Z_10 ));
    InMux I__13525 (
            .O(N__63732),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__13524 (
            .O(N__63729),
            .I(N__63726));
    LocalMux I__13523 (
            .O(N__63726),
            .I(N__63723));
    Odrv12 I__13522 (
            .O(N__63723),
            .I(\ppm_encoder_1.elevator_RNIT4BA6Z0Z_11 ));
    InMux I__13521 (
            .O(N__63720),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__13520 (
            .O(N__63717),
            .I(N__63714));
    LocalMux I__13519 (
            .O(N__63714),
            .I(N__63711));
    Span4Mux_h I__13518 (
            .O(N__63711),
            .I(N__63708));
    Odrv4 I__13517 (
            .O(N__63708),
            .I(\ppm_encoder_1.elevator_RNI2ABA6Z0Z_12 ));
    InMux I__13516 (
            .O(N__63705),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__13515 (
            .O(N__63702),
            .I(N__63699));
    LocalMux I__13514 (
            .O(N__63699),
            .I(N__63696));
    Span4Mux_v I__13513 (
            .O(N__63696),
            .I(N__63693));
    Odrv4 I__13512 (
            .O(N__63693),
            .I(\ppm_encoder_1.elevator_RNI7FBA6Z0Z_13 ));
    InMux I__13511 (
            .O(N__63690),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    CascadeMux I__13510 (
            .O(N__63687),
            .I(N__63684));
    InMux I__13509 (
            .O(N__63684),
            .I(N__63681));
    LocalMux I__13508 (
            .O(N__63681),
            .I(N__63678));
    Odrv4 I__13507 (
            .O(N__63678),
            .I(\ppm_encoder_1.aileron_esr_RNIG1J17Z0Z_14 ));
    InMux I__13506 (
            .O(N__63675),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__13505 (
            .O(N__63672),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__13504 (
            .O(N__63669),
            .I(N__63666));
    LocalMux I__13503 (
            .O(N__63666),
            .I(N__63663));
    Odrv12 I__13502 (
            .O(N__63663),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__13501 (
            .O(N__63660),
            .I(bfn_17_10_0_));
    InMux I__13500 (
            .O(N__63657),
            .I(N__63654));
    LocalMux I__13499 (
            .O(N__63654),
            .I(\ppm_encoder_1.aileron_RNI2Q3U4Z0Z_0 ));
    InMux I__13498 (
            .O(N__63651),
            .I(N__63648));
    LocalMux I__13497 (
            .O(N__63648),
            .I(N__63645));
    Odrv4 I__13496 (
            .O(N__63645),
            .I(\ppm_encoder_1.throttle_RNIFL0A6Z0Z_1 ));
    CascadeMux I__13495 (
            .O(N__63642),
            .I(N__63638));
    InMux I__13494 (
            .O(N__63641),
            .I(N__63635));
    InMux I__13493 (
            .O(N__63638),
            .I(N__63632));
    LocalMux I__13492 (
            .O(N__63635),
            .I(N__63629));
    LocalMux I__13491 (
            .O(N__63632),
            .I(N__63626));
    Span4Mux_v I__13490 (
            .O(N__63629),
            .I(N__63621));
    Span4Mux_v I__13489 (
            .O(N__63626),
            .I(N__63621));
    Odrv4 I__13488 (
            .O(N__63621),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    InMux I__13487 (
            .O(N__63618),
            .I(N__63615));
    LocalMux I__13486 (
            .O(N__63615),
            .I(N__63612));
    Span4Mux_v I__13485 (
            .O(N__63612),
            .I(N__63609));
    Odrv4 I__13484 (
            .O(N__63609),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__13483 (
            .O(N__63606),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__13482 (
            .O(N__63603),
            .I(N__63600));
    LocalMux I__13481 (
            .O(N__63600),
            .I(\ppm_encoder_1.aileron_RNIA24U4Z0Z_2 ));
    InMux I__13480 (
            .O(N__63597),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__13479 (
            .O(N__63594),
            .I(N__63591));
    LocalMux I__13478 (
            .O(N__63591),
            .I(\ppm_encoder_1.aileron_RNIE64U4Z0Z_3 ));
    InMux I__13477 (
            .O(N__63588),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__13476 (
            .O(N__63585),
            .I(N__63582));
    LocalMux I__13475 (
            .O(N__63582),
            .I(N__63579));
    Odrv4 I__13474 (
            .O(N__63579),
            .I(\ppm_encoder_1.elevator_RNI0L5L6Z0Z_4 ));
    InMux I__13473 (
            .O(N__63576),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__13472 (
            .O(N__63573),
            .I(N__63570));
    LocalMux I__13471 (
            .O(N__63570),
            .I(N__63567));
    Odrv4 I__13470 (
            .O(N__63567),
            .I(\ppm_encoder_1.elevator_RNI5Q5L6Z0Z_5 ));
    InMux I__13469 (
            .O(N__63564),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__13468 (
            .O(N__63561),
            .I(N__63558));
    LocalMux I__13467 (
            .O(N__63558),
            .I(N__63555));
    Span4Mux_h I__13466 (
            .O(N__63555),
            .I(N__63552));
    Odrv4 I__13465 (
            .O(N__63552),
            .I(\ppm_encoder_1.throttle_RNI1T1M6Z0Z_6 ));
    InMux I__13464 (
            .O(N__63549),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__13463 (
            .O(N__63546),
            .I(N__63543));
    LocalMux I__13462 (
            .O(N__63543),
            .I(N__63540));
    Span4Mux_h I__13461 (
            .O(N__63540),
            .I(N__63537));
    Odrv4 I__13460 (
            .O(N__63537),
            .I(\ppm_encoder_1.throttle_RNI622M6Z0Z_7 ));
    InMux I__13459 (
            .O(N__63534),
            .I(N__63530));
    CascadeMux I__13458 (
            .O(N__63533),
            .I(N__63527));
    LocalMux I__13457 (
            .O(N__63530),
            .I(N__63524));
    InMux I__13456 (
            .O(N__63527),
            .I(N__63521));
    Span4Mux_h I__13455 (
            .O(N__63524),
            .I(N__63516));
    LocalMux I__13454 (
            .O(N__63521),
            .I(N__63516));
    Span4Mux_h I__13453 (
            .O(N__63516),
            .I(N__63513));
    Span4Mux_v I__13452 (
            .O(N__63513),
            .I(N__63510));
    Odrv4 I__13451 (
            .O(N__63510),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    InMux I__13450 (
            .O(N__63507),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__13449 (
            .O(N__63504),
            .I(N__63495));
    InMux I__13448 (
            .O(N__63503),
            .I(N__63492));
    InMux I__13447 (
            .O(N__63502),
            .I(N__63485));
    InMux I__13446 (
            .O(N__63501),
            .I(N__63482));
    InMux I__13445 (
            .O(N__63500),
            .I(N__63479));
    InMux I__13444 (
            .O(N__63499),
            .I(N__63476));
    InMux I__13443 (
            .O(N__63498),
            .I(N__63473));
    LocalMux I__13442 (
            .O(N__63495),
            .I(N__63470));
    LocalMux I__13441 (
            .O(N__63492),
            .I(N__63467));
    InMux I__13440 (
            .O(N__63491),
            .I(N__63464));
    InMux I__13439 (
            .O(N__63490),
            .I(N__63459));
    InMux I__13438 (
            .O(N__63489),
            .I(N__63454));
    InMux I__13437 (
            .O(N__63488),
            .I(N__63454));
    LocalMux I__13436 (
            .O(N__63485),
            .I(N__63447));
    LocalMux I__13435 (
            .O(N__63482),
            .I(N__63447));
    LocalMux I__13434 (
            .O(N__63479),
            .I(N__63447));
    LocalMux I__13433 (
            .O(N__63476),
            .I(N__63434));
    LocalMux I__13432 (
            .O(N__63473),
            .I(N__63434));
    Span4Mux_h I__13431 (
            .O(N__63470),
            .I(N__63434));
    Span4Mux_h I__13430 (
            .O(N__63467),
            .I(N__63434));
    LocalMux I__13429 (
            .O(N__63464),
            .I(N__63434));
    InMux I__13428 (
            .O(N__63463),
            .I(N__63429));
    InMux I__13427 (
            .O(N__63462),
            .I(N__63426));
    LocalMux I__13426 (
            .O(N__63459),
            .I(N__63421));
    LocalMux I__13425 (
            .O(N__63454),
            .I(N__63421));
    Span4Mux_v I__13424 (
            .O(N__63447),
            .I(N__63416));
    InMux I__13423 (
            .O(N__63446),
            .I(N__63413));
    InMux I__13422 (
            .O(N__63445),
            .I(N__63410));
    Span4Mux_v I__13421 (
            .O(N__63434),
            .I(N__63407));
    InMux I__13420 (
            .O(N__63433),
            .I(N__63402));
    InMux I__13419 (
            .O(N__63432),
            .I(N__63402));
    LocalMux I__13418 (
            .O(N__63429),
            .I(N__63395));
    LocalMux I__13417 (
            .O(N__63426),
            .I(N__63395));
    Span4Mux_h I__13416 (
            .O(N__63421),
            .I(N__63395));
    InMux I__13415 (
            .O(N__63420),
            .I(N__63390));
    InMux I__13414 (
            .O(N__63419),
            .I(N__63390));
    Span4Mux_h I__13413 (
            .O(N__63416),
            .I(N__63385));
    LocalMux I__13412 (
            .O(N__63413),
            .I(N__63385));
    LocalMux I__13411 (
            .O(N__63410),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__13410 (
            .O(N__63407),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__13409 (
            .O(N__63402),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__13408 (
            .O(N__63395),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__13407 (
            .O(N__63390),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__13406 (
            .O(N__63385),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__13405 (
            .O(N__63372),
            .I(N__63365));
    InMux I__13404 (
            .O(N__63371),
            .I(N__63357));
    InMux I__13403 (
            .O(N__63370),
            .I(N__63352));
    InMux I__13402 (
            .O(N__63369),
            .I(N__63352));
    InMux I__13401 (
            .O(N__63368),
            .I(N__63349));
    LocalMux I__13400 (
            .O(N__63365),
            .I(N__63346));
    InMux I__13399 (
            .O(N__63364),
            .I(N__63343));
    InMux I__13398 (
            .O(N__63363),
            .I(N__63339));
    InMux I__13397 (
            .O(N__63362),
            .I(N__63336));
    InMux I__13396 (
            .O(N__63361),
            .I(N__63333));
    InMux I__13395 (
            .O(N__63360),
            .I(N__63330));
    LocalMux I__13394 (
            .O(N__63357),
            .I(N__63321));
    LocalMux I__13393 (
            .O(N__63352),
            .I(N__63321));
    LocalMux I__13392 (
            .O(N__63349),
            .I(N__63318));
    Span4Mux_h I__13391 (
            .O(N__63346),
            .I(N__63313));
    LocalMux I__13390 (
            .O(N__63343),
            .I(N__63313));
    InMux I__13389 (
            .O(N__63342),
            .I(N__63310));
    LocalMux I__13388 (
            .O(N__63339),
            .I(N__63307));
    LocalMux I__13387 (
            .O(N__63336),
            .I(N__63300));
    LocalMux I__13386 (
            .O(N__63333),
            .I(N__63300));
    LocalMux I__13385 (
            .O(N__63330),
            .I(N__63300));
    InMux I__13384 (
            .O(N__63329),
            .I(N__63295));
    InMux I__13383 (
            .O(N__63328),
            .I(N__63295));
    InMux I__13382 (
            .O(N__63327),
            .I(N__63292));
    InMux I__13381 (
            .O(N__63326),
            .I(N__63289));
    Span4Mux_v I__13380 (
            .O(N__63321),
            .I(N__63280));
    Span4Mux_h I__13379 (
            .O(N__63318),
            .I(N__63280));
    Span4Mux_v I__13378 (
            .O(N__63313),
            .I(N__63280));
    LocalMux I__13377 (
            .O(N__63310),
            .I(N__63280));
    Odrv4 I__13376 (
            .O(N__63307),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__13375 (
            .O(N__63300),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__13374 (
            .O(N__63295),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__13373 (
            .O(N__63292),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__13372 (
            .O(N__63289),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__13371 (
            .O(N__63280),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__13370 (
            .O(N__63267),
            .I(N__63260));
    InMux I__13369 (
            .O(N__63266),
            .I(N__63254));
    InMux I__13368 (
            .O(N__63265),
            .I(N__63251));
    InMux I__13367 (
            .O(N__63264),
            .I(N__63246));
    InMux I__13366 (
            .O(N__63263),
            .I(N__63243));
    LocalMux I__13365 (
            .O(N__63260),
            .I(N__63240));
    InMux I__13364 (
            .O(N__63259),
            .I(N__63235));
    InMux I__13363 (
            .O(N__63258),
            .I(N__63235));
    InMux I__13362 (
            .O(N__63257),
            .I(N__63232));
    LocalMux I__13361 (
            .O(N__63254),
            .I(N__63227));
    LocalMux I__13360 (
            .O(N__63251),
            .I(N__63227));
    InMux I__13359 (
            .O(N__63250),
            .I(N__63224));
    InMux I__13358 (
            .O(N__63249),
            .I(N__63219));
    LocalMux I__13357 (
            .O(N__63246),
            .I(N__63214));
    LocalMux I__13356 (
            .O(N__63243),
            .I(N__63205));
    Span4Mux_v I__13355 (
            .O(N__63240),
            .I(N__63205));
    LocalMux I__13354 (
            .O(N__63235),
            .I(N__63205));
    LocalMux I__13353 (
            .O(N__63232),
            .I(N__63205));
    Span4Mux_v I__13352 (
            .O(N__63227),
            .I(N__63200));
    LocalMux I__13351 (
            .O(N__63224),
            .I(N__63200));
    InMux I__13350 (
            .O(N__63223),
            .I(N__63197));
    InMux I__13349 (
            .O(N__63222),
            .I(N__63194));
    LocalMux I__13348 (
            .O(N__63219),
            .I(N__63191));
    InMux I__13347 (
            .O(N__63218),
            .I(N__63188));
    InMux I__13346 (
            .O(N__63217),
            .I(N__63185));
    Odrv4 I__13345 (
            .O(N__63214),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__13344 (
            .O(N__63205),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__13343 (
            .O(N__63200),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__13342 (
            .O(N__63197),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__13341 (
            .O(N__63194),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__13340 (
            .O(N__63191),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__13339 (
            .O(N__63188),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__13338 (
            .O(N__63185),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    CascadeMux I__13337 (
            .O(N__63168),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ));
    InMux I__13336 (
            .O(N__63165),
            .I(N__63157));
    InMux I__13335 (
            .O(N__63164),
            .I(N__63152));
    InMux I__13334 (
            .O(N__63163),
            .I(N__63149));
    InMux I__13333 (
            .O(N__63162),
            .I(N__63145));
    InMux I__13332 (
            .O(N__63161),
            .I(N__63138));
    InMux I__13331 (
            .O(N__63160),
            .I(N__63135));
    LocalMux I__13330 (
            .O(N__63157),
            .I(N__63132));
    InMux I__13329 (
            .O(N__63156),
            .I(N__63129));
    InMux I__13328 (
            .O(N__63155),
            .I(N__63126));
    LocalMux I__13327 (
            .O(N__63152),
            .I(N__63121));
    LocalMux I__13326 (
            .O(N__63149),
            .I(N__63121));
    InMux I__13325 (
            .O(N__63148),
            .I(N__63118));
    LocalMux I__13324 (
            .O(N__63145),
            .I(N__63113));
    InMux I__13323 (
            .O(N__63144),
            .I(N__63108));
    InMux I__13322 (
            .O(N__63143),
            .I(N__63108));
    InMux I__13321 (
            .O(N__63142),
            .I(N__63103));
    InMux I__13320 (
            .O(N__63141),
            .I(N__63103));
    LocalMux I__13319 (
            .O(N__63138),
            .I(N__63100));
    LocalMux I__13318 (
            .O(N__63135),
            .I(N__63091));
    Span4Mux_v I__13317 (
            .O(N__63132),
            .I(N__63091));
    LocalMux I__13316 (
            .O(N__63129),
            .I(N__63091));
    LocalMux I__13315 (
            .O(N__63126),
            .I(N__63091));
    Span4Mux_v I__13314 (
            .O(N__63121),
            .I(N__63086));
    LocalMux I__13313 (
            .O(N__63118),
            .I(N__63086));
    InMux I__13312 (
            .O(N__63117),
            .I(N__63081));
    InMux I__13311 (
            .O(N__63116),
            .I(N__63081));
    Odrv4 I__13310 (
            .O(N__63113),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__13309 (
            .O(N__63108),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__13308 (
            .O(N__63103),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__13307 (
            .O(N__63100),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__13306 (
            .O(N__63091),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__13305 (
            .O(N__63086),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__13304 (
            .O(N__63081),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    InMux I__13303 (
            .O(N__63066),
            .I(N__63063));
    LocalMux I__13302 (
            .O(N__63063),
            .I(\ppm_encoder_1.N_288 ));
    CascadeMux I__13301 (
            .O(N__63060),
            .I(N__63056));
    InMux I__13300 (
            .O(N__63059),
            .I(N__63051));
    InMux I__13299 (
            .O(N__63056),
            .I(N__63048));
    InMux I__13298 (
            .O(N__63055),
            .I(N__63041));
    InMux I__13297 (
            .O(N__63054),
            .I(N__63038));
    LocalMux I__13296 (
            .O(N__63051),
            .I(N__63029));
    LocalMux I__13295 (
            .O(N__63048),
            .I(N__63029));
    InMux I__13294 (
            .O(N__63047),
            .I(N__63026));
    InMux I__13293 (
            .O(N__63046),
            .I(N__63023));
    InMux I__13292 (
            .O(N__63045),
            .I(N__63020));
    InMux I__13291 (
            .O(N__63044),
            .I(N__63017));
    LocalMux I__13290 (
            .O(N__63041),
            .I(N__63014));
    LocalMux I__13289 (
            .O(N__63038),
            .I(N__63011));
    InMux I__13288 (
            .O(N__63037),
            .I(N__63008));
    InMux I__13287 (
            .O(N__63036),
            .I(N__63003));
    InMux I__13286 (
            .O(N__63035),
            .I(N__63003));
    InMux I__13285 (
            .O(N__63034),
            .I(N__63000));
    Span4Mux_h I__13284 (
            .O(N__63029),
            .I(N__62991));
    LocalMux I__13283 (
            .O(N__63026),
            .I(N__62988));
    LocalMux I__13282 (
            .O(N__63023),
            .I(N__62981));
    LocalMux I__13281 (
            .O(N__63020),
            .I(N__62981));
    LocalMux I__13280 (
            .O(N__63017),
            .I(N__62981));
    Span4Mux_h I__13279 (
            .O(N__63014),
            .I(N__62972));
    Span4Mux_v I__13278 (
            .O(N__63011),
            .I(N__62972));
    LocalMux I__13277 (
            .O(N__63008),
            .I(N__62972));
    LocalMux I__13276 (
            .O(N__63003),
            .I(N__62972));
    LocalMux I__13275 (
            .O(N__63000),
            .I(N__62969));
    InMux I__13274 (
            .O(N__62999),
            .I(N__62966));
    InMux I__13273 (
            .O(N__62998),
            .I(N__62963));
    CascadeMux I__13272 (
            .O(N__62997),
            .I(N__62960));
    CascadeMux I__13271 (
            .O(N__62996),
            .I(N__62957));
    CascadeMux I__13270 (
            .O(N__62995),
            .I(N__62953));
    CascadeMux I__13269 (
            .O(N__62994),
            .I(N__62949));
    Sp12to4 I__13268 (
            .O(N__62991),
            .I(N__62943));
    Span12Mux_h I__13267 (
            .O(N__62988),
            .I(N__62943));
    Span4Mux_v I__13266 (
            .O(N__62981),
            .I(N__62940));
    Span4Mux_v I__13265 (
            .O(N__62972),
            .I(N__62937));
    Span4Mux_h I__13264 (
            .O(N__62969),
            .I(N__62930));
    LocalMux I__13263 (
            .O(N__62966),
            .I(N__62930));
    LocalMux I__13262 (
            .O(N__62963),
            .I(N__62930));
    InMux I__13261 (
            .O(N__62960),
            .I(N__62927));
    InMux I__13260 (
            .O(N__62957),
            .I(N__62922));
    InMux I__13259 (
            .O(N__62956),
            .I(N__62922));
    InMux I__13258 (
            .O(N__62953),
            .I(N__62913));
    InMux I__13257 (
            .O(N__62952),
            .I(N__62913));
    InMux I__13256 (
            .O(N__62949),
            .I(N__62913));
    InMux I__13255 (
            .O(N__62948),
            .I(N__62913));
    Odrv12 I__13254 (
            .O(N__62943),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__13253 (
            .O(N__62940),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__13252 (
            .O(N__62937),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__13251 (
            .O(N__62930),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__13250 (
            .O(N__62927),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__13249 (
            .O(N__62922),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__13248 (
            .O(N__62913),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__13247 (
            .O(N__62898),
            .I(N__62895));
    LocalMux I__13246 (
            .O(N__62895),
            .I(N__62892));
    Span4Mux_h I__13245 (
            .O(N__62892),
            .I(N__62889));
    Odrv4 I__13244 (
            .O(N__62889),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__13243 (
            .O(N__62886),
            .I(N__62883));
    LocalMux I__13242 (
            .O(N__62883),
            .I(N__62880));
    Span4Mux_h I__13241 (
            .O(N__62880),
            .I(N__62876));
    InMux I__13240 (
            .O(N__62879),
            .I(N__62873));
    Span4Mux_v I__13239 (
            .O(N__62876),
            .I(N__62868));
    LocalMux I__13238 (
            .O(N__62873),
            .I(N__62868));
    Span4Mux_h I__13237 (
            .O(N__62868),
            .I(N__62865));
    Odrv4 I__13236 (
            .O(N__62865),
            .I(front_order_2));
    InMux I__13235 (
            .O(N__62862),
            .I(N__62859));
    LocalMux I__13234 (
            .O(N__62859),
            .I(N__62856));
    Span4Mux_h I__13233 (
            .O(N__62856),
            .I(N__62853));
    Odrv4 I__13232 (
            .O(N__62853),
            .I(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ));
    CascadeMux I__13231 (
            .O(N__62850),
            .I(N__62847));
    InMux I__13230 (
            .O(N__62847),
            .I(N__62842));
    InMux I__13229 (
            .O(N__62846),
            .I(N__62837));
    InMux I__13228 (
            .O(N__62845),
            .I(N__62837));
    LocalMux I__13227 (
            .O(N__62842),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    LocalMux I__13226 (
            .O(N__62837),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    InMux I__13225 (
            .O(N__62832),
            .I(N__62829));
    LocalMux I__13224 (
            .O(N__62829),
            .I(N__62826));
    Span4Mux_v I__13223 (
            .O(N__62826),
            .I(N__62823));
    Span4Mux_h I__13222 (
            .O(N__62823),
            .I(N__62820));
    Odrv4 I__13221 (
            .O(N__62820),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__13220 (
            .O(N__62817),
            .I(N__62814));
    LocalMux I__13219 (
            .O(N__62814),
            .I(N__62811));
    Span4Mux_v I__13218 (
            .O(N__62811),
            .I(N__62807));
    InMux I__13217 (
            .O(N__62810),
            .I(N__62804));
    Span4Mux_h I__13216 (
            .O(N__62807),
            .I(N__62799));
    LocalMux I__13215 (
            .O(N__62804),
            .I(N__62799));
    Span4Mux_h I__13214 (
            .O(N__62799),
            .I(N__62796));
    Span4Mux_h I__13213 (
            .O(N__62796),
            .I(N__62793));
    Odrv4 I__13212 (
            .O(N__62793),
            .I(throttle_order_2));
    CascadeMux I__13211 (
            .O(N__62790),
            .I(N__62785));
    InMux I__13210 (
            .O(N__62789),
            .I(N__62778));
    InMux I__13209 (
            .O(N__62788),
            .I(N__62778));
    InMux I__13208 (
            .O(N__62785),
            .I(N__62778));
    LocalMux I__13207 (
            .O(N__62778),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__13206 (
            .O(N__62775),
            .I(N__62772));
    LocalMux I__13205 (
            .O(N__62772),
            .I(N__62769));
    Odrv4 I__13204 (
            .O(N__62769),
            .I(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ));
    InMux I__13203 (
            .O(N__62766),
            .I(N__62761));
    InMux I__13202 (
            .O(N__62765),
            .I(N__62756));
    InMux I__13201 (
            .O(N__62764),
            .I(N__62756));
    LocalMux I__13200 (
            .O(N__62761),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    LocalMux I__13199 (
            .O(N__62756),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    CascadeMux I__13198 (
            .O(N__62751),
            .I(N__62746));
    CascadeMux I__13197 (
            .O(N__62750),
            .I(N__62743));
    CascadeMux I__13196 (
            .O(N__62749),
            .I(N__62740));
    InMux I__13195 (
            .O(N__62746),
            .I(N__62734));
    InMux I__13194 (
            .O(N__62743),
            .I(N__62727));
    InMux I__13193 (
            .O(N__62740),
            .I(N__62727));
    InMux I__13192 (
            .O(N__62739),
            .I(N__62727));
    CascadeMux I__13191 (
            .O(N__62738),
            .I(N__62724));
    CascadeMux I__13190 (
            .O(N__62737),
            .I(N__62721));
    LocalMux I__13189 (
            .O(N__62734),
            .I(N__62702));
    LocalMux I__13188 (
            .O(N__62727),
            .I(N__62702));
    InMux I__13187 (
            .O(N__62724),
            .I(N__62695));
    InMux I__13186 (
            .O(N__62721),
            .I(N__62695));
    InMux I__13185 (
            .O(N__62720),
            .I(N__62695));
    CascadeMux I__13184 (
            .O(N__62719),
            .I(N__62690));
    CascadeMux I__13183 (
            .O(N__62718),
            .I(N__62687));
    CascadeMux I__13182 (
            .O(N__62717),
            .I(N__62684));
    CascadeMux I__13181 (
            .O(N__62716),
            .I(N__62679));
    CascadeMux I__13180 (
            .O(N__62715),
            .I(N__62668));
    CascadeMux I__13179 (
            .O(N__62714),
            .I(N__62665));
    CascadeMux I__13178 (
            .O(N__62713),
            .I(N__62662));
    CascadeMux I__13177 (
            .O(N__62712),
            .I(N__62659));
    CascadeMux I__13176 (
            .O(N__62711),
            .I(N__62656));
    CascadeMux I__13175 (
            .O(N__62710),
            .I(N__62649));
    CascadeMux I__13174 (
            .O(N__62709),
            .I(N__62646));
    CascadeMux I__13173 (
            .O(N__62708),
            .I(N__62643));
    CascadeMux I__13172 (
            .O(N__62707),
            .I(N__62640));
    Span4Mux_v I__13171 (
            .O(N__62702),
            .I(N__62634));
    LocalMux I__13170 (
            .O(N__62695),
            .I(N__62634));
    CascadeMux I__13169 (
            .O(N__62694),
            .I(N__62629));
    InMux I__13168 (
            .O(N__62693),
            .I(N__62622));
    InMux I__13167 (
            .O(N__62690),
            .I(N__62622));
    InMux I__13166 (
            .O(N__62687),
            .I(N__62622));
    InMux I__13165 (
            .O(N__62684),
            .I(N__62619));
    InMux I__13164 (
            .O(N__62683),
            .I(N__62612));
    InMux I__13163 (
            .O(N__62682),
            .I(N__62612));
    InMux I__13162 (
            .O(N__62679),
            .I(N__62612));
    InMux I__13161 (
            .O(N__62678),
            .I(N__62605));
    InMux I__13160 (
            .O(N__62677),
            .I(N__62605));
    InMux I__13159 (
            .O(N__62676),
            .I(N__62605));
    CascadeMux I__13158 (
            .O(N__62675),
            .I(N__62601));
    CascadeMux I__13157 (
            .O(N__62674),
            .I(N__62598));
    CascadeMux I__13156 (
            .O(N__62673),
            .I(N__62594));
    InMux I__13155 (
            .O(N__62672),
            .I(N__62583));
    InMux I__13154 (
            .O(N__62671),
            .I(N__62583));
    InMux I__13153 (
            .O(N__62668),
            .I(N__62583));
    InMux I__13152 (
            .O(N__62665),
            .I(N__62578));
    InMux I__13151 (
            .O(N__62662),
            .I(N__62571));
    InMux I__13150 (
            .O(N__62659),
            .I(N__62571));
    InMux I__13149 (
            .O(N__62656),
            .I(N__62571));
    CascadeMux I__13148 (
            .O(N__62655),
            .I(N__62565));
    CascadeMux I__13147 (
            .O(N__62654),
            .I(N__62562));
    CascadeMux I__13146 (
            .O(N__62653),
            .I(N__62559));
    InMux I__13145 (
            .O(N__62652),
            .I(N__62545));
    InMux I__13144 (
            .O(N__62649),
            .I(N__62545));
    InMux I__13143 (
            .O(N__62646),
            .I(N__62545));
    InMux I__13142 (
            .O(N__62643),
            .I(N__62545));
    InMux I__13141 (
            .O(N__62640),
            .I(N__62545));
    InMux I__13140 (
            .O(N__62639),
            .I(N__62545));
    Span4Mux_h I__13139 (
            .O(N__62634),
            .I(N__62542));
    InMux I__13138 (
            .O(N__62633),
            .I(N__62535));
    InMux I__13137 (
            .O(N__62632),
            .I(N__62535));
    InMux I__13136 (
            .O(N__62629),
            .I(N__62535));
    LocalMux I__13135 (
            .O(N__62622),
            .I(N__62530));
    LocalMux I__13134 (
            .O(N__62619),
            .I(N__62530));
    LocalMux I__13133 (
            .O(N__62612),
            .I(N__62525));
    LocalMux I__13132 (
            .O(N__62605),
            .I(N__62525));
    InMux I__13131 (
            .O(N__62604),
            .I(N__62518));
    InMux I__13130 (
            .O(N__62601),
            .I(N__62518));
    InMux I__13129 (
            .O(N__62598),
            .I(N__62518));
    InMux I__13128 (
            .O(N__62597),
            .I(N__62509));
    InMux I__13127 (
            .O(N__62594),
            .I(N__62509));
    InMux I__13126 (
            .O(N__62593),
            .I(N__62509));
    InMux I__13125 (
            .O(N__62592),
            .I(N__62509));
    InMux I__13124 (
            .O(N__62591),
            .I(N__62504));
    InMux I__13123 (
            .O(N__62590),
            .I(N__62504));
    LocalMux I__13122 (
            .O(N__62583),
            .I(N__62501));
    InMux I__13121 (
            .O(N__62582),
            .I(N__62496));
    InMux I__13120 (
            .O(N__62581),
            .I(N__62496));
    LocalMux I__13119 (
            .O(N__62578),
            .I(N__62491));
    LocalMux I__13118 (
            .O(N__62571),
            .I(N__62491));
    InMux I__13117 (
            .O(N__62570),
            .I(N__62476));
    InMux I__13116 (
            .O(N__62569),
            .I(N__62476));
    InMux I__13115 (
            .O(N__62568),
            .I(N__62476));
    InMux I__13114 (
            .O(N__62565),
            .I(N__62476));
    InMux I__13113 (
            .O(N__62562),
            .I(N__62476));
    InMux I__13112 (
            .O(N__62559),
            .I(N__62476));
    InMux I__13111 (
            .O(N__62558),
            .I(N__62476));
    LocalMux I__13110 (
            .O(N__62545),
            .I(N__62471));
    Sp12to4 I__13109 (
            .O(N__62542),
            .I(N__62471));
    LocalMux I__13108 (
            .O(N__62535),
            .I(N__62464));
    Span4Mux_v I__13107 (
            .O(N__62530),
            .I(N__62464));
    Span4Mux_v I__13106 (
            .O(N__62525),
            .I(N__62464));
    LocalMux I__13105 (
            .O(N__62518),
            .I(N__62453));
    LocalMux I__13104 (
            .O(N__62509),
            .I(N__62453));
    LocalMux I__13103 (
            .O(N__62504),
            .I(N__62453));
    Sp12to4 I__13102 (
            .O(N__62501),
            .I(N__62453));
    LocalMux I__13101 (
            .O(N__62496),
            .I(N__62453));
    Span12Mux_h I__13100 (
            .O(N__62491),
            .I(N__62450));
    LocalMux I__13099 (
            .O(N__62476),
            .I(N__62443));
    Span12Mux_v I__13098 (
            .O(N__62471),
            .I(N__62443));
    Sp12to4 I__13097 (
            .O(N__62464),
            .I(N__62443));
    Span12Mux_h I__13096 (
            .O(N__62453),
            .I(N__62440));
    Span12Mux_v I__13095 (
            .O(N__62450),
            .I(N__62437));
    Span12Mux_h I__13094 (
            .O(N__62443),
            .I(N__62434));
    Span12Mux_v I__13093 (
            .O(N__62440),
            .I(N__62431));
    Odrv12 I__13092 (
            .O(N__62437),
            .I(pid_altitude_dv));
    Odrv12 I__13091 (
            .O(N__62434),
            .I(pid_altitude_dv));
    Odrv12 I__13090 (
            .O(N__62431),
            .I(pid_altitude_dv));
    InMux I__13089 (
            .O(N__62424),
            .I(N__62421));
    LocalMux I__13088 (
            .O(N__62421),
            .I(N__62418));
    Span4Mux_v I__13087 (
            .O(N__62418),
            .I(N__62415));
    Span4Mux_h I__13086 (
            .O(N__62415),
            .I(N__62411));
    InMux I__13085 (
            .O(N__62414),
            .I(N__62408));
    Odrv4 I__13084 (
            .O(N__62411),
            .I(scaler_4_data_6));
    LocalMux I__13083 (
            .O(N__62408),
            .I(scaler_4_data_6));
    InMux I__13082 (
            .O(N__62403),
            .I(N__62400));
    LocalMux I__13081 (
            .O(N__62400),
            .I(\pid_side.N_57_0 ));
    InMux I__13080 (
            .O(N__62397),
            .I(N__62394));
    LocalMux I__13079 (
            .O(N__62394),
            .I(\pid_side.N_129 ));
    CascadeMux I__13078 (
            .O(N__62391),
            .I(N__62386));
    InMux I__13077 (
            .O(N__62390),
            .I(N__62383));
    InMux I__13076 (
            .O(N__62389),
            .I(N__62380));
    InMux I__13075 (
            .O(N__62386),
            .I(N__62377));
    LocalMux I__13074 (
            .O(N__62383),
            .I(N__62374));
    LocalMux I__13073 (
            .O(N__62380),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__13072 (
            .O(N__62377),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__13071 (
            .O(N__62374),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__13070 (
            .O(N__62367),
            .I(N__62362));
    InMux I__13069 (
            .O(N__62366),
            .I(N__62359));
    InMux I__13068 (
            .O(N__62365),
            .I(N__62356));
    LocalMux I__13067 (
            .O(N__62362),
            .I(N__62353));
    LocalMux I__13066 (
            .O(N__62359),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__13065 (
            .O(N__62356),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__13064 (
            .O(N__62353),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__13063 (
            .O(N__62346),
            .I(N__62343));
    LocalMux I__13062 (
            .O(N__62343),
            .I(N__62340));
    Span4Mux_h I__13061 (
            .O(N__62340),
            .I(N__62337));
    Odrv4 I__13060 (
            .O(N__62337),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    IoInMux I__13059 (
            .O(N__62334),
            .I(N__62331));
    LocalMux I__13058 (
            .O(N__62331),
            .I(N__62328));
    IoSpan4Mux I__13057 (
            .O(N__62328),
            .I(N__62325));
    Span4Mux_s3_v I__13056 (
            .O(N__62325),
            .I(N__62322));
    Odrv4 I__13055 (
            .O(N__62322),
            .I(\pid_side.state_RNIL5IFZ0Z_0 ));
    InMux I__13054 (
            .O(N__62319),
            .I(N__62315));
    InMux I__13053 (
            .O(N__62318),
            .I(N__62312));
    LocalMux I__13052 (
            .O(N__62315),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    LocalMux I__13051 (
            .O(N__62312),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__13050 (
            .O(N__62307),
            .I(N__62303));
    InMux I__13049 (
            .O(N__62306),
            .I(N__62300));
    LocalMux I__13048 (
            .O(N__62303),
            .I(N__62297));
    LocalMux I__13047 (
            .O(N__62300),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    Odrv4 I__13046 (
            .O(N__62297),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    CascadeMux I__13045 (
            .O(N__62292),
            .I(N__62288));
    CascadeMux I__13044 (
            .O(N__62291),
            .I(N__62285));
    InMux I__13043 (
            .O(N__62288),
            .I(N__62282));
    InMux I__13042 (
            .O(N__62285),
            .I(N__62279));
    LocalMux I__13041 (
            .O(N__62282),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    LocalMux I__13040 (
            .O(N__62279),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    InMux I__13039 (
            .O(N__62274),
            .I(N__62271));
    LocalMux I__13038 (
            .O(N__62271),
            .I(N__62267));
    InMux I__13037 (
            .O(N__62270),
            .I(N__62264));
    Span12Mux_v I__13036 (
            .O(N__62267),
            .I(N__62259));
    LocalMux I__13035 (
            .O(N__62264),
            .I(N__62259));
    Span12Mux_v I__13034 (
            .O(N__62259),
            .I(N__62256));
    Odrv12 I__13033 (
            .O(N__62256),
            .I(xy_kd_1));
    InMux I__13032 (
            .O(N__62253),
            .I(N__62250));
    LocalMux I__13031 (
            .O(N__62250),
            .I(\pid_side.N_58_0 ));
    InMux I__13030 (
            .O(N__62247),
            .I(N__62244));
    LocalMux I__13029 (
            .O(N__62244),
            .I(\pid_side.N_36_0 ));
    CascadeMux I__13028 (
            .O(N__62241),
            .I(\pid_side.N_36_0_cascade_ ));
    CascadeMux I__13027 (
            .O(N__62238),
            .I(\pid_side.N_57_0_cascade_ ));
    InMux I__13026 (
            .O(N__62235),
            .I(N__62232));
    LocalMux I__13025 (
            .O(N__62232),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_24 ));
    InMux I__13024 (
            .O(N__62229),
            .I(N__62223));
    InMux I__13023 (
            .O(N__62228),
            .I(N__62223));
    LocalMux I__13022 (
            .O(N__62223),
            .I(\pid_side.N_29_1 ));
    InMux I__13021 (
            .O(N__62220),
            .I(N__62217));
    LocalMux I__13020 (
            .O(N__62217),
            .I(N__62213));
    InMux I__13019 (
            .O(N__62216),
            .I(N__62210));
    Odrv4 I__13018 (
            .O(N__62213),
            .I(\pid_side.N_32_0 ));
    LocalMux I__13017 (
            .O(N__62210),
            .I(\pid_side.N_32_0 ));
    CascadeMux I__13016 (
            .O(N__62205),
            .I(N__62202));
    InMux I__13015 (
            .O(N__62202),
            .I(N__62199));
    LocalMux I__13014 (
            .O(N__62199),
            .I(N__62196));
    Span4Mux_v I__13013 (
            .O(N__62196),
            .I(N__62193));
    Span4Mux_v I__13012 (
            .O(N__62193),
            .I(N__62190));
    Odrv4 I__13011 (
            .O(N__62190),
            .I(\pid_side.error_i_regZ0Z_8 ));
    InMux I__13010 (
            .O(N__62187),
            .I(N__62184));
    LocalMux I__13009 (
            .O(N__62184),
            .I(N__62181));
    Span4Mux_h I__13008 (
            .O(N__62181),
            .I(N__62178));
    Odrv4 I__13007 (
            .O(N__62178),
            .I(\pid_side.N_60_0 ));
    InMux I__13006 (
            .O(N__62175),
            .I(N__62172));
    LocalMux I__13005 (
            .O(N__62172),
            .I(\pid_side.m0_2_03 ));
    CascadeMux I__13004 (
            .O(N__62169),
            .I(\pid_side.N_60_0_cascade_ ));
    CascadeMux I__13003 (
            .O(N__62166),
            .I(N__62162));
    CascadeMux I__13002 (
            .O(N__62165),
            .I(N__62159));
    InMux I__13001 (
            .O(N__62162),
            .I(N__62156));
    InMux I__13000 (
            .O(N__62159),
            .I(N__62153));
    LocalMux I__12999 (
            .O(N__62156),
            .I(N__62148));
    LocalMux I__12998 (
            .O(N__62153),
            .I(N__62145));
    InMux I__12997 (
            .O(N__62152),
            .I(N__62142));
    InMux I__12996 (
            .O(N__62151),
            .I(N__62134));
    Span4Mux_v I__12995 (
            .O(N__62148),
            .I(N__62127));
    Span4Mux_v I__12994 (
            .O(N__62145),
            .I(N__62127));
    LocalMux I__12993 (
            .O(N__62142),
            .I(N__62127));
    InMux I__12992 (
            .O(N__62141),
            .I(N__62124));
    CascadeMux I__12991 (
            .O(N__62140),
            .I(N__62121));
    CascadeMux I__12990 (
            .O(N__62139),
            .I(N__62118));
    CascadeMux I__12989 (
            .O(N__62138),
            .I(N__62115));
    CascadeMux I__12988 (
            .O(N__62137),
            .I(N__62112));
    LocalMux I__12987 (
            .O(N__62134),
            .I(N__62109));
    Span4Mux_h I__12986 (
            .O(N__62127),
            .I(N__62104));
    LocalMux I__12985 (
            .O(N__62124),
            .I(N__62104));
    InMux I__12984 (
            .O(N__62121),
            .I(N__62098));
    InMux I__12983 (
            .O(N__62118),
            .I(N__62098));
    InMux I__12982 (
            .O(N__62115),
            .I(N__62093));
    InMux I__12981 (
            .O(N__62112),
            .I(N__62093));
    Span4Mux_v I__12980 (
            .O(N__62109),
            .I(N__62088));
    Span4Mux_h I__12979 (
            .O(N__62104),
            .I(N__62088));
    InMux I__12978 (
            .O(N__62103),
            .I(N__62085));
    LocalMux I__12977 (
            .O(N__62098),
            .I(N__62080));
    LocalMux I__12976 (
            .O(N__62093),
            .I(N__62080));
    Span4Mux_v I__12975 (
            .O(N__62088),
            .I(N__62077));
    LocalMux I__12974 (
            .O(N__62085),
            .I(pid_side_N_166_mux));
    Odrv4 I__12973 (
            .O(N__62080),
            .I(pid_side_N_166_mux));
    Odrv4 I__12972 (
            .O(N__62077),
            .I(pid_side_N_166_mux));
    CascadeMux I__12971 (
            .O(N__62070),
            .I(\pid_side.error_i_reg_9_rn_1_12_cascade_ ));
    CascadeMux I__12970 (
            .O(N__62067),
            .I(N__62064));
    InMux I__12969 (
            .O(N__62064),
            .I(N__62061));
    LocalMux I__12968 (
            .O(N__62061),
            .I(N__62058));
    Span4Mux_v I__12967 (
            .O(N__62058),
            .I(N__62055));
    Span4Mux_v I__12966 (
            .O(N__62055),
            .I(N__62052));
    Odrv4 I__12965 (
            .O(N__62052),
            .I(\pid_side.error_i_regZ0Z_12 ));
    InMux I__12964 (
            .O(N__62049),
            .I(N__62045));
    InMux I__12963 (
            .O(N__62048),
            .I(N__62041));
    LocalMux I__12962 (
            .O(N__62045),
            .I(N__62038));
    InMux I__12961 (
            .O(N__62044),
            .I(N__62035));
    LocalMux I__12960 (
            .O(N__62041),
            .I(\pid_side.N_15_0 ));
    Odrv4 I__12959 (
            .O(N__62038),
            .I(\pid_side.N_15_0 ));
    LocalMux I__12958 (
            .O(N__62035),
            .I(\pid_side.N_15_0 ));
    CascadeMux I__12957 (
            .O(N__62028),
            .I(\pid_side.N_27_1_cascade_ ));
    InMux I__12956 (
            .O(N__62025),
            .I(N__62019));
    InMux I__12955 (
            .O(N__62024),
            .I(N__62016));
    CascadeMux I__12954 (
            .O(N__62023),
            .I(N__62013));
    InMux I__12953 (
            .O(N__62022),
            .I(N__62009));
    LocalMux I__12952 (
            .O(N__62019),
            .I(N__62004));
    LocalMux I__12951 (
            .O(N__62016),
            .I(N__62004));
    InMux I__12950 (
            .O(N__62013),
            .I(N__61999));
    InMux I__12949 (
            .O(N__62012),
            .I(N__61999));
    LocalMux I__12948 (
            .O(N__62009),
            .I(N__61994));
    Span4Mux_v I__12947 (
            .O(N__62004),
            .I(N__61994));
    LocalMux I__12946 (
            .O(N__61999),
            .I(\pid_side.N_63 ));
    Odrv4 I__12945 (
            .O(N__61994),
            .I(\pid_side.N_63 ));
    InMux I__12944 (
            .O(N__61989),
            .I(N__61986));
    LocalMux I__12943 (
            .O(N__61986),
            .I(\pid_side.error_i_reg_esr_RNO_3Z0Z_24 ));
    InMux I__12942 (
            .O(N__61983),
            .I(N__61980));
    LocalMux I__12941 (
            .O(N__61980),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_24 ));
    InMux I__12940 (
            .O(N__61977),
            .I(N__61974));
    LocalMux I__12939 (
            .O(N__61974),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_24 ));
    InMux I__12938 (
            .O(N__61971),
            .I(N__61968));
    LocalMux I__12937 (
            .O(N__61968),
            .I(\pid_side.N_27_1 ));
    InMux I__12936 (
            .O(N__61965),
            .I(N__61960));
    InMux I__12935 (
            .O(N__61964),
            .I(N__61955));
    InMux I__12934 (
            .O(N__61963),
            .I(N__61955));
    LocalMux I__12933 (
            .O(N__61960),
            .I(\pid_side.N_28_1 ));
    LocalMux I__12932 (
            .O(N__61955),
            .I(\pid_side.N_28_1 ));
    InMux I__12931 (
            .O(N__61950),
            .I(N__61947));
    LocalMux I__12930 (
            .O(N__61947),
            .I(\pid_side.N_25_0 ));
    CascadeMux I__12929 (
            .O(N__61944),
            .I(\pid_side.N_25_0_cascade_ ));
    InMux I__12928 (
            .O(N__61941),
            .I(N__61938));
    LocalMux I__12927 (
            .O(N__61938),
            .I(N__61933));
    InMux I__12926 (
            .O(N__61937),
            .I(N__61928));
    InMux I__12925 (
            .O(N__61936),
            .I(N__61928));
    Odrv4 I__12924 (
            .O(N__61933),
            .I(\pid_side.N_38_1 ));
    LocalMux I__12923 (
            .O(N__61928),
            .I(\pid_side.N_38_1 ));
    InMux I__12922 (
            .O(N__61923),
            .I(N__61920));
    LocalMux I__12921 (
            .O(N__61920),
            .I(\pid_side.m4_2_03 ));
    CascadeMux I__12920 (
            .O(N__61917),
            .I(\pid_side.error_i_reg_9_rn_0_16_cascade_ ));
    InMux I__12919 (
            .O(N__61914),
            .I(N__61907));
    InMux I__12918 (
            .O(N__61913),
            .I(N__61902));
    InMux I__12917 (
            .O(N__61912),
            .I(N__61902));
    InMux I__12916 (
            .O(N__61911),
            .I(N__61899));
    InMux I__12915 (
            .O(N__61910),
            .I(N__61896));
    LocalMux I__12914 (
            .O(N__61907),
            .I(N__61893));
    LocalMux I__12913 (
            .O(N__61902),
            .I(N__61888));
    LocalMux I__12912 (
            .O(N__61899),
            .I(N__61885));
    LocalMux I__12911 (
            .O(N__61896),
            .I(N__61882));
    Span4Mux_v I__12910 (
            .O(N__61893),
            .I(N__61879));
    InMux I__12909 (
            .O(N__61892),
            .I(N__61876));
    InMux I__12908 (
            .O(N__61891),
            .I(N__61873));
    Span4Mux_h I__12907 (
            .O(N__61888),
            .I(N__61870));
    Span4Mux_h I__12906 (
            .O(N__61885),
            .I(N__61863));
    Span4Mux_v I__12905 (
            .O(N__61882),
            .I(N__61863));
    Span4Mux_h I__12904 (
            .O(N__61879),
            .I(N__61863));
    LocalMux I__12903 (
            .O(N__61876),
            .I(pid_front_error_i_reg_9_sn_19));
    LocalMux I__12902 (
            .O(N__61873),
            .I(pid_front_error_i_reg_9_sn_19));
    Odrv4 I__12901 (
            .O(N__61870),
            .I(pid_front_error_i_reg_9_sn_19));
    Odrv4 I__12900 (
            .O(N__61863),
            .I(pid_front_error_i_reg_9_sn_19));
    CascadeMux I__12899 (
            .O(N__61854),
            .I(N__61851));
    InMux I__12898 (
            .O(N__61851),
            .I(N__61848));
    LocalMux I__12897 (
            .O(N__61848),
            .I(N__61845));
    Span4Mux_v I__12896 (
            .O(N__61845),
            .I(N__61842));
    Odrv4 I__12895 (
            .O(N__61842),
            .I(\pid_side.error_i_regZ0Z_16 ));
    InMux I__12894 (
            .O(N__61839),
            .I(N__61835));
    InMux I__12893 (
            .O(N__61838),
            .I(N__61830));
    LocalMux I__12892 (
            .O(N__61835),
            .I(N__61827));
    CascadeMux I__12891 (
            .O(N__61834),
            .I(N__61824));
    CascadeMux I__12890 (
            .O(N__61833),
            .I(N__61821));
    LocalMux I__12889 (
            .O(N__61830),
            .I(N__61818));
    Span4Mux_v I__12888 (
            .O(N__61827),
            .I(N__61815));
    InMux I__12887 (
            .O(N__61824),
            .I(N__61811));
    InMux I__12886 (
            .O(N__61821),
            .I(N__61806));
    Span4Mux_v I__12885 (
            .O(N__61818),
            .I(N__61802));
    Span4Mux_h I__12884 (
            .O(N__61815),
            .I(N__61799));
    CascadeMux I__12883 (
            .O(N__61814),
            .I(N__61796));
    LocalMux I__12882 (
            .O(N__61811),
            .I(N__61793));
    InMux I__12881 (
            .O(N__61810),
            .I(N__61788));
    InMux I__12880 (
            .O(N__61809),
            .I(N__61788));
    LocalMux I__12879 (
            .O(N__61806),
            .I(N__61785));
    InMux I__12878 (
            .O(N__61805),
            .I(N__61782));
    Span4Mux_h I__12877 (
            .O(N__61802),
            .I(N__61779));
    Span4Mux_h I__12876 (
            .O(N__61799),
            .I(N__61776));
    InMux I__12875 (
            .O(N__61796),
            .I(N__61773));
    Span4Mux_v I__12874 (
            .O(N__61793),
            .I(N__61766));
    LocalMux I__12873 (
            .O(N__61788),
            .I(N__61766));
    Span4Mux_v I__12872 (
            .O(N__61785),
            .I(N__61766));
    LocalMux I__12871 (
            .O(N__61782),
            .I(N__61761));
    Sp12to4 I__12870 (
            .O(N__61779),
            .I(N__61761));
    Span4Mux_h I__12869 (
            .O(N__61776),
            .I(N__61758));
    LocalMux I__12868 (
            .O(N__61773),
            .I(drone_H_disp_front_0));
    Odrv4 I__12867 (
            .O(N__61766),
            .I(drone_H_disp_front_0));
    Odrv12 I__12866 (
            .O(N__61761),
            .I(drone_H_disp_front_0));
    Odrv4 I__12865 (
            .O(N__61758),
            .I(drone_H_disp_front_0));
    CascadeMux I__12864 (
            .O(N__61749),
            .I(N__61746));
    InMux I__12863 (
            .O(N__61746),
            .I(N__61739));
    InMux I__12862 (
            .O(N__61745),
            .I(N__61739));
    InMux I__12861 (
            .O(N__61744),
            .I(N__61735));
    LocalMux I__12860 (
            .O(N__61739),
            .I(N__61732));
    InMux I__12859 (
            .O(N__61738),
            .I(N__61729));
    LocalMux I__12858 (
            .O(N__61735),
            .I(N__61724));
    Span4Mux_v I__12857 (
            .O(N__61732),
            .I(N__61724));
    LocalMux I__12856 (
            .O(N__61729),
            .I(N__61721));
    Span4Mux_h I__12855 (
            .O(N__61724),
            .I(N__61716));
    Span4Mux_v I__12854 (
            .O(N__61721),
            .I(N__61716));
    Odrv4 I__12853 (
            .O(N__61716),
            .I(\pid_front.m0_0_03 ));
    CascadeMux I__12852 (
            .O(N__61713),
            .I(\pid_front.m0_0_03_cascade_ ));
    InMux I__12851 (
            .O(N__61710),
            .I(N__61704));
    InMux I__12850 (
            .O(N__61709),
            .I(N__61704));
    LocalMux I__12849 (
            .O(N__61704),
            .I(N__61701));
    Span4Mux_h I__12848 (
            .O(N__61701),
            .I(N__61698));
    Sp12to4 I__12847 (
            .O(N__61698),
            .I(N__61695));
    Odrv12 I__12846 (
            .O(N__61695),
            .I(\pid_front.un4_error_i_reg_22_nsZ0Z_1 ));
    InMux I__12845 (
            .O(N__61692),
            .I(N__61685));
    InMux I__12844 (
            .O(N__61691),
            .I(N__61685));
    InMux I__12843 (
            .O(N__61690),
            .I(N__61682));
    LocalMux I__12842 (
            .O(N__61685),
            .I(N__61679));
    LocalMux I__12841 (
            .O(N__61682),
            .I(\pid_side.m0_0_03 ));
    Odrv4 I__12840 (
            .O(N__61679),
            .I(\pid_side.m0_0_03 ));
    InMux I__12839 (
            .O(N__61674),
            .I(N__61666));
    InMux I__12838 (
            .O(N__61673),
            .I(N__61661));
    InMux I__12837 (
            .O(N__61672),
            .I(N__61656));
    InMux I__12836 (
            .O(N__61671),
            .I(N__61656));
    CascadeMux I__12835 (
            .O(N__61670),
            .I(N__61652));
    InMux I__12834 (
            .O(N__61669),
            .I(N__61649));
    LocalMux I__12833 (
            .O(N__61666),
            .I(N__61646));
    InMux I__12832 (
            .O(N__61665),
            .I(N__61643));
    InMux I__12831 (
            .O(N__61664),
            .I(N__61640));
    LocalMux I__12830 (
            .O(N__61661),
            .I(N__61629));
    LocalMux I__12829 (
            .O(N__61656),
            .I(N__61629));
    InMux I__12828 (
            .O(N__61655),
            .I(N__61626));
    InMux I__12827 (
            .O(N__61652),
            .I(N__61623));
    LocalMux I__12826 (
            .O(N__61649),
            .I(N__61614));
    Span4Mux_v I__12825 (
            .O(N__61646),
            .I(N__61614));
    LocalMux I__12824 (
            .O(N__61643),
            .I(N__61614));
    LocalMux I__12823 (
            .O(N__61640),
            .I(N__61614));
    InMux I__12822 (
            .O(N__61639),
            .I(N__61609));
    InMux I__12821 (
            .O(N__61638),
            .I(N__61609));
    InMux I__12820 (
            .O(N__61637),
            .I(N__61606));
    InMux I__12819 (
            .O(N__61636),
            .I(N__61602));
    InMux I__12818 (
            .O(N__61635),
            .I(N__61597));
    InMux I__12817 (
            .O(N__61634),
            .I(N__61597));
    Span4Mux_v I__12816 (
            .O(N__61629),
            .I(N__61592));
    LocalMux I__12815 (
            .O(N__61626),
            .I(N__61592));
    LocalMux I__12814 (
            .O(N__61623),
            .I(N__61584));
    Sp12to4 I__12813 (
            .O(N__61614),
            .I(N__61584));
    LocalMux I__12812 (
            .O(N__61609),
            .I(N__61584));
    LocalMux I__12811 (
            .O(N__61606),
            .I(N__61581));
    InMux I__12810 (
            .O(N__61605),
            .I(N__61578));
    LocalMux I__12809 (
            .O(N__61602),
            .I(N__61573));
    LocalMux I__12808 (
            .O(N__61597),
            .I(N__61573));
    Span4Mux_h I__12807 (
            .O(N__61592),
            .I(N__61570));
    InMux I__12806 (
            .O(N__61591),
            .I(N__61567));
    Span12Mux_s6_v I__12805 (
            .O(N__61584),
            .I(N__61562));
    Span12Mux_v I__12804 (
            .O(N__61581),
            .I(N__61562));
    LocalMux I__12803 (
            .O(N__61578),
            .I(N__61559));
    Odrv4 I__12802 (
            .O(N__61573),
            .I(xy_ki_fast_2));
    Odrv4 I__12801 (
            .O(N__61570),
            .I(xy_ki_fast_2));
    LocalMux I__12800 (
            .O(N__61567),
            .I(xy_ki_fast_2));
    Odrv12 I__12799 (
            .O(N__61562),
            .I(xy_ki_fast_2));
    Odrv4 I__12798 (
            .O(N__61559),
            .I(xy_ki_fast_2));
    CascadeMux I__12797 (
            .O(N__61548),
            .I(\pid_side.m0_0_03_cascade_ ));
    CascadeMux I__12796 (
            .O(N__61545),
            .I(\pid_side.N_32_0_cascade_ ));
    InMux I__12795 (
            .O(N__61542),
            .I(N__61538));
    InMux I__12794 (
            .O(N__61541),
            .I(N__61535));
    LocalMux I__12793 (
            .O(N__61538),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    LocalMux I__12792 (
            .O(N__61535),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    CascadeMux I__12791 (
            .O(N__61530),
            .I(\pid_side.m29_2_03_0_cascade_ ));
    CascadeMux I__12790 (
            .O(N__61527),
            .I(N__61524));
    InMux I__12789 (
            .O(N__61524),
            .I(N__61521));
    LocalMux I__12788 (
            .O(N__61521),
            .I(N__61518));
    Odrv4 I__12787 (
            .O(N__61518),
            .I(\pid_side.error_i_regZ0Z_25 ));
    CascadeMux I__12786 (
            .O(N__61515),
            .I(\pid_side.N_117_cascade_ ));
    InMux I__12785 (
            .O(N__61512),
            .I(N__61509));
    LocalMux I__12784 (
            .O(N__61509),
            .I(N__61506));
    Odrv4 I__12783 (
            .O(N__61506),
            .I(\pid_side.N_116_0 ));
    CascadeMux I__12782 (
            .O(N__61503),
            .I(N__61500));
    InMux I__12781 (
            .O(N__61500),
            .I(N__61497));
    LocalMux I__12780 (
            .O(N__61497),
            .I(N__61494));
    Span4Mux_v I__12779 (
            .O(N__61494),
            .I(N__61491));
    Odrv4 I__12778 (
            .O(N__61491),
            .I(\pid_side.error_i_regZ0Z_5 ));
    InMux I__12777 (
            .O(N__61488),
            .I(N__61485));
    LocalMux I__12776 (
            .O(N__61485),
            .I(N__61482));
    Odrv12 I__12775 (
            .O(N__61482),
            .I(\pid_side.N_41_0 ));
    InMux I__12774 (
            .O(N__61479),
            .I(N__61474));
    InMux I__12773 (
            .O(N__61478),
            .I(N__61471));
    InMux I__12772 (
            .O(N__61477),
            .I(N__61468));
    LocalMux I__12771 (
            .O(N__61474),
            .I(\pid_side.N_39_1 ));
    LocalMux I__12770 (
            .O(N__61471),
            .I(\pid_side.N_39_1 ));
    LocalMux I__12769 (
            .O(N__61468),
            .I(\pid_side.N_39_1 ));
    CascadeMux I__12768 (
            .O(N__61461),
            .I(N__61458));
    InMux I__12767 (
            .O(N__61458),
            .I(N__61455));
    LocalMux I__12766 (
            .O(N__61455),
            .I(N__61452));
    Span4Mux_v I__12765 (
            .O(N__61452),
            .I(N__61449));
    Odrv4 I__12764 (
            .O(N__61449),
            .I(\pid_side.error_i_regZ0Z_10 ));
    CascadeMux I__12763 (
            .O(N__61446),
            .I(N__61443));
    InMux I__12762 (
            .O(N__61443),
            .I(N__61440));
    LocalMux I__12761 (
            .O(N__61440),
            .I(N__61437));
    Span4Mux_v I__12760 (
            .O(N__61437),
            .I(N__61434));
    Odrv4 I__12759 (
            .O(N__61434),
            .I(\pid_side.error_i_regZ0Z_4 ));
    InMux I__12758 (
            .O(N__61431),
            .I(N__61428));
    LocalMux I__12757 (
            .O(N__61428),
            .I(N__61425));
    Odrv4 I__12756 (
            .O(N__61425),
            .I(\pid_side.N_55_0 ));
    InMux I__12755 (
            .O(N__61422),
            .I(N__61419));
    LocalMux I__12754 (
            .O(N__61419),
            .I(N__61416));
    Span4Mux_h I__12753 (
            .O(N__61416),
            .I(N__61413));
    Odrv4 I__12752 (
            .O(N__61413),
            .I(\pid_side.N_110 ));
    InMux I__12751 (
            .O(N__61410),
            .I(N__61407));
    LocalMux I__12750 (
            .O(N__61407),
            .I(N__61404));
    Span4Mux_h I__12749 (
            .O(N__61404),
            .I(N__61401));
    Span4Mux_v I__12748 (
            .O(N__61401),
            .I(N__61398));
    Odrv4 I__12747 (
            .O(N__61398),
            .I(\pid_side.error_i_regZ0Z_6 ));
    InMux I__12746 (
            .O(N__61395),
            .I(N__61391));
    InMux I__12745 (
            .O(N__61394),
            .I(N__61388));
    LocalMux I__12744 (
            .O(N__61391),
            .I(N__61383));
    LocalMux I__12743 (
            .O(N__61388),
            .I(N__61383));
    Odrv4 I__12742 (
            .O(N__61383),
            .I(\pid_side.un1_pid_prereg_370_1 ));
    InMux I__12741 (
            .O(N__61380),
            .I(N__61375));
    InMux I__12740 (
            .O(N__61379),
            .I(N__61372));
    InMux I__12739 (
            .O(N__61378),
            .I(N__61369));
    LocalMux I__12738 (
            .O(N__61375),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    LocalMux I__12737 (
            .O(N__61372),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    LocalMux I__12736 (
            .O(N__61369),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    InMux I__12735 (
            .O(N__61362),
            .I(N__61353));
    InMux I__12734 (
            .O(N__61361),
            .I(N__61353));
    InMux I__12733 (
            .O(N__61360),
            .I(N__61348));
    InMux I__12732 (
            .O(N__61359),
            .I(N__61348));
    InMux I__12731 (
            .O(N__61358),
            .I(N__61345));
    LocalMux I__12730 (
            .O(N__61353),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    LocalMux I__12729 (
            .O(N__61348),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    LocalMux I__12728 (
            .O(N__61345),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    CascadeMux I__12727 (
            .O(N__61338),
            .I(\pid_side.un1_pid_prereg_0_25_cascade_ ));
    InMux I__12726 (
            .O(N__61335),
            .I(N__61331));
    InMux I__12725 (
            .O(N__61334),
            .I(N__61328));
    LocalMux I__12724 (
            .O(N__61331),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    LocalMux I__12723 (
            .O(N__61328),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    InMux I__12722 (
            .O(N__61323),
            .I(N__61320));
    LocalMux I__12721 (
            .O(N__61320),
            .I(\pid_side.m11_0_ns_1 ));
    CascadeMux I__12720 (
            .O(N__61317),
            .I(\pid_side.m88_0_ns_1_cascade_ ));
    CascadeMux I__12719 (
            .O(N__61314),
            .I(\pid_side.N_89_0_cascade_ ));
    CascadeMux I__12718 (
            .O(N__61311),
            .I(\pid_side.N_116_0_cascade_ ));
    InMux I__12717 (
            .O(N__61308),
            .I(N__61305));
    LocalMux I__12716 (
            .O(N__61305),
            .I(N__61302));
    Odrv4 I__12715 (
            .O(N__61302),
            .I(\pid_side.error_i_reg_9_rn_2_13 ));
    InMux I__12714 (
            .O(N__61299),
            .I(N__61295));
    InMux I__12713 (
            .O(N__61298),
            .I(N__61292));
    LocalMux I__12712 (
            .O(N__61295),
            .I(\pid_side.un1_pid_prereg_0_11 ));
    LocalMux I__12711 (
            .O(N__61292),
            .I(\pid_side.un1_pid_prereg_0_11 ));
    InMux I__12710 (
            .O(N__61287),
            .I(N__61281));
    InMux I__12709 (
            .O(N__61286),
            .I(N__61281));
    LocalMux I__12708 (
            .O(N__61281),
            .I(\pid_side.un1_pid_prereg_0_10 ));
    CascadeMux I__12707 (
            .O(N__61278),
            .I(\pid_side.un1_pid_prereg_0_12_cascade_ ));
    InMux I__12706 (
            .O(N__61275),
            .I(N__61271));
    InMux I__12705 (
            .O(N__61274),
            .I(N__61268));
    LocalMux I__12704 (
            .O(N__61271),
            .I(N__61262));
    LocalMux I__12703 (
            .O(N__61268),
            .I(N__61262));
    InMux I__12702 (
            .O(N__61267),
            .I(N__61259));
    Odrv4 I__12701 (
            .O(N__61262),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    LocalMux I__12700 (
            .O(N__61259),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    CascadeMux I__12699 (
            .O(N__61254),
            .I(N__61250));
    CascadeMux I__12698 (
            .O(N__61253),
            .I(N__61246));
    InMux I__12697 (
            .O(N__61250),
            .I(N__61241));
    InMux I__12696 (
            .O(N__61249),
            .I(N__61241));
    InMux I__12695 (
            .O(N__61246),
            .I(N__61238));
    LocalMux I__12694 (
            .O(N__61241),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    LocalMux I__12693 (
            .O(N__61238),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    CascadeMux I__12692 (
            .O(N__61233),
            .I(\pid_side.un1_pid_prereg_0_23_cascade_ ));
    InMux I__12691 (
            .O(N__61230),
            .I(N__61225));
    InMux I__12690 (
            .O(N__61229),
            .I(N__61220));
    InMux I__12689 (
            .O(N__61228),
            .I(N__61220));
    LocalMux I__12688 (
            .O(N__61225),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    LocalMux I__12687 (
            .O(N__61220),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    InMux I__12686 (
            .O(N__61215),
            .I(N__61208));
    InMux I__12685 (
            .O(N__61214),
            .I(N__61208));
    InMux I__12684 (
            .O(N__61213),
            .I(N__61205));
    LocalMux I__12683 (
            .O(N__61208),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    LocalMux I__12682 (
            .O(N__61205),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    InMux I__12681 (
            .O(N__61200),
            .I(N__61196));
    InMux I__12680 (
            .O(N__61199),
            .I(N__61193));
    LocalMux I__12679 (
            .O(N__61196),
            .I(\pid_side.un1_pid_prereg_0_23 ));
    LocalMux I__12678 (
            .O(N__61193),
            .I(\pid_side.un1_pid_prereg_0_23 ));
    CascadeMux I__12677 (
            .O(N__61188),
            .I(\pid_side.un1_pid_prereg_0_24_cascade_ ));
    CascadeMux I__12676 (
            .O(N__61185),
            .I(\pid_side.un1_pid_prereg_0_10_cascade_ ));
    InMux I__12675 (
            .O(N__61182),
            .I(N__61177));
    InMux I__12674 (
            .O(N__61181),
            .I(N__61172));
    InMux I__12673 (
            .O(N__61180),
            .I(N__61172));
    LocalMux I__12672 (
            .O(N__61177),
            .I(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ));
    LocalMux I__12671 (
            .O(N__61172),
            .I(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ));
    InMux I__12670 (
            .O(N__61167),
            .I(N__61163));
    InMux I__12669 (
            .O(N__61166),
            .I(N__61160));
    LocalMux I__12668 (
            .O(N__61163),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    LocalMux I__12667 (
            .O(N__61160),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    InMux I__12666 (
            .O(N__61155),
            .I(N__61152));
    LocalMux I__12665 (
            .O(N__61152),
            .I(N__61147));
    InMux I__12664 (
            .O(N__61151),
            .I(N__61142));
    InMux I__12663 (
            .O(N__61150),
            .I(N__61142));
    Odrv4 I__12662 (
            .O(N__61147),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    LocalMux I__12661 (
            .O(N__61142),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    CascadeMux I__12660 (
            .O(N__61137),
            .I(\pid_side.un1_pid_prereg_0_16_cascade_ ));
    InMux I__12659 (
            .O(N__61134),
            .I(N__61129));
    InMux I__12658 (
            .O(N__61133),
            .I(N__61124));
    InMux I__12657 (
            .O(N__61132),
            .I(N__61124));
    LocalMux I__12656 (
            .O(N__61129),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    LocalMux I__12655 (
            .O(N__61124),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    InMux I__12654 (
            .O(N__61119),
            .I(N__61116));
    LocalMux I__12653 (
            .O(N__61116),
            .I(N__61112));
    InMux I__12652 (
            .O(N__61115),
            .I(N__61109));
    Odrv4 I__12651 (
            .O(N__61112),
            .I(\pid_side.un1_pid_prereg_0_16 ));
    LocalMux I__12650 (
            .O(N__61109),
            .I(\pid_side.un1_pid_prereg_0_16 ));
    CascadeMux I__12649 (
            .O(N__61104),
            .I(\pid_side.un1_pid_prereg_0_11_cascade_ ));
    InMux I__12648 (
            .O(N__61101),
            .I(N__61096));
    InMux I__12647 (
            .O(N__61100),
            .I(N__61091));
    InMux I__12646 (
            .O(N__61099),
            .I(N__61091));
    LocalMux I__12645 (
            .O(N__61096),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    LocalMux I__12644 (
            .O(N__61091),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    InMux I__12643 (
            .O(N__61086),
            .I(N__61082));
    InMux I__12642 (
            .O(N__61085),
            .I(N__61079));
    LocalMux I__12641 (
            .O(N__61082),
            .I(N__61076));
    LocalMux I__12640 (
            .O(N__61079),
            .I(N__61073));
    Odrv12 I__12639 (
            .O(N__61076),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    Odrv4 I__12638 (
            .O(N__61073),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    InMux I__12637 (
            .O(N__61068),
            .I(N__61065));
    LocalMux I__12636 (
            .O(N__61065),
            .I(\pid_side.un1_pid_prereg_97 ));
    CascadeMux I__12635 (
            .O(N__61062),
            .I(\pid_side.un1_pid_prereg_0_18_cascade_ ));
    CascadeMux I__12634 (
            .O(N__61059),
            .I(\pid_side.un1_pid_prereg_0_14_cascade_ ));
    InMux I__12633 (
            .O(N__61056),
            .I(N__61051));
    InMux I__12632 (
            .O(N__61055),
            .I(N__61048));
    InMux I__12631 (
            .O(N__61054),
            .I(N__61045));
    LocalMux I__12630 (
            .O(N__61051),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    LocalMux I__12629 (
            .O(N__61048),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    LocalMux I__12628 (
            .O(N__61045),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    InMux I__12627 (
            .O(N__61038),
            .I(N__61034));
    InMux I__12626 (
            .O(N__61037),
            .I(N__61030));
    LocalMux I__12625 (
            .O(N__61034),
            .I(N__61027));
    InMux I__12624 (
            .O(N__61033),
            .I(N__61024));
    LocalMux I__12623 (
            .O(N__61030),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    Odrv4 I__12622 (
            .O(N__61027),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    LocalMux I__12621 (
            .O(N__61024),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    CascadeMux I__12620 (
            .O(N__61017),
            .I(\pid_side.un1_pid_prereg_0_1_cascade_ ));
    InMux I__12619 (
            .O(N__61014),
            .I(N__61011));
    LocalMux I__12618 (
            .O(N__61011),
            .I(N__61007));
    InMux I__12617 (
            .O(N__61010),
            .I(N__61004));
    Odrv4 I__12616 (
            .O(N__61007),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    LocalMux I__12615 (
            .O(N__61004),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    CascadeMux I__12614 (
            .O(N__60999),
            .I(\pid_side.un1_pid_prereg_0_0_cascade_ ));
    InMux I__12613 (
            .O(N__60996),
            .I(N__60992));
    InMux I__12612 (
            .O(N__60995),
            .I(N__60989));
    LocalMux I__12611 (
            .O(N__60992),
            .I(\pid_side.un1_pid_prereg_0_1 ));
    LocalMux I__12610 (
            .O(N__60989),
            .I(\pid_side.un1_pid_prereg_0_1 ));
    InMux I__12609 (
            .O(N__60984),
            .I(N__60980));
    InMux I__12608 (
            .O(N__60983),
            .I(N__60977));
    LocalMux I__12607 (
            .O(N__60980),
            .I(\pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12 ));
    LocalMux I__12606 (
            .O(N__60977),
            .I(\pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12 ));
    InMux I__12605 (
            .O(N__60972),
            .I(N__60968));
    InMux I__12604 (
            .O(N__60971),
            .I(N__60965));
    LocalMux I__12603 (
            .O(N__60968),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ));
    LocalMux I__12602 (
            .O(N__60965),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ));
    CascadeMux I__12601 (
            .O(N__60960),
            .I(\pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12_cascade_ ));
    CascadeMux I__12600 (
            .O(N__60957),
            .I(\pid_side.error_d_reg_prev_esr_RNIG7B43Z0Z_12_cascade_ ));
    CascadeMux I__12599 (
            .O(N__60954),
            .I(\pid_side.un1_pid_prereg_0_19_cascade_ ));
    CascadeMux I__12598 (
            .O(N__60951),
            .I(N__60948));
    InMux I__12597 (
            .O(N__60948),
            .I(N__60942));
    InMux I__12596 (
            .O(N__60947),
            .I(N__60942));
    LocalMux I__12595 (
            .O(N__60942),
            .I(\pid_side.error_d_reg_prevZ0Z_3 ));
    InMux I__12594 (
            .O(N__60939),
            .I(N__60936));
    LocalMux I__12593 (
            .O(N__60936),
            .I(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ));
    InMux I__12592 (
            .O(N__60933),
            .I(N__60928));
    InMux I__12591 (
            .O(N__60932),
            .I(N__60923));
    InMux I__12590 (
            .O(N__60931),
            .I(N__60923));
    LocalMux I__12589 (
            .O(N__60928),
            .I(N__60920));
    LocalMux I__12588 (
            .O(N__60923),
            .I(N__60917));
    Odrv4 I__12587 (
            .O(N__60920),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ));
    Odrv4 I__12586 (
            .O(N__60917),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ));
    CascadeMux I__12585 (
            .O(N__60912),
            .I(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ));
    CascadeMux I__12584 (
            .O(N__60909),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14_cascade_ ));
    CascadeMux I__12583 (
            .O(N__60906),
            .I(\pid_side.un1_pid_prereg_0_2_cascade_ ));
    CascadeMux I__12582 (
            .O(N__60903),
            .I(\pid_side.un1_pid_prereg_0_3_cascade_ ));
    InMux I__12581 (
            .O(N__60900),
            .I(N__60894));
    InMux I__12580 (
            .O(N__60899),
            .I(N__60894));
    LocalMux I__12579 (
            .O(N__60894),
            .I(N__60890));
    InMux I__12578 (
            .O(N__60893),
            .I(N__60887));
    Span4Mux_h I__12577 (
            .O(N__60890),
            .I(N__60884));
    LocalMux I__12576 (
            .O(N__60887),
            .I(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ));
    Odrv4 I__12575 (
            .O(N__60884),
            .I(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ));
    CascadeMux I__12574 (
            .O(N__60879),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ));
    InMux I__12573 (
            .O(N__60876),
            .I(N__60873));
    LocalMux I__12572 (
            .O(N__60873),
            .I(N__60868));
    InMux I__12571 (
            .O(N__60872),
            .I(N__60863));
    InMux I__12570 (
            .O(N__60871),
            .I(N__60863));
    Odrv4 I__12569 (
            .O(N__60868),
            .I(\pid_side.N_99 ));
    LocalMux I__12568 (
            .O(N__60863),
            .I(\pid_side.N_99 ));
    InMux I__12567 (
            .O(N__60858),
            .I(N__60855));
    LocalMux I__12566 (
            .O(N__60855),
            .I(\pid_side.N_11_i ));
    InMux I__12565 (
            .O(N__60852),
            .I(N__60849));
    LocalMux I__12564 (
            .O(N__60849),
            .I(N__60846));
    Span4Mux_h I__12563 (
            .O(N__60846),
            .I(N__60842));
    InMux I__12562 (
            .O(N__60845),
            .I(N__60839));
    Odrv4 I__12561 (
            .O(N__60842),
            .I(side_order_12));
    LocalMux I__12560 (
            .O(N__60839),
            .I(side_order_12));
    InMux I__12559 (
            .O(N__60834),
            .I(N__60831));
    LocalMux I__12558 (
            .O(N__60831),
            .I(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ));
    CascadeMux I__12557 (
            .O(N__60828),
            .I(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ));
    InMux I__12556 (
            .O(N__60825),
            .I(N__60820));
    InMux I__12555 (
            .O(N__60824),
            .I(N__60815));
    InMux I__12554 (
            .O(N__60823),
            .I(N__60815));
    LocalMux I__12553 (
            .O(N__60820),
            .I(N__60812));
    LocalMux I__12552 (
            .O(N__60815),
            .I(N__60809));
    Odrv4 I__12551 (
            .O(N__60812),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    Odrv4 I__12550 (
            .O(N__60809),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    InMux I__12549 (
            .O(N__60804),
            .I(N__60800));
    InMux I__12548 (
            .O(N__60803),
            .I(N__60797));
    LocalMux I__12547 (
            .O(N__60800),
            .I(N__60794));
    LocalMux I__12546 (
            .O(N__60797),
            .I(N__60791));
    Span4Mux_v I__12545 (
            .O(N__60794),
            .I(N__60786));
    Span4Mux_h I__12544 (
            .O(N__60791),
            .I(N__60786));
    Odrv4 I__12543 (
            .O(N__60786),
            .I(side_order_11));
    InMux I__12542 (
            .O(N__60783),
            .I(N__60780));
    LocalMux I__12541 (
            .O(N__60780),
            .I(N__60777));
    Span4Mux_v I__12540 (
            .O(N__60777),
            .I(N__60774));
    Odrv4 I__12539 (
            .O(N__60774),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__12538 (
            .O(N__60771),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__12537 (
            .O(N__60768),
            .I(N__60765));
    LocalMux I__12536 (
            .O(N__60765),
            .I(N__60762));
    Odrv4 I__12535 (
            .O(N__60762),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__12534 (
            .O(N__60759),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__12533 (
            .O(N__60756),
            .I(N__60753));
    LocalMux I__12532 (
            .O(N__60753),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__12531 (
            .O(N__60750),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__12530 (
            .O(N__60747),
            .I(\ppm_encoder_1.un1_aileron_cry_13 ));
    InMux I__12529 (
            .O(N__60744),
            .I(N__60741));
    LocalMux I__12528 (
            .O(N__60741),
            .I(N__60737));
    InMux I__12527 (
            .O(N__60740),
            .I(N__60734));
    Sp12to4 I__12526 (
            .O(N__60737),
            .I(N__60729));
    LocalMux I__12525 (
            .O(N__60734),
            .I(N__60729));
    Odrv12 I__12524 (
            .O(N__60729),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CEMux I__12523 (
            .O(N__60726),
            .I(N__60720));
    CEMux I__12522 (
            .O(N__60725),
            .I(N__60717));
    CEMux I__12521 (
            .O(N__60724),
            .I(N__60714));
    CEMux I__12520 (
            .O(N__60723),
            .I(N__60710));
    LocalMux I__12519 (
            .O(N__60720),
            .I(N__60707));
    LocalMux I__12518 (
            .O(N__60717),
            .I(N__60702));
    LocalMux I__12517 (
            .O(N__60714),
            .I(N__60702));
    CEMux I__12516 (
            .O(N__60713),
            .I(N__60699));
    LocalMux I__12515 (
            .O(N__60710),
            .I(N__60696));
    Span4Mux_v I__12514 (
            .O(N__60707),
            .I(N__60693));
    Span4Mux_v I__12513 (
            .O(N__60702),
            .I(N__60688));
    LocalMux I__12512 (
            .O(N__60699),
            .I(N__60688));
    Span4Mux_h I__12511 (
            .O(N__60696),
            .I(N__60685));
    Span4Mux_h I__12510 (
            .O(N__60693),
            .I(N__60682));
    Span4Mux_h I__12509 (
            .O(N__60688),
            .I(N__60679));
    Span4Mux_v I__12508 (
            .O(N__60685),
            .I(N__60676));
    Odrv4 I__12507 (
            .O(N__60682),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__12506 (
            .O(N__60679),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__12505 (
            .O(N__60676),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    InMux I__12504 (
            .O(N__60669),
            .I(N__60665));
    InMux I__12503 (
            .O(N__60668),
            .I(N__60662));
    LocalMux I__12502 (
            .O(N__60665),
            .I(N__60657));
    LocalMux I__12501 (
            .O(N__60662),
            .I(N__60657));
    Span4Mux_v I__12500 (
            .O(N__60657),
            .I(N__60649));
    InMux I__12499 (
            .O(N__60656),
            .I(N__60646));
    InMux I__12498 (
            .O(N__60655),
            .I(N__60643));
    CascadeMux I__12497 (
            .O(N__60654),
            .I(N__60639));
    CascadeMux I__12496 (
            .O(N__60653),
            .I(N__60636));
    CascadeMux I__12495 (
            .O(N__60652),
            .I(N__60632));
    Span4Mux_v I__12494 (
            .O(N__60649),
            .I(N__60622));
    LocalMux I__12493 (
            .O(N__60646),
            .I(N__60622));
    LocalMux I__12492 (
            .O(N__60643),
            .I(N__60622));
    InMux I__12491 (
            .O(N__60642),
            .I(N__60618));
    InMux I__12490 (
            .O(N__60639),
            .I(N__60613));
    InMux I__12489 (
            .O(N__60636),
            .I(N__60613));
    InMux I__12488 (
            .O(N__60635),
            .I(N__60606));
    InMux I__12487 (
            .O(N__60632),
            .I(N__60606));
    InMux I__12486 (
            .O(N__60631),
            .I(N__60606));
    InMux I__12485 (
            .O(N__60630),
            .I(N__60603));
    CascadeMux I__12484 (
            .O(N__60629),
            .I(N__60599));
    Span4Mux_v I__12483 (
            .O(N__60622),
            .I(N__60590));
    InMux I__12482 (
            .O(N__60621),
            .I(N__60587));
    LocalMux I__12481 (
            .O(N__60618),
            .I(N__60583));
    LocalMux I__12480 (
            .O(N__60613),
            .I(N__60576));
    LocalMux I__12479 (
            .O(N__60606),
            .I(N__60576));
    LocalMux I__12478 (
            .O(N__60603),
            .I(N__60576));
    InMux I__12477 (
            .O(N__60602),
            .I(N__60573));
    InMux I__12476 (
            .O(N__60599),
            .I(N__60567));
    CascadeMux I__12475 (
            .O(N__60598),
            .I(N__60564));
    CascadeMux I__12474 (
            .O(N__60597),
            .I(N__60561));
    CascadeMux I__12473 (
            .O(N__60596),
            .I(N__60557));
    CascadeMux I__12472 (
            .O(N__60595),
            .I(N__60554));
    CascadeMux I__12471 (
            .O(N__60594),
            .I(N__60551));
    CascadeMux I__12470 (
            .O(N__60593),
            .I(N__60548));
    Span4Mux_s1_h I__12469 (
            .O(N__60590),
            .I(N__60542));
    LocalMux I__12468 (
            .O(N__60587),
            .I(N__60542));
    CascadeMux I__12467 (
            .O(N__60586),
            .I(N__60539));
    Span4Mux_s3_h I__12466 (
            .O(N__60583),
            .I(N__60533));
    Span4Mux_v I__12465 (
            .O(N__60576),
            .I(N__60530));
    LocalMux I__12464 (
            .O(N__60573),
            .I(N__60527));
    InMux I__12463 (
            .O(N__60572),
            .I(N__60523));
    IoInMux I__12462 (
            .O(N__60571),
            .I(N__60517));
    InMux I__12461 (
            .O(N__60570),
            .I(N__60514));
    LocalMux I__12460 (
            .O(N__60567),
            .I(N__60511));
    InMux I__12459 (
            .O(N__60564),
            .I(N__60500));
    InMux I__12458 (
            .O(N__60561),
            .I(N__60500));
    InMux I__12457 (
            .O(N__60560),
            .I(N__60500));
    InMux I__12456 (
            .O(N__60557),
            .I(N__60500));
    InMux I__12455 (
            .O(N__60554),
            .I(N__60500));
    InMux I__12454 (
            .O(N__60551),
            .I(N__60495));
    InMux I__12453 (
            .O(N__60548),
            .I(N__60495));
    CascadeMux I__12452 (
            .O(N__60547),
            .I(N__60491));
    Span4Mux_v I__12451 (
            .O(N__60542),
            .I(N__60488));
    InMux I__12450 (
            .O(N__60539),
            .I(N__60485));
    CascadeMux I__12449 (
            .O(N__60538),
            .I(N__60481));
    CascadeMux I__12448 (
            .O(N__60537),
            .I(N__60478));
    CascadeMux I__12447 (
            .O(N__60536),
            .I(N__60475));
    Span4Mux_v I__12446 (
            .O(N__60533),
            .I(N__60468));
    Span4Mux_v I__12445 (
            .O(N__60530),
            .I(N__60468));
    Span4Mux_s3_h I__12444 (
            .O(N__60527),
            .I(N__60468));
    CascadeMux I__12443 (
            .O(N__60526),
            .I(N__60465));
    LocalMux I__12442 (
            .O(N__60523),
            .I(N__60462));
    InMux I__12441 (
            .O(N__60522),
            .I(N__60459));
    InMux I__12440 (
            .O(N__60521),
            .I(N__60456));
    CascadeMux I__12439 (
            .O(N__60520),
            .I(N__60450));
    LocalMux I__12438 (
            .O(N__60517),
            .I(N__60444));
    LocalMux I__12437 (
            .O(N__60514),
            .I(N__60441));
    Span4Mux_h I__12436 (
            .O(N__60511),
            .I(N__60438));
    LocalMux I__12435 (
            .O(N__60500),
            .I(N__60433));
    LocalMux I__12434 (
            .O(N__60495),
            .I(N__60433));
    InMux I__12433 (
            .O(N__60494),
            .I(N__60428));
    InMux I__12432 (
            .O(N__60491),
            .I(N__60428));
    Span4Mux_h I__12431 (
            .O(N__60488),
            .I(N__60425));
    LocalMux I__12430 (
            .O(N__60485),
            .I(N__60422));
    InMux I__12429 (
            .O(N__60484),
            .I(N__60415));
    InMux I__12428 (
            .O(N__60481),
            .I(N__60415));
    InMux I__12427 (
            .O(N__60478),
            .I(N__60415));
    InMux I__12426 (
            .O(N__60475),
            .I(N__60412));
    Span4Mux_h I__12425 (
            .O(N__60468),
            .I(N__60409));
    InMux I__12424 (
            .O(N__60465),
            .I(N__60406));
    Span4Mux_v I__12423 (
            .O(N__60462),
            .I(N__60401));
    LocalMux I__12422 (
            .O(N__60459),
            .I(N__60401));
    LocalMux I__12421 (
            .O(N__60456),
            .I(N__60398));
    InMux I__12420 (
            .O(N__60455),
            .I(N__60395));
    InMux I__12419 (
            .O(N__60454),
            .I(N__60392));
    InMux I__12418 (
            .O(N__60453),
            .I(N__60389));
    InMux I__12417 (
            .O(N__60450),
            .I(N__60386));
    CascadeMux I__12416 (
            .O(N__60449),
            .I(N__60383));
    CascadeMux I__12415 (
            .O(N__60448),
            .I(N__60380));
    CascadeMux I__12414 (
            .O(N__60447),
            .I(N__60377));
    Sp12to4 I__12413 (
            .O(N__60444),
            .I(N__60370));
    Span12Mux_s4_h I__12412 (
            .O(N__60441),
            .I(N__60367));
    Sp12to4 I__12411 (
            .O(N__60438),
            .I(N__60364));
    Span4Mux_h I__12410 (
            .O(N__60433),
            .I(N__60359));
    LocalMux I__12409 (
            .O(N__60428),
            .I(N__60359));
    Span4Mux_h I__12408 (
            .O(N__60425),
            .I(N__60356));
    Span4Mux_h I__12407 (
            .O(N__60422),
            .I(N__60349));
    LocalMux I__12406 (
            .O(N__60415),
            .I(N__60349));
    LocalMux I__12405 (
            .O(N__60412),
            .I(N__60349));
    Span4Mux_h I__12404 (
            .O(N__60409),
            .I(N__60344));
    LocalMux I__12403 (
            .O(N__60406),
            .I(N__60344));
    Sp12to4 I__12402 (
            .O(N__60401),
            .I(N__60335));
    Sp12to4 I__12401 (
            .O(N__60398),
            .I(N__60335));
    LocalMux I__12400 (
            .O(N__60395),
            .I(N__60335));
    LocalMux I__12399 (
            .O(N__60392),
            .I(N__60335));
    LocalMux I__12398 (
            .O(N__60389),
            .I(N__60332));
    LocalMux I__12397 (
            .O(N__60386),
            .I(N__60329));
    InMux I__12396 (
            .O(N__60383),
            .I(N__60326));
    InMux I__12395 (
            .O(N__60380),
            .I(N__60321));
    InMux I__12394 (
            .O(N__60377),
            .I(N__60321));
    CascadeMux I__12393 (
            .O(N__60376),
            .I(N__60318));
    CascadeMux I__12392 (
            .O(N__60375),
            .I(N__60315));
    CascadeMux I__12391 (
            .O(N__60374),
            .I(N__60312));
    CascadeMux I__12390 (
            .O(N__60373),
            .I(N__60309));
    Span12Mux_v I__12389 (
            .O(N__60370),
            .I(N__60302));
    Span12Mux_h I__12388 (
            .O(N__60367),
            .I(N__60302));
    Span12Mux_h I__12387 (
            .O(N__60364),
            .I(N__60302));
    Span4Mux_v I__12386 (
            .O(N__60359),
            .I(N__60299));
    Span4Mux_h I__12385 (
            .O(N__60356),
            .I(N__60294));
    Span4Mux_v I__12384 (
            .O(N__60349),
            .I(N__60294));
    Span4Mux_h I__12383 (
            .O(N__60344),
            .I(N__60291));
    Span12Mux_v I__12382 (
            .O(N__60335),
            .I(N__60280));
    Span12Mux_s0_h I__12381 (
            .O(N__60332),
            .I(N__60280));
    Span12Mux_v I__12380 (
            .O(N__60329),
            .I(N__60280));
    LocalMux I__12379 (
            .O(N__60326),
            .I(N__60280));
    LocalMux I__12378 (
            .O(N__60321),
            .I(N__60280));
    InMux I__12377 (
            .O(N__60318),
            .I(N__60277));
    InMux I__12376 (
            .O(N__60315),
            .I(N__60272));
    InMux I__12375 (
            .O(N__60312),
            .I(N__60272));
    InMux I__12374 (
            .O(N__60309),
            .I(N__60269));
    Odrv12 I__12373 (
            .O(N__60302),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12372 (
            .O(N__60299),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12371 (
            .O(N__60294),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12370 (
            .O(N__60291),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12369 (
            .O(N__60280),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12368 (
            .O(N__60277),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12367 (
            .O(N__60272),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12366 (
            .O(N__60269),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__12365 (
            .O(N__60252),
            .I(N__60249));
    InMux I__12364 (
            .O(N__60249),
            .I(N__60246));
    LocalMux I__12363 (
            .O(N__60246),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a4_4 ));
    InMux I__12362 (
            .O(N__60243),
            .I(N__60240));
    LocalMux I__12361 (
            .O(N__60240),
            .I(\pid_side.source_pid10lt4_0 ));
    InMux I__12360 (
            .O(N__60237),
            .I(N__60234));
    LocalMux I__12359 (
            .O(N__60234),
            .I(N__60231));
    Odrv4 I__12358 (
            .O(N__60231),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a4_3 ));
    InMux I__12357 (
            .O(N__60228),
            .I(N__60225));
    LocalMux I__12356 (
            .O(N__60225),
            .I(\pid_side.un11lto30_i_a2_0_and ));
    InMux I__12355 (
            .O(N__60222),
            .I(N__60219));
    LocalMux I__12354 (
            .O(N__60219),
            .I(N__60216));
    Odrv12 I__12353 (
            .O(N__60216),
            .I(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ));
    InMux I__12352 (
            .O(N__60213),
            .I(\ppm_encoder_1.un1_aileron_cry_2 ));
    InMux I__12351 (
            .O(N__60210),
            .I(N__60207));
    LocalMux I__12350 (
            .O(N__60207),
            .I(N__60203));
    InMux I__12349 (
            .O(N__60206),
            .I(N__60200));
    Span4Mux_h I__12348 (
            .O(N__60203),
            .I(N__60197));
    LocalMux I__12347 (
            .O(N__60200),
            .I(side_order_4));
    Odrv4 I__12346 (
            .O(N__60197),
            .I(side_order_4));
    InMux I__12345 (
            .O(N__60192),
            .I(N__60189));
    LocalMux I__12344 (
            .O(N__60189),
            .I(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ));
    InMux I__12343 (
            .O(N__60186),
            .I(\ppm_encoder_1.un1_aileron_cry_3 ));
    InMux I__12342 (
            .O(N__60183),
            .I(N__60179));
    InMux I__12341 (
            .O(N__60182),
            .I(N__60176));
    LocalMux I__12340 (
            .O(N__60179),
            .I(N__60173));
    LocalMux I__12339 (
            .O(N__60176),
            .I(N__60170));
    Span4Mux_v I__12338 (
            .O(N__60173),
            .I(N__60167));
    Span4Mux_h I__12337 (
            .O(N__60170),
            .I(N__60164));
    Odrv4 I__12336 (
            .O(N__60167),
            .I(side_order_5));
    Odrv4 I__12335 (
            .O(N__60164),
            .I(side_order_5));
    InMux I__12334 (
            .O(N__60159),
            .I(N__60156));
    LocalMux I__12333 (
            .O(N__60156),
            .I(N__60153));
    Odrv4 I__12332 (
            .O(N__60153),
            .I(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ));
    InMux I__12331 (
            .O(N__60150),
            .I(\ppm_encoder_1.un1_aileron_cry_4 ));
    CascadeMux I__12330 (
            .O(N__60147),
            .I(N__60144));
    InMux I__12329 (
            .O(N__60144),
            .I(N__60140));
    InMux I__12328 (
            .O(N__60143),
            .I(N__60137));
    LocalMux I__12327 (
            .O(N__60140),
            .I(N__60134));
    LocalMux I__12326 (
            .O(N__60137),
            .I(N__60131));
    Sp12to4 I__12325 (
            .O(N__60134),
            .I(N__60128));
    Span4Mux_v I__12324 (
            .O(N__60131),
            .I(N__60125));
    Odrv12 I__12323 (
            .O(N__60128),
            .I(side_order_6));
    Odrv4 I__12322 (
            .O(N__60125),
            .I(side_order_6));
    InMux I__12321 (
            .O(N__60120),
            .I(N__60117));
    LocalMux I__12320 (
            .O(N__60117),
            .I(N__60114));
    Span4Mux_h I__12319 (
            .O(N__60114),
            .I(N__60111));
    Odrv4 I__12318 (
            .O(N__60111),
            .I(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ));
    InMux I__12317 (
            .O(N__60108),
            .I(\ppm_encoder_1.un1_aileron_cry_5 ));
    CascadeMux I__12316 (
            .O(N__60105),
            .I(N__60102));
    InMux I__12315 (
            .O(N__60102),
            .I(N__60098));
    InMux I__12314 (
            .O(N__60101),
            .I(N__60095));
    LocalMux I__12313 (
            .O(N__60098),
            .I(N__60092));
    LocalMux I__12312 (
            .O(N__60095),
            .I(N__60089));
    Span4Mux_v I__12311 (
            .O(N__60092),
            .I(N__60086));
    Span4Mux_v I__12310 (
            .O(N__60089),
            .I(N__60083));
    Odrv4 I__12309 (
            .O(N__60086),
            .I(side_order_7));
    Odrv4 I__12308 (
            .O(N__60083),
            .I(side_order_7));
    InMux I__12307 (
            .O(N__60078),
            .I(N__60075));
    LocalMux I__12306 (
            .O(N__60075),
            .I(N__60072));
    Span4Mux_h I__12305 (
            .O(N__60072),
            .I(N__60069));
    Odrv4 I__12304 (
            .O(N__60069),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__12303 (
            .O(N__60066),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__12302 (
            .O(N__60063),
            .I(N__60059));
    InMux I__12301 (
            .O(N__60062),
            .I(N__60056));
    LocalMux I__12300 (
            .O(N__60059),
            .I(N__60053));
    LocalMux I__12299 (
            .O(N__60056),
            .I(N__60050));
    Span4Mux_h I__12298 (
            .O(N__60053),
            .I(N__60047));
    Odrv12 I__12297 (
            .O(N__60050),
            .I(side_order_8));
    Odrv4 I__12296 (
            .O(N__60047),
            .I(side_order_8));
    InMux I__12295 (
            .O(N__60042),
            .I(N__60039));
    LocalMux I__12294 (
            .O(N__60039),
            .I(N__60036));
    Span4Mux_h I__12293 (
            .O(N__60036),
            .I(N__60033));
    Odrv4 I__12292 (
            .O(N__60033),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__12291 (
            .O(N__60030),
            .I(bfn_16_11_0_));
    InMux I__12290 (
            .O(N__60027),
            .I(N__60024));
    LocalMux I__12289 (
            .O(N__60024),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__12288 (
            .O(N__60021),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__12287 (
            .O(N__60018),
            .I(N__60015));
    LocalMux I__12286 (
            .O(N__60015),
            .I(N__60011));
    InMux I__12285 (
            .O(N__60014),
            .I(N__60008));
    Span4Mux_v I__12284 (
            .O(N__60011),
            .I(N__60003));
    LocalMux I__12283 (
            .O(N__60008),
            .I(N__60003));
    Span4Mux_v I__12282 (
            .O(N__60003),
            .I(N__60000));
    Odrv4 I__12281 (
            .O(N__60000),
            .I(side_order_10));
    InMux I__12280 (
            .O(N__59997),
            .I(N__59994));
    LocalMux I__12279 (
            .O(N__59994),
            .I(N__59991));
    Odrv4 I__12278 (
            .O(N__59991),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__12277 (
            .O(N__59988),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__12276 (
            .O(N__59985),
            .I(N__59981));
    CascadeMux I__12275 (
            .O(N__59984),
            .I(N__59977));
    LocalMux I__12274 (
            .O(N__59981),
            .I(N__59974));
    InMux I__12273 (
            .O(N__59980),
            .I(N__59971));
    InMux I__12272 (
            .O(N__59977),
            .I(N__59968));
    Span4Mux_v I__12271 (
            .O(N__59974),
            .I(N__59965));
    LocalMux I__12270 (
            .O(N__59971),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    LocalMux I__12269 (
            .O(N__59968),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__12268 (
            .O(N__59965),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__12267 (
            .O(N__59958),
            .I(N__59953));
    InMux I__12266 (
            .O(N__59957),
            .I(N__59948));
    InMux I__12265 (
            .O(N__59956),
            .I(N__59943));
    LocalMux I__12264 (
            .O(N__59953),
            .I(N__59940));
    InMux I__12263 (
            .O(N__59952),
            .I(N__59937));
    InMux I__12262 (
            .O(N__59951),
            .I(N__59930));
    LocalMux I__12261 (
            .O(N__59948),
            .I(N__59927));
    InMux I__12260 (
            .O(N__59947),
            .I(N__59922));
    InMux I__12259 (
            .O(N__59946),
            .I(N__59922));
    LocalMux I__12258 (
            .O(N__59943),
            .I(N__59919));
    Span4Mux_h I__12257 (
            .O(N__59940),
            .I(N__59916));
    LocalMux I__12256 (
            .O(N__59937),
            .I(N__59913));
    InMux I__12255 (
            .O(N__59936),
            .I(N__59910));
    InMux I__12254 (
            .O(N__59935),
            .I(N__59907));
    InMux I__12253 (
            .O(N__59934),
            .I(N__59904));
    InMux I__12252 (
            .O(N__59933),
            .I(N__59901));
    LocalMux I__12251 (
            .O(N__59930),
            .I(N__59896));
    Span4Mux_h I__12250 (
            .O(N__59927),
            .I(N__59896));
    LocalMux I__12249 (
            .O(N__59922),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__12248 (
            .O(N__59919),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__12247 (
            .O(N__59916),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__12246 (
            .O(N__59913),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__12245 (
            .O(N__59910),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__12244 (
            .O(N__59907),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__12243 (
            .O(N__59904),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__12242 (
            .O(N__59901),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__12241 (
            .O(N__59896),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    CascadeMux I__12240 (
            .O(N__59877),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ));
    InMux I__12239 (
            .O(N__59874),
            .I(N__59871));
    LocalMux I__12238 (
            .O(N__59871),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10 ));
    CascadeMux I__12237 (
            .O(N__59868),
            .I(N__59863));
    CascadeMux I__12236 (
            .O(N__59867),
            .I(N__59860));
    InMux I__12235 (
            .O(N__59866),
            .I(N__59855));
    InMux I__12234 (
            .O(N__59863),
            .I(N__59855));
    InMux I__12233 (
            .O(N__59860),
            .I(N__59852));
    LocalMux I__12232 (
            .O(N__59855),
            .I(N__59849));
    LocalMux I__12231 (
            .O(N__59852),
            .I(N__59846));
    Span4Mux_h I__12230 (
            .O(N__59849),
            .I(N__59843));
    Odrv4 I__12229 (
            .O(N__59846),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__12228 (
            .O(N__59843),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    CascadeMux I__12227 (
            .O(N__59838),
            .I(N__59833));
    InMux I__12226 (
            .O(N__59837),
            .I(N__59830));
    InMux I__12225 (
            .O(N__59836),
            .I(N__59825));
    InMux I__12224 (
            .O(N__59833),
            .I(N__59825));
    LocalMux I__12223 (
            .O(N__59830),
            .I(N__59822));
    LocalMux I__12222 (
            .O(N__59825),
            .I(N__59819));
    Odrv4 I__12221 (
            .O(N__59822),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__12220 (
            .O(N__59819),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    CascadeMux I__12219 (
            .O(N__59814),
            .I(\ppm_encoder_1.N_296_cascade_ ));
    InMux I__12218 (
            .O(N__59811),
            .I(N__59808));
    LocalMux I__12217 (
            .O(N__59808),
            .I(N__59805));
    Span4Mux_h I__12216 (
            .O(N__59805),
            .I(N__59802));
    Odrv4 I__12215 (
            .O(N__59802),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__12214 (
            .O(N__59799),
            .I(N__59790));
    InMux I__12213 (
            .O(N__59798),
            .I(N__59790));
    InMux I__12212 (
            .O(N__59797),
            .I(N__59790));
    LocalMux I__12211 (
            .O(N__59790),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__12210 (
            .O(N__59787),
            .I(N__59784));
    LocalMux I__12209 (
            .O(N__59784),
            .I(N__59780));
    InMux I__12208 (
            .O(N__59783),
            .I(N__59777));
    Span4Mux_h I__12207 (
            .O(N__59780),
            .I(N__59774));
    LocalMux I__12206 (
            .O(N__59777),
            .I(N__59771));
    Span4Mux_v I__12205 (
            .O(N__59774),
            .I(N__59768));
    Span4Mux_h I__12204 (
            .O(N__59771),
            .I(N__59765));
    Odrv4 I__12203 (
            .O(N__59768),
            .I(side_order_0));
    Odrv4 I__12202 (
            .O(N__59765),
            .I(side_order_0));
    InMux I__12201 (
            .O(N__59760),
            .I(N__59757));
    LocalMux I__12200 (
            .O(N__59757),
            .I(N__59754));
    Span4Mux_h I__12199 (
            .O(N__59754),
            .I(N__59751));
    Odrv4 I__12198 (
            .O(N__59751),
            .I(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ));
    InMux I__12197 (
            .O(N__59748),
            .I(\ppm_encoder_1.un1_aileron_cry_0 ));
    InMux I__12196 (
            .O(N__59745),
            .I(\ppm_encoder_1.un1_aileron_cry_1 ));
    CascadeMux I__12195 (
            .O(N__59742),
            .I(\ppm_encoder_1.un1_init_pulses_10_0_cascade_ ));
    InMux I__12194 (
            .O(N__59739),
            .I(N__59736));
    LocalMux I__12193 (
            .O(N__59736),
            .I(N__59733));
    Odrv4 I__12192 (
            .O(N__59733),
            .I(\ppm_encoder_1.N_289 ));
    CascadeMux I__12191 (
            .O(N__59730),
            .I(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ));
    InMux I__12190 (
            .O(N__59727),
            .I(N__59724));
    LocalMux I__12189 (
            .O(N__59724),
            .I(N__59721));
    Span4Mux_h I__12188 (
            .O(N__59721),
            .I(N__59718));
    Odrv4 I__12187 (
            .O(N__59718),
            .I(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ));
    InMux I__12186 (
            .O(N__59715),
            .I(N__59712));
    LocalMux I__12185 (
            .O(N__59712),
            .I(N__59708));
    InMux I__12184 (
            .O(N__59711),
            .I(N__59705));
    Span4Mux_v I__12183 (
            .O(N__59708),
            .I(N__59700));
    LocalMux I__12182 (
            .O(N__59705),
            .I(N__59700));
    Span4Mux_h I__12181 (
            .O(N__59700),
            .I(N__59697));
    Odrv4 I__12180 (
            .O(N__59697),
            .I(front_order_3));
    InMux I__12179 (
            .O(N__59694),
            .I(N__59685));
    InMux I__12178 (
            .O(N__59693),
            .I(N__59685));
    InMux I__12177 (
            .O(N__59692),
            .I(N__59685));
    LocalMux I__12176 (
            .O(N__59685),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    InMux I__12175 (
            .O(N__59682),
            .I(N__59679));
    LocalMux I__12174 (
            .O(N__59679),
            .I(N__59676));
    Span4Mux_h I__12173 (
            .O(N__59676),
            .I(N__59673));
    Odrv4 I__12172 (
            .O(N__59673),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    CascadeMux I__12171 (
            .O(N__59670),
            .I(N__59667));
    InMux I__12170 (
            .O(N__59667),
            .I(N__59664));
    LocalMux I__12169 (
            .O(N__59664),
            .I(N__59660));
    InMux I__12168 (
            .O(N__59663),
            .I(N__59657));
    Span4Mux_v I__12167 (
            .O(N__59660),
            .I(N__59654));
    LocalMux I__12166 (
            .O(N__59657),
            .I(N__59651));
    Span4Mux_h I__12165 (
            .O(N__59654),
            .I(N__59646));
    Span4Mux_v I__12164 (
            .O(N__59651),
            .I(N__59646));
    Span4Mux_h I__12163 (
            .O(N__59646),
            .I(N__59643));
    Odrv4 I__12162 (
            .O(N__59643),
            .I(throttle_order_3));
    CascadeMux I__12161 (
            .O(N__59640),
            .I(N__59635));
    InMux I__12160 (
            .O(N__59639),
            .I(N__59628));
    InMux I__12159 (
            .O(N__59638),
            .I(N__59628));
    InMux I__12158 (
            .O(N__59635),
            .I(N__59628));
    LocalMux I__12157 (
            .O(N__59628),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__12156 (
            .O(N__59625),
            .I(N__59622));
    LocalMux I__12155 (
            .O(N__59622),
            .I(N__59617));
    InMux I__12154 (
            .O(N__59621),
            .I(N__59612));
    InMux I__12153 (
            .O(N__59620),
            .I(N__59612));
    Odrv4 I__12152 (
            .O(N__59617),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    LocalMux I__12151 (
            .O(N__59612),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    CascadeMux I__12150 (
            .O(N__59607),
            .I(N__59604));
    InMux I__12149 (
            .O(N__59604),
            .I(N__59600));
    InMux I__12148 (
            .O(N__59603),
            .I(N__59597));
    LocalMux I__12147 (
            .O(N__59600),
            .I(N__59594));
    LocalMux I__12146 (
            .O(N__59597),
            .I(N__59589));
    Span4Mux_h I__12145 (
            .O(N__59594),
            .I(N__59589));
    Span4Mux_v I__12144 (
            .O(N__59589),
            .I(N__59586));
    Odrv4 I__12143 (
            .O(N__59586),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    InMux I__12142 (
            .O(N__59583),
            .I(N__59580));
    LocalMux I__12141 (
            .O(N__59580),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    InMux I__12140 (
            .O(N__59577),
            .I(N__59574));
    LocalMux I__12139 (
            .O(N__59574),
            .I(N__59571));
    Span4Mux_v I__12138 (
            .O(N__59571),
            .I(N__59568));
    Odrv4 I__12137 (
            .O(N__59568),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    InMux I__12136 (
            .O(N__59565),
            .I(N__59562));
    LocalMux I__12135 (
            .O(N__59562),
            .I(N__59559));
    Span4Mux_h I__12134 (
            .O(N__59559),
            .I(N__59555));
    InMux I__12133 (
            .O(N__59558),
            .I(N__59552));
    Span4Mux_v I__12132 (
            .O(N__59555),
            .I(N__59547));
    LocalMux I__12131 (
            .O(N__59552),
            .I(N__59547));
    Span4Mux_h I__12130 (
            .O(N__59547),
            .I(N__59544));
    Odrv4 I__12129 (
            .O(N__59544),
            .I(front_order_0));
    InMux I__12128 (
            .O(N__59541),
            .I(N__59538));
    LocalMux I__12127 (
            .O(N__59538),
            .I(N__59534));
    InMux I__12126 (
            .O(N__59537),
            .I(N__59531));
    Span4Mux_h I__12125 (
            .O(N__59534),
            .I(N__59528));
    LocalMux I__12124 (
            .O(N__59531),
            .I(N__59525));
    Span4Mux_v I__12123 (
            .O(N__59528),
            .I(N__59522));
    Span4Mux_h I__12122 (
            .O(N__59525),
            .I(N__59519));
    Sp12to4 I__12121 (
            .O(N__59522),
            .I(N__59516));
    Span4Mux_h I__12120 (
            .O(N__59519),
            .I(N__59513));
    Odrv12 I__12119 (
            .O(N__59516),
            .I(throttle_order_0));
    Odrv4 I__12118 (
            .O(N__59513),
            .I(throttle_order_0));
    InMux I__12117 (
            .O(N__59508),
            .I(N__59503));
    InMux I__12116 (
            .O(N__59507),
            .I(N__59498));
    InMux I__12115 (
            .O(N__59506),
            .I(N__59498));
    LocalMux I__12114 (
            .O(N__59503),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    LocalMux I__12113 (
            .O(N__59498),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    CascadeMux I__12112 (
            .O(N__59493),
            .I(N__59488));
    InMux I__12111 (
            .O(N__59492),
            .I(N__59485));
    InMux I__12110 (
            .O(N__59491),
            .I(N__59480));
    InMux I__12109 (
            .O(N__59488),
            .I(N__59480));
    LocalMux I__12108 (
            .O(N__59485),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    LocalMux I__12107 (
            .O(N__59480),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    InMux I__12106 (
            .O(N__59475),
            .I(N__59472));
    LocalMux I__12105 (
            .O(N__59472),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0 ));
    InMux I__12104 (
            .O(N__59469),
            .I(N__59463));
    InMux I__12103 (
            .O(N__59468),
            .I(N__59456));
    InMux I__12102 (
            .O(N__59467),
            .I(N__59456));
    InMux I__12101 (
            .O(N__59466),
            .I(N__59456));
    LocalMux I__12100 (
            .O(N__59463),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    LocalMux I__12099 (
            .O(N__59456),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    CascadeMux I__12098 (
            .O(N__59451),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ));
    CascadeMux I__12097 (
            .O(N__59448),
            .I(N__59445));
    InMux I__12096 (
            .O(N__59445),
            .I(N__59442));
    LocalMux I__12095 (
            .O(N__59442),
            .I(N__59439));
    Span4Mux_h I__12094 (
            .O(N__59439),
            .I(N__59436));
    Span4Mux_v I__12093 (
            .O(N__59436),
            .I(N__59433));
    Span4Mux_h I__12092 (
            .O(N__59433),
            .I(N__59430));
    Odrv4 I__12091 (
            .O(N__59430),
            .I(\pid_front.error_i_regZ0Z_5 ));
    CEMux I__12090 (
            .O(N__59427),
            .I(N__59419));
    CEMux I__12089 (
            .O(N__59426),
            .I(N__59416));
    CEMux I__12088 (
            .O(N__59425),
            .I(N__59413));
    CEMux I__12087 (
            .O(N__59424),
            .I(N__59410));
    CEMux I__12086 (
            .O(N__59423),
            .I(N__59407));
    CEMux I__12085 (
            .O(N__59422),
            .I(N__59404));
    LocalMux I__12084 (
            .O(N__59419),
            .I(N__59400));
    LocalMux I__12083 (
            .O(N__59416),
            .I(N__59397));
    LocalMux I__12082 (
            .O(N__59413),
            .I(N__59394));
    LocalMux I__12081 (
            .O(N__59410),
            .I(N__59391));
    LocalMux I__12080 (
            .O(N__59407),
            .I(N__59386));
    LocalMux I__12079 (
            .O(N__59404),
            .I(N__59386));
    CEMux I__12078 (
            .O(N__59403),
            .I(N__59383));
    Span4Mux_h I__12077 (
            .O(N__59400),
            .I(N__59378));
    Span4Mux_h I__12076 (
            .O(N__59397),
            .I(N__59378));
    Span4Mux_v I__12075 (
            .O(N__59394),
            .I(N__59368));
    Span4Mux_v I__12074 (
            .O(N__59391),
            .I(N__59368));
    Span4Mux_v I__12073 (
            .O(N__59386),
            .I(N__59368));
    LocalMux I__12072 (
            .O(N__59383),
            .I(N__59368));
    Span4Mux_v I__12071 (
            .O(N__59378),
            .I(N__59364));
    CEMux I__12070 (
            .O(N__59377),
            .I(N__59360));
    Span4Mux_h I__12069 (
            .O(N__59368),
            .I(N__59357));
    CEMux I__12068 (
            .O(N__59367),
            .I(N__59354));
    IoSpan4Mux I__12067 (
            .O(N__59364),
            .I(N__59351));
    CEMux I__12066 (
            .O(N__59363),
            .I(N__59348));
    LocalMux I__12065 (
            .O(N__59360),
            .I(N__59342));
    Span4Mux_h I__12064 (
            .O(N__59357),
            .I(N__59337));
    LocalMux I__12063 (
            .O(N__59354),
            .I(N__59337));
    Span4Mux_s2_v I__12062 (
            .O(N__59351),
            .I(N__59331));
    LocalMux I__12061 (
            .O(N__59348),
            .I(N__59331));
    CEMux I__12060 (
            .O(N__59347),
            .I(N__59328));
    CEMux I__12059 (
            .O(N__59346),
            .I(N__59324));
    CEMux I__12058 (
            .O(N__59345),
            .I(N__59321));
    Span4Mux_h I__12057 (
            .O(N__59342),
            .I(N__59318));
    Span4Mux_v I__12056 (
            .O(N__59337),
            .I(N__59315));
    CEMux I__12055 (
            .O(N__59336),
            .I(N__59312));
    Span4Mux_v I__12054 (
            .O(N__59331),
            .I(N__59309));
    LocalMux I__12053 (
            .O(N__59328),
            .I(N__59306));
    CEMux I__12052 (
            .O(N__59327),
            .I(N__59303));
    LocalMux I__12051 (
            .O(N__59324),
            .I(N__59298));
    LocalMux I__12050 (
            .O(N__59321),
            .I(N__59298));
    Span4Mux_v I__12049 (
            .O(N__59318),
            .I(N__59295));
    Span4Mux_h I__12048 (
            .O(N__59315),
            .I(N__59292));
    LocalMux I__12047 (
            .O(N__59312),
            .I(N__59289));
    Span4Mux_h I__12046 (
            .O(N__59309),
            .I(N__59286));
    Span4Mux_h I__12045 (
            .O(N__59306),
            .I(N__59283));
    LocalMux I__12044 (
            .O(N__59303),
            .I(N__59278));
    Sp12to4 I__12043 (
            .O(N__59298),
            .I(N__59278));
    Span4Mux_h I__12042 (
            .O(N__59295),
            .I(N__59275));
    Sp12to4 I__12041 (
            .O(N__59292),
            .I(N__59270));
    Span12Mux_h I__12040 (
            .O(N__59289),
            .I(N__59270));
    Span4Mux_v I__12039 (
            .O(N__59286),
            .I(N__59267));
    Sp12to4 I__12038 (
            .O(N__59283),
            .I(N__59262));
    Span12Mux_s7_v I__12037 (
            .O(N__59278),
            .I(N__59262));
    Span4Mux_v I__12036 (
            .O(N__59275),
            .I(N__59259));
    Span12Mux_v I__12035 (
            .O(N__59270),
            .I(N__59256));
    Span4Mux_v I__12034 (
            .O(N__59267),
            .I(N__59253));
    Odrv12 I__12033 (
            .O(N__59262),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__12032 (
            .O(N__59259),
            .I(\pid_front.state_ns_0_0 ));
    Odrv12 I__12031 (
            .O(N__59256),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__12030 (
            .O(N__59253),
            .I(\pid_front.state_ns_0_0 ));
    InMux I__12029 (
            .O(N__59244),
            .I(N__59241));
    LocalMux I__12028 (
            .O(N__59241),
            .I(N__59236));
    InMux I__12027 (
            .O(N__59240),
            .I(N__59233));
    InMux I__12026 (
            .O(N__59239),
            .I(N__59230));
    Span4Mux_h I__12025 (
            .O(N__59236),
            .I(N__59225));
    LocalMux I__12024 (
            .O(N__59233),
            .I(N__59225));
    LocalMux I__12023 (
            .O(N__59230),
            .I(N__59221));
    Sp12to4 I__12022 (
            .O(N__59225),
            .I(N__59218));
    InMux I__12021 (
            .O(N__59224),
            .I(N__59215));
    Span4Mux_v I__12020 (
            .O(N__59221),
            .I(N__59212));
    Span12Mux_v I__12019 (
            .O(N__59218),
            .I(N__59207));
    LocalMux I__12018 (
            .O(N__59215),
            .I(N__59207));
    Odrv4 I__12017 (
            .O(N__59212),
            .I(pid_side_error_i_reg_9_sn_27));
    Odrv12 I__12016 (
            .O(N__59207),
            .I(pid_side_error_i_reg_9_sn_27));
    InMux I__12015 (
            .O(N__59202),
            .I(N__59195));
    InMux I__12014 (
            .O(N__59201),
            .I(N__59190));
    InMux I__12013 (
            .O(N__59200),
            .I(N__59190));
    InMux I__12012 (
            .O(N__59199),
            .I(N__59187));
    InMux I__12011 (
            .O(N__59198),
            .I(N__59184));
    LocalMux I__12010 (
            .O(N__59195),
            .I(N__59179));
    LocalMux I__12009 (
            .O(N__59190),
            .I(N__59179));
    LocalMux I__12008 (
            .O(N__59187),
            .I(N__59172));
    LocalMux I__12007 (
            .O(N__59184),
            .I(N__59172));
    Span4Mux_h I__12006 (
            .O(N__59179),
            .I(N__59172));
    Odrv4 I__12005 (
            .O(N__59172),
            .I(\pid_front.m2_0_03_3_i_0 ));
    InMux I__12004 (
            .O(N__59169),
            .I(N__59166));
    LocalMux I__12003 (
            .O(N__59166),
            .I(\pid_front.N_55_0 ));
    InMux I__12002 (
            .O(N__59163),
            .I(N__59160));
    LocalMux I__12001 (
            .O(N__59160),
            .I(N__59156));
    InMux I__12000 (
            .O(N__59159),
            .I(N__59153));
    Span4Mux_h I__11999 (
            .O(N__59156),
            .I(N__59149));
    LocalMux I__11998 (
            .O(N__59153),
            .I(N__59146));
    InMux I__11997 (
            .O(N__59152),
            .I(N__59143));
    Span4Mux_h I__11996 (
            .O(N__59149),
            .I(N__59140));
    Span4Mux_h I__11995 (
            .O(N__59146),
            .I(N__59137));
    LocalMux I__11994 (
            .O(N__59143),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__11993 (
            .O(N__59140),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__11992 (
            .O(N__59137),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__11991 (
            .O(N__59130),
            .I(N__59125));
    CascadeMux I__11990 (
            .O(N__59129),
            .I(N__59122));
    CascadeMux I__11989 (
            .O(N__59128),
            .I(N__59119));
    LocalMux I__11988 (
            .O(N__59125),
            .I(N__59116));
    InMux I__11987 (
            .O(N__59122),
            .I(N__59113));
    InMux I__11986 (
            .O(N__59119),
            .I(N__59110));
    Span4Mux_v I__11985 (
            .O(N__59116),
            .I(N__59107));
    LocalMux I__11984 (
            .O(N__59113),
            .I(N__59104));
    LocalMux I__11983 (
            .O(N__59110),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    Odrv4 I__11982 (
            .O(N__59107),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    Odrv12 I__11981 (
            .O(N__59104),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__11980 (
            .O(N__59097),
            .I(N__59094));
    LocalMux I__11979 (
            .O(N__59094),
            .I(N__59091));
    Span4Mux_v I__11978 (
            .O(N__59091),
            .I(N__59088));
    Odrv4 I__11977 (
            .O(N__59088),
            .I(\ppm_encoder_1.N_290 ));
    InMux I__11976 (
            .O(N__59085),
            .I(N__59079));
    InMux I__11975 (
            .O(N__59084),
            .I(N__59074));
    InMux I__11974 (
            .O(N__59083),
            .I(N__59074));
    InMux I__11973 (
            .O(N__59082),
            .I(N__59071));
    LocalMux I__11972 (
            .O(N__59079),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__11971 (
            .O(N__59074),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__11970 (
            .O(N__59071),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    InMux I__11969 (
            .O(N__59064),
            .I(N__59060));
    InMux I__11968 (
            .O(N__59063),
            .I(N__59057));
    LocalMux I__11967 (
            .O(N__59060),
            .I(N__59053));
    LocalMux I__11966 (
            .O(N__59057),
            .I(N__59050));
    InMux I__11965 (
            .O(N__59056),
            .I(N__59047));
    Span4Mux_h I__11964 (
            .O(N__59053),
            .I(N__59044));
    Span4Mux_h I__11963 (
            .O(N__59050),
            .I(N__59041));
    LocalMux I__11962 (
            .O(N__59047),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__11961 (
            .O(N__59044),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__11960 (
            .O(N__59041),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    CascadeMux I__11959 (
            .O(N__59034),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGAZ0Z_0_cascade_ ));
    CascadeMux I__11958 (
            .O(N__59031),
            .I(\ppm_encoder_1.throttle_m_1_cascade_ ));
    InMux I__11957 (
            .O(N__59028),
            .I(N__59025));
    LocalMux I__11956 (
            .O(N__59025),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1 ));
    InMux I__11955 (
            .O(N__59022),
            .I(N__59018));
    InMux I__11954 (
            .O(N__59021),
            .I(N__59015));
    LocalMux I__11953 (
            .O(N__59018),
            .I(\pid_front.N_110 ));
    LocalMux I__11952 (
            .O(N__59015),
            .I(\pid_front.N_110 ));
    CascadeMux I__11951 (
            .O(N__59010),
            .I(N__59007));
    InMux I__11950 (
            .O(N__59007),
            .I(N__59004));
    LocalMux I__11949 (
            .O(N__59004),
            .I(N__59001));
    Span4Mux_v I__11948 (
            .O(N__59001),
            .I(N__58998));
    Span4Mux_h I__11947 (
            .O(N__58998),
            .I(N__58995));
    Odrv4 I__11946 (
            .O(N__58995),
            .I(\pid_front.error_i_regZ0Z_6 ));
    InMux I__11945 (
            .O(N__58992),
            .I(N__58989));
    LocalMux I__11944 (
            .O(N__58989),
            .I(N__58983));
    InMux I__11943 (
            .O(N__58988),
            .I(N__58980));
    InMux I__11942 (
            .O(N__58987),
            .I(N__58975));
    InMux I__11941 (
            .O(N__58986),
            .I(N__58975));
    Span4Mux_h I__11940 (
            .O(N__58983),
            .I(N__58970));
    LocalMux I__11939 (
            .O(N__58980),
            .I(N__58970));
    LocalMux I__11938 (
            .O(N__58975),
            .I(\pid_front.N_15_0 ));
    Odrv4 I__11937 (
            .O(N__58970),
            .I(\pid_front.N_15_0 ));
    InMux I__11936 (
            .O(N__58965),
            .I(N__58962));
    LocalMux I__11935 (
            .O(N__58962),
            .I(N__58959));
    Odrv4 I__11934 (
            .O(N__58959),
            .I(\pid_front.N_32_0 ));
    CascadeMux I__11933 (
            .O(N__58956),
            .I(\pid_front.N_32_0_cascade_ ));
    InMux I__11932 (
            .O(N__58953),
            .I(N__58950));
    LocalMux I__11931 (
            .O(N__58950),
            .I(N__58946));
    InMux I__11930 (
            .O(N__58949),
            .I(N__58943));
    Odrv4 I__11929 (
            .O(N__58946),
            .I(\pid_front.N_29_1 ));
    LocalMux I__11928 (
            .O(N__58943),
            .I(\pid_front.N_29_1 ));
    CascadeMux I__11927 (
            .O(N__58938),
            .I(N__58935));
    InMux I__11926 (
            .O(N__58935),
            .I(N__58932));
    LocalMux I__11925 (
            .O(N__58932),
            .I(N__58929));
    Span4Mux_v I__11924 (
            .O(N__58929),
            .I(N__58926));
    Span4Mux_h I__11923 (
            .O(N__58926),
            .I(N__58923));
    Odrv4 I__11922 (
            .O(N__58923),
            .I(\pid_front.error_i_regZ0Z_8 ));
    InMux I__11921 (
            .O(N__58920),
            .I(N__58917));
    LocalMux I__11920 (
            .O(N__58917),
            .I(N__58914));
    Span12Mux_s6_v I__11919 (
            .O(N__58914),
            .I(N__58908));
    InMux I__11918 (
            .O(N__58913),
            .I(N__58903));
    InMux I__11917 (
            .O(N__58912),
            .I(N__58903));
    InMux I__11916 (
            .O(N__58911),
            .I(N__58900));
    Odrv12 I__11915 (
            .O(N__58908),
            .I(\pid_front.m1_0_03 ));
    LocalMux I__11914 (
            .O(N__58903),
            .I(\pid_front.m1_0_03 ));
    LocalMux I__11913 (
            .O(N__58900),
            .I(\pid_front.m1_0_03 ));
    CascadeMux I__11912 (
            .O(N__58893),
            .I(\pid_front.N_117_cascade_ ));
    InMux I__11911 (
            .O(N__58890),
            .I(N__58887));
    LocalMux I__11910 (
            .O(N__58887),
            .I(N__58884));
    Odrv12 I__11909 (
            .O(N__58884),
            .I(\pid_front.N_116_0 ));
    InMux I__11908 (
            .O(N__58881),
            .I(N__58876));
    InMux I__11907 (
            .O(N__58880),
            .I(N__58871));
    InMux I__11906 (
            .O(N__58879),
            .I(N__58871));
    LocalMux I__11905 (
            .O(N__58876),
            .I(\pid_side.N_15_1 ));
    LocalMux I__11904 (
            .O(N__58871),
            .I(\pid_side.N_15_1 ));
    InMux I__11903 (
            .O(N__58866),
            .I(N__58860));
    InMux I__11902 (
            .O(N__58865),
            .I(N__58857));
    InMux I__11901 (
            .O(N__58864),
            .I(N__58852));
    InMux I__11900 (
            .O(N__58863),
            .I(N__58852));
    LocalMux I__11899 (
            .O(N__58860),
            .I(\pid_side.N_39_0 ));
    LocalMux I__11898 (
            .O(N__58857),
            .I(\pid_side.N_39_0 ));
    LocalMux I__11897 (
            .O(N__58852),
            .I(\pid_side.N_39_0 ));
    CascadeMux I__11896 (
            .O(N__58845),
            .I(N__58842));
    InMux I__11895 (
            .O(N__58842),
            .I(N__58839));
    LocalMux I__11894 (
            .O(N__58839),
            .I(N__58836));
    Odrv12 I__11893 (
            .O(N__58836),
            .I(\pid_side.error_i_regZ0Z_3 ));
    CascadeMux I__11892 (
            .O(N__58833),
            .I(\pid_side.m5_2_03_cascade_ ));
    InMux I__11891 (
            .O(N__58830),
            .I(N__58827));
    LocalMux I__11890 (
            .O(N__58827),
            .I(N__58824));
    Odrv12 I__11889 (
            .O(N__58824),
            .I(\pid_side.error_i_regZ0Z_17 ));
    InMux I__11888 (
            .O(N__58821),
            .I(N__58818));
    LocalMux I__11887 (
            .O(N__58818),
            .I(N__58815));
    Odrv12 I__11886 (
            .O(N__58815),
            .I(\pid_side.m27_2_03_0 ));
    InMux I__11885 (
            .O(N__58812),
            .I(N__58809));
    LocalMux I__11884 (
            .O(N__58809),
            .I(\pid_side.m11_2_03_3_i_0 ));
    InMux I__11883 (
            .O(N__58806),
            .I(N__58803));
    LocalMux I__11882 (
            .O(N__58803),
            .I(N__58800));
    Span12Mux_s10_h I__11881 (
            .O(N__58800),
            .I(N__58797));
    Odrv12 I__11880 (
            .O(N__58797),
            .I(\pid_side.error_i_regZ0Z_23 ));
    InMux I__11879 (
            .O(N__58794),
            .I(N__58791));
    LocalMux I__11878 (
            .O(N__58791),
            .I(N__58788));
    Span4Mux_v I__11877 (
            .O(N__58788),
            .I(N__58785));
    Odrv4 I__11876 (
            .O(N__58785),
            .I(\pid_side.error_i_regZ0Z_24 ));
    InMux I__11875 (
            .O(N__58782),
            .I(N__58779));
    LocalMux I__11874 (
            .O(N__58779),
            .I(\pid_side.m136_ns_1 ));
    CascadeMux I__11873 (
            .O(N__58776),
            .I(\pid_side.N_110_cascade_ ));
    InMux I__11872 (
            .O(N__58773),
            .I(N__58769));
    InMux I__11871 (
            .O(N__58772),
            .I(N__58764));
    LocalMux I__11870 (
            .O(N__58769),
            .I(N__58761));
    InMux I__11869 (
            .O(N__58768),
            .I(N__58756));
    InMux I__11868 (
            .O(N__58767),
            .I(N__58756));
    LocalMux I__11867 (
            .O(N__58764),
            .I(N__58748));
    Span4Mux_v I__11866 (
            .O(N__58761),
            .I(N__58748));
    LocalMux I__11865 (
            .O(N__58756),
            .I(N__58748));
    InMux I__11864 (
            .O(N__58755),
            .I(N__58745));
    Odrv4 I__11863 (
            .O(N__58748),
            .I(\pid_side.m2_0_03_3_i_0 ));
    LocalMux I__11862 (
            .O(N__58745),
            .I(\pid_side.m2_0_03_3_i_0 ));
    InMux I__11861 (
            .O(N__58740),
            .I(N__58737));
    LocalMux I__11860 (
            .O(N__58737),
            .I(\pid_side.m7_2_03 ));
    InMux I__11859 (
            .O(N__58734),
            .I(N__58731));
    LocalMux I__11858 (
            .O(N__58731),
            .I(N__58728));
    Odrv4 I__11857 (
            .O(N__58728),
            .I(\pid_side.error_i_reg_9_rn_0_19 ));
    InMux I__11856 (
            .O(N__58725),
            .I(N__58722));
    LocalMux I__11855 (
            .O(N__58722),
            .I(N__58719));
    Odrv4 I__11854 (
            .O(N__58719),
            .I(\pid_side.N_53_0 ));
    CascadeMux I__11853 (
            .O(N__58716),
            .I(\pid_side.N_53_0_cascade_ ));
    InMux I__11852 (
            .O(N__58713),
            .I(N__58710));
    LocalMux I__11851 (
            .O(N__58710),
            .I(N__58707));
    Odrv4 I__11850 (
            .O(N__58707),
            .I(\pid_side.error_i_reg_9_rn_0_27 ));
    InMux I__11849 (
            .O(N__58704),
            .I(N__58701));
    LocalMux I__11848 (
            .O(N__58701),
            .I(\pid_side.error_cry_0_c_RNI9I2AZ0Z2 ));
    InMux I__11847 (
            .O(N__58698),
            .I(N__58695));
    LocalMux I__11846 (
            .O(N__58695),
            .I(N__58692));
    Span4Mux_h I__11845 (
            .O(N__58692),
            .I(N__58689));
    Odrv4 I__11844 (
            .O(N__58689),
            .I(\pid_side.m104_ns_sx ));
    CascadeMux I__11843 (
            .O(N__58686),
            .I(\pid_side.m104_ns_sx_cascade_ ));
    CascadeMux I__11842 (
            .O(N__58683),
            .I(N__58680));
    InMux I__11841 (
            .O(N__58680),
            .I(N__58675));
    InMux I__11840 (
            .O(N__58679),
            .I(N__58672));
    InMux I__11839 (
            .O(N__58678),
            .I(N__58669));
    LocalMux I__11838 (
            .O(N__58675),
            .I(N__58666));
    LocalMux I__11837 (
            .O(N__58672),
            .I(\pid_side.N_49_0 ));
    LocalMux I__11836 (
            .O(N__58669),
            .I(\pid_side.N_49_0 ));
    Odrv4 I__11835 (
            .O(N__58666),
            .I(\pid_side.N_49_0 ));
    InMux I__11834 (
            .O(N__58659),
            .I(N__58655));
    CascadeMux I__11833 (
            .O(N__58658),
            .I(N__58652));
    LocalMux I__11832 (
            .O(N__58655),
            .I(N__58649));
    InMux I__11831 (
            .O(N__58652),
            .I(N__58646));
    Span4Mux_v I__11830 (
            .O(N__58649),
            .I(N__58643));
    LocalMux I__11829 (
            .O(N__58646),
            .I(N__58640));
    Odrv4 I__11828 (
            .O(N__58643),
            .I(\pid_side.error_i_regZ0Z_0 ));
    Odrv12 I__11827 (
            .O(N__58640),
            .I(\pid_side.error_i_regZ0Z_0 ));
    CascadeMux I__11826 (
            .O(N__58635),
            .I(N__58632));
    InMux I__11825 (
            .O(N__58632),
            .I(N__58629));
    LocalMux I__11824 (
            .O(N__58629),
            .I(N__58626));
    Odrv12 I__11823 (
            .O(N__58626),
            .I(\pid_side.error_i_regZ0Z_1 ));
    CascadeMux I__11822 (
            .O(N__58623),
            .I(N__58620));
    InMux I__11821 (
            .O(N__58620),
            .I(N__58617));
    LocalMux I__11820 (
            .O(N__58617),
            .I(N__58614));
    Odrv12 I__11819 (
            .O(N__58614),
            .I(\pid_side.error_i_regZ0Z_2 ));
    InMux I__11818 (
            .O(N__58611),
            .I(N__58605));
    InMux I__11817 (
            .O(N__58610),
            .I(N__58605));
    LocalMux I__11816 (
            .O(N__58605),
            .I(\pid_side.N_50_1 ));
    InMux I__11815 (
            .O(N__58602),
            .I(N__58599));
    LocalMux I__11814 (
            .O(N__58599),
            .I(N__58596));
    Odrv12 I__11813 (
            .O(N__58596),
            .I(\pid_side.error_i_regZ0Z_19 ));
    CascadeMux I__11812 (
            .O(N__58593),
            .I(N__58590));
    InMux I__11811 (
            .O(N__58590),
            .I(N__58587));
    LocalMux I__11810 (
            .O(N__58587),
            .I(N__58584));
    Odrv12 I__11809 (
            .O(N__58584),
            .I(\pid_side.error_i_regZ0Z_18 ));
    CascadeMux I__11808 (
            .O(N__58581),
            .I(\pid_side.N_3_cascade_ ));
    CascadeMux I__11807 (
            .O(N__58578),
            .I(\pid_side.m2_0_03_3_i_0_cascade_ ));
    CascadeMux I__11806 (
            .O(N__58575),
            .I(\pid_side.m6_2_03_cascade_ ));
    InMux I__11805 (
            .O(N__58572),
            .I(N__58569));
    LocalMux I__11804 (
            .O(N__58569),
            .I(\pid_side.error_i_reg_9_rn_0_18 ));
    CascadeMux I__11803 (
            .O(N__58566),
            .I(\pid_side.m51_0_ns_1_cascade_ ));
    CascadeMux I__11802 (
            .O(N__58563),
            .I(\pid_side.N_39_0_cascade_ ));
    InMux I__11801 (
            .O(N__58560),
            .I(N__58554));
    InMux I__11800 (
            .O(N__58559),
            .I(N__58554));
    LocalMux I__11799 (
            .O(N__58554),
            .I(\dron_frame_decoder_1.drone_H_disp_side_4 ));
    SRMux I__11798 (
            .O(N__58551),
            .I(N__58547));
    SRMux I__11797 (
            .O(N__58550),
            .I(N__58544));
    LocalMux I__11796 (
            .O(N__58547),
            .I(N__58541));
    LocalMux I__11795 (
            .O(N__58544),
            .I(N__58538));
    Span4Mux_v I__11794 (
            .O(N__58541),
            .I(N__58535));
    Span4Mux_v I__11793 (
            .O(N__58538),
            .I(N__58532));
    Span4Mux_h I__11792 (
            .O(N__58535),
            .I(N__58529));
    Span4Mux_v I__11791 (
            .O(N__58532),
            .I(N__58526));
    Span4Mux_v I__11790 (
            .O(N__58529),
            .I(N__58521));
    Span4Mux_h I__11789 (
            .O(N__58526),
            .I(N__58521));
    Odrv4 I__11788 (
            .O(N__58521),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    CascadeMux I__11787 (
            .O(N__58518),
            .I(N__58514));
    InMux I__11786 (
            .O(N__58517),
            .I(N__58499));
    InMux I__11785 (
            .O(N__58514),
            .I(N__58499));
    InMux I__11784 (
            .O(N__58513),
            .I(N__58496));
    CascadeMux I__11783 (
            .O(N__58512),
            .I(N__58492));
    CascadeMux I__11782 (
            .O(N__58511),
            .I(N__58489));
    CascadeMux I__11781 (
            .O(N__58510),
            .I(N__58486));
    CascadeMux I__11780 (
            .O(N__58509),
            .I(N__58480));
    CascadeMux I__11779 (
            .O(N__58508),
            .I(N__58477));
    CascadeMux I__11778 (
            .O(N__58507),
            .I(N__58474));
    CascadeMux I__11777 (
            .O(N__58506),
            .I(N__58471));
    CascadeMux I__11776 (
            .O(N__58505),
            .I(N__58467));
    CascadeMux I__11775 (
            .O(N__58504),
            .I(N__58464));
    LocalMux I__11774 (
            .O(N__58499),
            .I(N__58461));
    LocalMux I__11773 (
            .O(N__58496),
            .I(N__58458));
    InMux I__11772 (
            .O(N__58495),
            .I(N__58449));
    InMux I__11771 (
            .O(N__58492),
            .I(N__58449));
    InMux I__11770 (
            .O(N__58489),
            .I(N__58449));
    InMux I__11769 (
            .O(N__58486),
            .I(N__58449));
    CascadeMux I__11768 (
            .O(N__58485),
            .I(N__58446));
    CascadeMux I__11767 (
            .O(N__58484),
            .I(N__58443));
    InMux I__11766 (
            .O(N__58483),
            .I(N__58434));
    InMux I__11765 (
            .O(N__58480),
            .I(N__58434));
    InMux I__11764 (
            .O(N__58477),
            .I(N__58434));
    InMux I__11763 (
            .O(N__58474),
            .I(N__58434));
    InMux I__11762 (
            .O(N__58471),
            .I(N__58425));
    InMux I__11761 (
            .O(N__58470),
            .I(N__58425));
    InMux I__11760 (
            .O(N__58467),
            .I(N__58425));
    InMux I__11759 (
            .O(N__58464),
            .I(N__58425));
    Span4Mux_h I__11758 (
            .O(N__58461),
            .I(N__58422));
    Span4Mux_h I__11757 (
            .O(N__58458),
            .I(N__58419));
    LocalMux I__11756 (
            .O(N__58449),
            .I(N__58416));
    InMux I__11755 (
            .O(N__58446),
            .I(N__58411));
    InMux I__11754 (
            .O(N__58443),
            .I(N__58411));
    LocalMux I__11753 (
            .O(N__58434),
            .I(N__58405));
    LocalMux I__11752 (
            .O(N__58425),
            .I(N__58405));
    Span4Mux_v I__11751 (
            .O(N__58422),
            .I(N__58402));
    Span4Mux_v I__11750 (
            .O(N__58419),
            .I(N__58398));
    Span4Mux_h I__11749 (
            .O(N__58416),
            .I(N__58393));
    LocalMux I__11748 (
            .O(N__58411),
            .I(N__58393));
    InMux I__11747 (
            .O(N__58410),
            .I(N__58390));
    Span4Mux_v I__11746 (
            .O(N__58405),
            .I(N__58386));
    Sp12to4 I__11745 (
            .O(N__58402),
            .I(N__58383));
    InMux I__11744 (
            .O(N__58401),
            .I(N__58380));
    Span4Mux_h I__11743 (
            .O(N__58398),
            .I(N__58373));
    Span4Mux_v I__11742 (
            .O(N__58393),
            .I(N__58373));
    LocalMux I__11741 (
            .O(N__58390),
            .I(N__58373));
    InMux I__11740 (
            .O(N__58389),
            .I(N__58370));
    Span4Mux_h I__11739 (
            .O(N__58386),
            .I(N__58367));
    Span12Mux_h I__11738 (
            .O(N__58383),
            .I(N__58362));
    LocalMux I__11737 (
            .O(N__58380),
            .I(N__58362));
    Span4Mux_h I__11736 (
            .O(N__58373),
            .I(N__58359));
    LocalMux I__11735 (
            .O(N__58370),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__11734 (
            .O(N__58367),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv12 I__11733 (
            .O(N__58362),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__11732 (
            .O(N__58359),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    InMux I__11731 (
            .O(N__58350),
            .I(N__58343));
    InMux I__11730 (
            .O(N__58349),
            .I(N__58335));
    InMux I__11729 (
            .O(N__58348),
            .I(N__58328));
    InMux I__11728 (
            .O(N__58347),
            .I(N__58328));
    InMux I__11727 (
            .O(N__58346),
            .I(N__58328));
    LocalMux I__11726 (
            .O(N__58343),
            .I(N__58325));
    InMux I__11725 (
            .O(N__58342),
            .I(N__58322));
    InMux I__11724 (
            .O(N__58341),
            .I(N__58313));
    InMux I__11723 (
            .O(N__58340),
            .I(N__58313));
    InMux I__11722 (
            .O(N__58339),
            .I(N__58313));
    InMux I__11721 (
            .O(N__58338),
            .I(N__58313));
    LocalMux I__11720 (
            .O(N__58335),
            .I(N__58306));
    LocalMux I__11719 (
            .O(N__58328),
            .I(N__58306));
    Span4Mux_v I__11718 (
            .O(N__58325),
            .I(N__58298));
    LocalMux I__11717 (
            .O(N__58322),
            .I(N__58295));
    LocalMux I__11716 (
            .O(N__58313),
            .I(N__58292));
    InMux I__11715 (
            .O(N__58312),
            .I(N__58287));
    InMux I__11714 (
            .O(N__58311),
            .I(N__58287));
    Span4Mux_h I__11713 (
            .O(N__58306),
            .I(N__58284));
    InMux I__11712 (
            .O(N__58305),
            .I(N__58281));
    InMux I__11711 (
            .O(N__58304),
            .I(N__58277));
    CascadeMux I__11710 (
            .O(N__58303),
            .I(N__58273));
    CascadeMux I__11709 (
            .O(N__58302),
            .I(N__58270));
    CascadeMux I__11708 (
            .O(N__58301),
            .I(N__58266));
    Span4Mux_h I__11707 (
            .O(N__58298),
            .I(N__58261));
    Span4Mux_h I__11706 (
            .O(N__58295),
            .I(N__58252));
    Span4Mux_v I__11705 (
            .O(N__58292),
            .I(N__58252));
    LocalMux I__11704 (
            .O(N__58287),
            .I(N__58252));
    Span4Mux_h I__11703 (
            .O(N__58284),
            .I(N__58252));
    LocalMux I__11702 (
            .O(N__58281),
            .I(N__58249));
    CascadeMux I__11701 (
            .O(N__58280),
            .I(N__58246));
    LocalMux I__11700 (
            .O(N__58277),
            .I(N__58243));
    InMux I__11699 (
            .O(N__58276),
            .I(N__58228));
    InMux I__11698 (
            .O(N__58273),
            .I(N__58228));
    InMux I__11697 (
            .O(N__58270),
            .I(N__58228));
    InMux I__11696 (
            .O(N__58269),
            .I(N__58228));
    InMux I__11695 (
            .O(N__58266),
            .I(N__58228));
    InMux I__11694 (
            .O(N__58265),
            .I(N__58228));
    InMux I__11693 (
            .O(N__58264),
            .I(N__58228));
    Span4Mux_v I__11692 (
            .O(N__58261),
            .I(N__58225));
    Span4Mux_v I__11691 (
            .O(N__58252),
            .I(N__58220));
    Span4Mux_h I__11690 (
            .O(N__58249),
            .I(N__58220));
    InMux I__11689 (
            .O(N__58246),
            .I(N__58217));
    Odrv12 I__11688 (
            .O(N__58243),
            .I(uart_drone_data_rdy));
    LocalMux I__11687 (
            .O(N__58228),
            .I(uart_drone_data_rdy));
    Odrv4 I__11686 (
            .O(N__58225),
            .I(uart_drone_data_rdy));
    Odrv4 I__11685 (
            .O(N__58220),
            .I(uart_drone_data_rdy));
    LocalMux I__11684 (
            .O(N__58217),
            .I(uart_drone_data_rdy));
    CascadeMux I__11683 (
            .O(N__58206),
            .I(\pid_side.m45_0_ns_1_cascade_ ));
    CascadeMux I__11682 (
            .O(N__58203),
            .I(\pid_side.N_46_1_cascade_ ));
    InMux I__11681 (
            .O(N__58200),
            .I(N__58197));
    LocalMux I__11680 (
            .O(N__58197),
            .I(N__58194));
    Span4Mux_h I__11679 (
            .O(N__58194),
            .I(N__58190));
    InMux I__11678 (
            .O(N__58193),
            .I(N__58187));
    Odrv4 I__11677 (
            .O(N__58190),
            .I(\pid_side.N_46_1 ));
    LocalMux I__11676 (
            .O(N__58187),
            .I(\pid_side.N_46_1 ));
    CascadeMux I__11675 (
            .O(N__58182),
            .I(\pid_side.N_50_1_cascade_ ));
    CascadeMux I__11674 (
            .O(N__58179),
            .I(N__58176));
    InMux I__11673 (
            .O(N__58176),
            .I(N__58173));
    LocalMux I__11672 (
            .O(N__58173),
            .I(N__58170));
    Odrv12 I__11671 (
            .O(N__58170),
            .I(\pid_side.error_i_regZ0Z_11 ));
    CascadeMux I__11670 (
            .O(N__58167),
            .I(N__58163));
    InMux I__11669 (
            .O(N__58166),
            .I(N__58158));
    InMux I__11668 (
            .O(N__58163),
            .I(N__58158));
    LocalMux I__11667 (
            .O(N__58158),
            .I(N__58155));
    Odrv4 I__11666 (
            .O(N__58155),
            .I(\pid_side.error_i_regZ0Z_27 ));
    InMux I__11665 (
            .O(N__58152),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26 ));
    CascadeMux I__11664 (
            .O(N__58149),
            .I(N__58143));
    CascadeMux I__11663 (
            .O(N__58148),
            .I(N__58139));
    InMux I__11662 (
            .O(N__58147),
            .I(N__58123));
    InMux I__11661 (
            .O(N__58146),
            .I(N__58123));
    InMux I__11660 (
            .O(N__58143),
            .I(N__58123));
    InMux I__11659 (
            .O(N__58142),
            .I(N__58123));
    InMux I__11658 (
            .O(N__58139),
            .I(N__58123));
    CascadeMux I__11657 (
            .O(N__58138),
            .I(N__58120));
    CascadeMux I__11656 (
            .O(N__58137),
            .I(N__58116));
    CascadeMux I__11655 (
            .O(N__58136),
            .I(N__58112));
    CascadeMux I__11654 (
            .O(N__58135),
            .I(N__58108));
    CascadeMux I__11653 (
            .O(N__58134),
            .I(N__58103));
    LocalMux I__11652 (
            .O(N__58123),
            .I(N__58099));
    InMux I__11651 (
            .O(N__58120),
            .I(N__58082));
    InMux I__11650 (
            .O(N__58119),
            .I(N__58082));
    InMux I__11649 (
            .O(N__58116),
            .I(N__58082));
    InMux I__11648 (
            .O(N__58115),
            .I(N__58082));
    InMux I__11647 (
            .O(N__58112),
            .I(N__58082));
    InMux I__11646 (
            .O(N__58111),
            .I(N__58082));
    InMux I__11645 (
            .O(N__58108),
            .I(N__58082));
    InMux I__11644 (
            .O(N__58107),
            .I(N__58082));
    InMux I__11643 (
            .O(N__58106),
            .I(N__58075));
    InMux I__11642 (
            .O(N__58103),
            .I(N__58075));
    InMux I__11641 (
            .O(N__58102),
            .I(N__58075));
    Odrv4 I__11640 (
            .O(N__58099),
            .I(\pid_side.error_i_acummZ0Z_13 ));
    LocalMux I__11639 (
            .O(N__58082),
            .I(\pid_side.error_i_acummZ0Z_13 ));
    LocalMux I__11638 (
            .O(N__58075),
            .I(\pid_side.error_i_acummZ0Z_13 ));
    InMux I__11637 (
            .O(N__58068),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__11636 (
            .O(N__58065),
            .I(N__58059));
    InMux I__11635 (
            .O(N__58064),
            .I(N__58059));
    LocalMux I__11634 (
            .O(N__58059),
            .I(\pid_side.error_i_acumm_preregZ0Z_27 ));
    CascadeMux I__11633 (
            .O(N__58056),
            .I(N__58052));
    InMux I__11632 (
            .O(N__58055),
            .I(N__58047));
    InMux I__11631 (
            .O(N__58052),
            .I(N__58047));
    LocalMux I__11630 (
            .O(N__58047),
            .I(\pid_side.error_i_acumm_preregZ0Z_25 ));
    InMux I__11629 (
            .O(N__58044),
            .I(N__58041));
    LocalMux I__11628 (
            .O(N__58041),
            .I(N__58038));
    Span4Mux_h I__11627 (
            .O(N__58038),
            .I(N__58033));
    InMux I__11626 (
            .O(N__58037),
            .I(N__58030));
    CascadeMux I__11625 (
            .O(N__58036),
            .I(N__58026));
    Span4Mux_h I__11624 (
            .O(N__58033),
            .I(N__58023));
    LocalMux I__11623 (
            .O(N__58030),
            .I(N__58020));
    InMux I__11622 (
            .O(N__58029),
            .I(N__58015));
    InMux I__11621 (
            .O(N__58026),
            .I(N__58015));
    Span4Mux_v I__11620 (
            .O(N__58023),
            .I(N__58010));
    Span4Mux_v I__11619 (
            .O(N__58020),
            .I(N__58010));
    LocalMux I__11618 (
            .O(N__58015),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    Odrv4 I__11617 (
            .O(N__58010),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    InMux I__11616 (
            .O(N__58005),
            .I(N__58001));
    InMux I__11615 (
            .O(N__58004),
            .I(N__57998));
    LocalMux I__11614 (
            .O(N__58001),
            .I(N__57992));
    LocalMux I__11613 (
            .O(N__57998),
            .I(N__57988));
    InMux I__11612 (
            .O(N__57997),
            .I(N__57985));
    InMux I__11611 (
            .O(N__57996),
            .I(N__57980));
    InMux I__11610 (
            .O(N__57995),
            .I(N__57980));
    Span4Mux_v I__11609 (
            .O(N__57992),
            .I(N__57975));
    InMux I__11608 (
            .O(N__57991),
            .I(N__57972));
    Span4Mux_h I__11607 (
            .O(N__57988),
            .I(N__57969));
    LocalMux I__11606 (
            .O(N__57985),
            .I(N__57964));
    LocalMux I__11605 (
            .O(N__57980),
            .I(N__57964));
    InMux I__11604 (
            .O(N__57979),
            .I(N__57959));
    InMux I__11603 (
            .O(N__57978),
            .I(N__57959));
    Span4Mux_h I__11602 (
            .O(N__57975),
            .I(N__57956));
    LocalMux I__11601 (
            .O(N__57972),
            .I(N__57953));
    Sp12to4 I__11600 (
            .O(N__57969),
            .I(N__57948));
    Sp12to4 I__11599 (
            .O(N__57964),
            .I(N__57948));
    LocalMux I__11598 (
            .O(N__57959),
            .I(N__57945));
    Span4Mux_v I__11597 (
            .O(N__57956),
            .I(N__57940));
    Span4Mux_v I__11596 (
            .O(N__57953),
            .I(N__57940));
    Span12Mux_v I__11595 (
            .O(N__57948),
            .I(N__57937));
    Span4Mux_h I__11594 (
            .O(N__57945),
            .I(N__57934));
    Odrv4 I__11593 (
            .O(N__57940),
            .I(uart_drone_data_1));
    Odrv12 I__11592 (
            .O(N__57937),
            .I(uart_drone_data_1));
    Odrv4 I__11591 (
            .O(N__57934),
            .I(uart_drone_data_1));
    CascadeMux I__11590 (
            .O(N__57927),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_1_0_cascade_ ));
    InMux I__11589 (
            .O(N__57924),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__11588 (
            .O(N__57921),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__11587 (
            .O(N__57918),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__11586 (
            .O(N__57915),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__11585 (
            .O(N__57912),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__11584 (
            .O(N__57909),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_22 ));
    InMux I__11583 (
            .O(N__57906),
            .I(bfn_15_18_0_));
    InMux I__11582 (
            .O(N__57903),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_24 ));
    InMux I__11581 (
            .O(N__57900),
            .I(N__57897));
    LocalMux I__11580 (
            .O(N__57897),
            .I(N__57894));
    Odrv4 I__11579 (
            .O(N__57894),
            .I(\pid_side.error_i_regZ0Z_26 ));
    InMux I__11578 (
            .O(N__57891),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_25 ));
    InMux I__11577 (
            .O(N__57888),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__11576 (
            .O(N__57885),
            .I(N__57882));
    LocalMux I__11575 (
            .O(N__57882),
            .I(\pid_side.error_i_acummZ0Z_10 ));
    InMux I__11574 (
            .O(N__57879),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__11573 (
            .O(N__57876),
            .I(N__57873));
    LocalMux I__11572 (
            .O(N__57873),
            .I(\pid_side.error_i_acummZ0Z_11 ));
    InMux I__11571 (
            .O(N__57870),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__11570 (
            .O(N__57867),
            .I(N__57864));
    LocalMux I__11569 (
            .O(N__57864),
            .I(N__57861));
    Span4Mux_v I__11568 (
            .O(N__57861),
            .I(N__57858));
    Odrv4 I__11567 (
            .O(N__57858),
            .I(\pid_side.error_i_acummZ0Z_12 ));
    InMux I__11566 (
            .O(N__57855),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_11 ));
    CascadeMux I__11565 (
            .O(N__57852),
            .I(N__57849));
    InMux I__11564 (
            .O(N__57849),
            .I(N__57846));
    LocalMux I__11563 (
            .O(N__57846),
            .I(N__57843));
    Span4Mux_h I__11562 (
            .O(N__57843),
            .I(N__57840));
    Odrv4 I__11561 (
            .O(N__57840),
            .I(\pid_side.error_i_regZ0Z_13 ));
    InMux I__11560 (
            .O(N__57837),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__11559 (
            .O(N__57834),
            .I(N__57831));
    LocalMux I__11558 (
            .O(N__57831),
            .I(N__57828));
    Span4Mux_v I__11557 (
            .O(N__57828),
            .I(N__57825));
    Span4Mux_v I__11556 (
            .O(N__57825),
            .I(N__57822));
    Odrv4 I__11555 (
            .O(N__57822),
            .I(\pid_side.error_i_regZ0Z_14 ));
    InMux I__11554 (
            .O(N__57819),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_13 ));
    CascadeMux I__11553 (
            .O(N__57816),
            .I(N__57813));
    InMux I__11552 (
            .O(N__57813),
            .I(N__57810));
    LocalMux I__11551 (
            .O(N__57810),
            .I(N__57807));
    Span4Mux_h I__11550 (
            .O(N__57807),
            .I(N__57804));
    Span4Mux_v I__11549 (
            .O(N__57804),
            .I(N__57801));
    Odrv4 I__11548 (
            .O(N__57801),
            .I(\pid_side.error_i_regZ0Z_15 ));
    InMux I__11547 (
            .O(N__57798),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__11546 (
            .O(N__57795),
            .I(bfn_15_17_0_));
    InMux I__11545 (
            .O(N__57792),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__11544 (
            .O(N__57789),
            .I(N__57786));
    LocalMux I__11543 (
            .O(N__57786),
            .I(\pid_side.error_i_acummZ0Z_1 ));
    InMux I__11542 (
            .O(N__57783),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__11541 (
            .O(N__57780),
            .I(N__57777));
    LocalMux I__11540 (
            .O(N__57777),
            .I(\pid_side.error_i_acummZ0Z_2 ));
    InMux I__11539 (
            .O(N__57774),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__11538 (
            .O(N__57771),
            .I(N__57768));
    LocalMux I__11537 (
            .O(N__57768),
            .I(\pid_side.error_i_acummZ0Z_3 ));
    InMux I__11536 (
            .O(N__57765),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__11535 (
            .O(N__57762),
            .I(N__57759));
    LocalMux I__11534 (
            .O(N__57759),
            .I(\pid_side.error_i_acummZ0Z_4 ));
    InMux I__11533 (
            .O(N__57756),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__11532 (
            .O(N__57753),
            .I(N__57750));
    LocalMux I__11531 (
            .O(N__57750),
            .I(N__57747));
    Odrv4 I__11530 (
            .O(N__57747),
            .I(\pid_side.error_i_acummZ0Z_5 ));
    InMux I__11529 (
            .O(N__57744),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4 ));
    CascadeMux I__11528 (
            .O(N__57741),
            .I(N__57738));
    InMux I__11527 (
            .O(N__57738),
            .I(N__57735));
    LocalMux I__11526 (
            .O(N__57735),
            .I(\pid_side.error_i_acummZ0Z_6 ));
    InMux I__11525 (
            .O(N__57732),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__11524 (
            .O(N__57729),
            .I(N__57726));
    LocalMux I__11523 (
            .O(N__57726),
            .I(N__57723));
    Span4Mux_v I__11522 (
            .O(N__57723),
            .I(N__57720));
    Odrv4 I__11521 (
            .O(N__57720),
            .I(\pid_side.error_i_regZ0Z_7 ));
    CascadeMux I__11520 (
            .O(N__57717),
            .I(N__57714));
    InMux I__11519 (
            .O(N__57714),
            .I(N__57711));
    LocalMux I__11518 (
            .O(N__57711),
            .I(\pid_side.error_i_acummZ0Z_7 ));
    InMux I__11517 (
            .O(N__57708),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__11516 (
            .O(N__57705),
            .I(N__57702));
    LocalMux I__11515 (
            .O(N__57702),
            .I(N__57699));
    Odrv4 I__11514 (
            .O(N__57699),
            .I(\pid_side.error_i_acummZ0Z_8 ));
    InMux I__11513 (
            .O(N__57696),
            .I(bfn_15_16_0_));
    InMux I__11512 (
            .O(N__57693),
            .I(N__57690));
    LocalMux I__11511 (
            .O(N__57690),
            .I(N__57687));
    Odrv4 I__11510 (
            .O(N__57687),
            .I(\pid_side.error_i_acummZ0Z_9 ));
    InMux I__11509 (
            .O(N__57684),
            .I(N__57681));
    LocalMux I__11508 (
            .O(N__57681),
            .I(N__57677));
    InMux I__11507 (
            .O(N__57680),
            .I(N__57674));
    Span4Mux_v I__11506 (
            .O(N__57677),
            .I(N__57668));
    LocalMux I__11505 (
            .O(N__57674),
            .I(N__57668));
    InMux I__11504 (
            .O(N__57673),
            .I(N__57665));
    Span4Mux_v I__11503 (
            .O(N__57668),
            .I(N__57662));
    LocalMux I__11502 (
            .O(N__57665),
            .I(xy_ki_5));
    Odrv4 I__11501 (
            .O(N__57662),
            .I(xy_ki_5));
    InMux I__11500 (
            .O(N__57657),
            .I(N__57653));
    InMux I__11499 (
            .O(N__57656),
            .I(N__57650));
    LocalMux I__11498 (
            .O(N__57653),
            .I(N__57647));
    LocalMux I__11497 (
            .O(N__57650),
            .I(N__57644));
    Span4Mux_v I__11496 (
            .O(N__57647),
            .I(N__57638));
    Span4Mux_h I__11495 (
            .O(N__57644),
            .I(N__57638));
    InMux I__11494 (
            .O(N__57643),
            .I(N__57635));
    Span4Mux_v I__11493 (
            .O(N__57638),
            .I(N__57632));
    LocalMux I__11492 (
            .O(N__57635),
            .I(xy_ki_6));
    Odrv4 I__11491 (
            .O(N__57632),
            .I(xy_ki_6));
    CascadeMux I__11490 (
            .O(N__57627),
            .I(N__57623));
    InMux I__11489 (
            .O(N__57626),
            .I(N__57620));
    InMux I__11488 (
            .O(N__57623),
            .I(N__57617));
    LocalMux I__11487 (
            .O(N__57620),
            .I(N__57614));
    LocalMux I__11486 (
            .O(N__57617),
            .I(N__57611));
    Span4Mux_v I__11485 (
            .O(N__57614),
            .I(N__57605));
    Span4Mux_h I__11484 (
            .O(N__57611),
            .I(N__57605));
    InMux I__11483 (
            .O(N__57610),
            .I(N__57602));
    Sp12to4 I__11482 (
            .O(N__57605),
            .I(N__57599));
    LocalMux I__11481 (
            .O(N__57602),
            .I(xy_ki_7));
    Odrv12 I__11480 (
            .O(N__57599),
            .I(xy_ki_7));
    InMux I__11479 (
            .O(N__57594),
            .I(N__57590));
    InMux I__11478 (
            .O(N__57593),
            .I(N__57587));
    LocalMux I__11477 (
            .O(N__57590),
            .I(N__57584));
    LocalMux I__11476 (
            .O(N__57587),
            .I(\pid_side.un11lto30_i_a2_5_and ));
    Odrv4 I__11475 (
            .O(N__57584),
            .I(\pid_side.un11lto30_i_a2_5_and ));
    InMux I__11474 (
            .O(N__57579),
            .I(N__57574));
    InMux I__11473 (
            .O(N__57578),
            .I(N__57571));
    InMux I__11472 (
            .O(N__57577),
            .I(N__57568));
    LocalMux I__11471 (
            .O(N__57574),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    LocalMux I__11470 (
            .O(N__57571),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    LocalMux I__11469 (
            .O(N__57568),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    CascadeMux I__11468 (
            .O(N__57561),
            .I(\pid_side.un11lto30_i_a2_5_and_cascade_ ));
    InMux I__11467 (
            .O(N__57558),
            .I(N__57553));
    InMux I__11466 (
            .O(N__57557),
            .I(N__57550));
    InMux I__11465 (
            .O(N__57556),
            .I(N__57547));
    LocalMux I__11464 (
            .O(N__57553),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    LocalMux I__11463 (
            .O(N__57550),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    LocalMux I__11462 (
            .O(N__57547),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    InMux I__11461 (
            .O(N__57540),
            .I(N__57537));
    LocalMux I__11460 (
            .O(N__57537),
            .I(N__57533));
    InMux I__11459 (
            .O(N__57536),
            .I(N__57530));
    Odrv12 I__11458 (
            .O(N__57533),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    LocalMux I__11457 (
            .O(N__57530),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    InMux I__11456 (
            .O(N__57525),
            .I(bfn_15_13_0_));
    InMux I__11455 (
            .O(N__57522),
            .I(N__57519));
    LocalMux I__11454 (
            .O(N__57519),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_o2_sx ));
    InMux I__11453 (
            .O(N__57516),
            .I(N__57513));
    LocalMux I__11452 (
            .O(N__57513),
            .I(\pid_side.N_102 ));
    InMux I__11451 (
            .O(N__57510),
            .I(N__57507));
    LocalMux I__11450 (
            .O(N__57507),
            .I(\pid_side.N_389 ));
    InMux I__11449 (
            .O(N__57504),
            .I(N__57501));
    LocalMux I__11448 (
            .O(N__57501),
            .I(N__57498));
    Span4Mux_h I__11447 (
            .O(N__57498),
            .I(N__57495));
    Span4Mux_h I__11446 (
            .O(N__57495),
            .I(N__57492));
    Odrv4 I__11445 (
            .O(N__57492),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__11444 (
            .O(N__57489),
            .I(\pid_side.pid_prereg_esr_RNIVRQ8Z0Z_20_cascade_ ));
    InMux I__11443 (
            .O(N__57486),
            .I(N__57483));
    LocalMux I__11442 (
            .O(N__57483),
            .I(N__57479));
    InMux I__11441 (
            .O(N__57482),
            .I(N__57476));
    Span4Mux_v I__11440 (
            .O(N__57479),
            .I(N__57473));
    LocalMux I__11439 (
            .O(N__57476),
            .I(N__57470));
    Odrv4 I__11438 (
            .O(N__57473),
            .I(front_order_10));
    Odrv12 I__11437 (
            .O(N__57470),
            .I(front_order_10));
    InMux I__11436 (
            .O(N__57465),
            .I(N__57462));
    LocalMux I__11435 (
            .O(N__57462),
            .I(N__57459));
    Span4Mux_h I__11434 (
            .O(N__57459),
            .I(N__57456));
    Odrv4 I__11433 (
            .O(N__57456),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__11432 (
            .O(N__57453),
            .I(N__57450));
    LocalMux I__11431 (
            .O(N__57450),
            .I(N__57447));
    Odrv4 I__11430 (
            .O(N__57447),
            .I(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ));
    InMux I__11429 (
            .O(N__57444),
            .I(N__57441));
    LocalMux I__11428 (
            .O(N__57441),
            .I(N__57437));
    InMux I__11427 (
            .O(N__57440),
            .I(N__57434));
    Span4Mux_h I__11426 (
            .O(N__57437),
            .I(N__57429));
    LocalMux I__11425 (
            .O(N__57434),
            .I(N__57429));
    Span4Mux_h I__11424 (
            .O(N__57429),
            .I(N__57426));
    Odrv4 I__11423 (
            .O(N__57426),
            .I(front_order_4));
    InMux I__11422 (
            .O(N__57423),
            .I(N__57420));
    LocalMux I__11421 (
            .O(N__57420),
            .I(N__57417));
    Odrv12 I__11420 (
            .O(N__57417),
            .I(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ));
    InMux I__11419 (
            .O(N__57414),
            .I(N__57410));
    InMux I__11418 (
            .O(N__57413),
            .I(N__57407));
    LocalMux I__11417 (
            .O(N__57410),
            .I(N__57404));
    LocalMux I__11416 (
            .O(N__57407),
            .I(N__57401));
    Span4Mux_v I__11415 (
            .O(N__57404),
            .I(N__57398));
    Span4Mux_v I__11414 (
            .O(N__57401),
            .I(N__57395));
    Odrv4 I__11413 (
            .O(N__57398),
            .I(front_order_5));
    Odrv4 I__11412 (
            .O(N__57395),
            .I(front_order_5));
    CascadeMux I__11411 (
            .O(N__57390),
            .I(N__57386));
    InMux I__11410 (
            .O(N__57389),
            .I(N__57380));
    InMux I__11409 (
            .O(N__57386),
            .I(N__57380));
    InMux I__11408 (
            .O(N__57385),
            .I(N__57377));
    LocalMux I__11407 (
            .O(N__57380),
            .I(N__57374));
    LocalMux I__11406 (
            .O(N__57377),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    Odrv12 I__11405 (
            .O(N__57374),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    CascadeMux I__11404 (
            .O(N__57369),
            .I(\ppm_encoder_1.N_299_cascade_ ));
    InMux I__11403 (
            .O(N__57366),
            .I(N__57363));
    LocalMux I__11402 (
            .O(N__57363),
            .I(N__57360));
    Span4Mux_h I__11401 (
            .O(N__57360),
            .I(N__57357));
    Span4Mux_v I__11400 (
            .O(N__57357),
            .I(N__57354));
    Odrv4 I__11399 (
            .O(N__57354),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__11398 (
            .O(N__57351),
            .I(N__57342));
    InMux I__11397 (
            .O(N__57350),
            .I(N__57342));
    InMux I__11396 (
            .O(N__57349),
            .I(N__57342));
    LocalMux I__11395 (
            .O(N__57342),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__11394 (
            .O(N__57339),
            .I(N__57336));
    LocalMux I__11393 (
            .O(N__57336),
            .I(N__57332));
    InMux I__11392 (
            .O(N__57335),
            .I(N__57329));
    Span4Mux_h I__11391 (
            .O(N__57332),
            .I(N__57326));
    LocalMux I__11390 (
            .O(N__57329),
            .I(N__57323));
    Odrv4 I__11389 (
            .O(N__57326),
            .I(front_order_13));
    Odrv4 I__11388 (
            .O(N__57323),
            .I(front_order_13));
    InMux I__11387 (
            .O(N__57318),
            .I(N__57315));
    LocalMux I__11386 (
            .O(N__57315),
            .I(N__57312));
    Span4Mux_h I__11385 (
            .O(N__57312),
            .I(N__57309));
    Odrv4 I__11384 (
            .O(N__57309),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    CascadeMux I__11383 (
            .O(N__57306),
            .I(N__57301));
    InMux I__11382 (
            .O(N__57305),
            .I(N__57294));
    InMux I__11381 (
            .O(N__57304),
            .I(N__57294));
    InMux I__11380 (
            .O(N__57301),
            .I(N__57294));
    LocalMux I__11379 (
            .O(N__57294),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__11378 (
            .O(N__57291),
            .I(N__57288));
    LocalMux I__11377 (
            .O(N__57288),
            .I(N__57284));
    InMux I__11376 (
            .O(N__57287),
            .I(N__57281));
    Span4Mux_h I__11375 (
            .O(N__57284),
            .I(N__57276));
    LocalMux I__11374 (
            .O(N__57281),
            .I(N__57276));
    Span4Mux_h I__11373 (
            .O(N__57276),
            .I(N__57273));
    Span4Mux_h I__11372 (
            .O(N__57273),
            .I(N__57270));
    Odrv4 I__11371 (
            .O(N__57270),
            .I(throttle_order_13));
    CascadeMux I__11370 (
            .O(N__57267),
            .I(N__57264));
    InMux I__11369 (
            .O(N__57264),
            .I(N__57261));
    LocalMux I__11368 (
            .O(N__57261),
            .I(N__57258));
    Span4Mux_h I__11367 (
            .O(N__57258),
            .I(N__57255));
    Odrv4 I__11366 (
            .O(N__57255),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    CascadeMux I__11365 (
            .O(N__57252),
            .I(N__57247));
    InMux I__11364 (
            .O(N__57251),
            .I(N__57240));
    InMux I__11363 (
            .O(N__57250),
            .I(N__57240));
    InMux I__11362 (
            .O(N__57247),
            .I(N__57240));
    LocalMux I__11361 (
            .O(N__57240),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    InMux I__11360 (
            .O(N__57237),
            .I(N__57232));
    InMux I__11359 (
            .O(N__57236),
            .I(N__57227));
    InMux I__11358 (
            .O(N__57235),
            .I(N__57227));
    LocalMux I__11357 (
            .O(N__57232),
            .I(N__57224));
    LocalMux I__11356 (
            .O(N__57227),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    Odrv4 I__11355 (
            .O(N__57224),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__11354 (
            .O(N__57219),
            .I(N__57216));
    LocalMux I__11353 (
            .O(N__57216),
            .I(N__57213));
    Span4Mux_h I__11352 (
            .O(N__57213),
            .I(N__57210));
    Span4Mux_v I__11351 (
            .O(N__57210),
            .I(N__57207));
    Odrv4 I__11350 (
            .O(N__57207),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__11349 (
            .O(N__57204),
            .I(N__57199));
    InMux I__11348 (
            .O(N__57203),
            .I(N__57194));
    InMux I__11347 (
            .O(N__57202),
            .I(N__57194));
    LocalMux I__11346 (
            .O(N__57199),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__11345 (
            .O(N__57194),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__11344 (
            .O(N__57189),
            .I(N__57186));
    InMux I__11343 (
            .O(N__57186),
            .I(N__57182));
    InMux I__11342 (
            .O(N__57185),
            .I(N__57179));
    LocalMux I__11341 (
            .O(N__57182),
            .I(N__57176));
    LocalMux I__11340 (
            .O(N__57179),
            .I(N__57173));
    Span4Mux_h I__11339 (
            .O(N__57176),
            .I(N__57168));
    Span4Mux_h I__11338 (
            .O(N__57173),
            .I(N__57168));
    Odrv4 I__11337 (
            .O(N__57168),
            .I(front_order_1));
    InMux I__11336 (
            .O(N__57165),
            .I(N__57162));
    LocalMux I__11335 (
            .O(N__57162),
            .I(N__57159));
    Odrv4 I__11334 (
            .O(N__57159),
            .I(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ));
    InMux I__11333 (
            .O(N__57156),
            .I(N__57151));
    InMux I__11332 (
            .O(N__57155),
            .I(N__57148));
    InMux I__11331 (
            .O(N__57154),
            .I(N__57145));
    LocalMux I__11330 (
            .O(N__57151),
            .I(N__57142));
    LocalMux I__11329 (
            .O(N__57148),
            .I(N__57139));
    LocalMux I__11328 (
            .O(N__57145),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    Odrv4 I__11327 (
            .O(N__57142),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    Odrv12 I__11326 (
            .O(N__57139),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    CascadeMux I__11325 (
            .O(N__57132),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ));
    CascadeMux I__11324 (
            .O(N__57129),
            .I(N__57125));
    InMux I__11323 (
            .O(N__57128),
            .I(N__57120));
    InMux I__11322 (
            .O(N__57125),
            .I(N__57120));
    LocalMux I__11321 (
            .O(N__57120),
            .I(N__57117));
    Span4Mux_h I__11320 (
            .O(N__57117),
            .I(N__57114));
    Odrv4 I__11319 (
            .O(N__57114),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__11318 (
            .O(N__57111),
            .I(\ppm_encoder_1.N_300_cascade_ ));
    InMux I__11317 (
            .O(N__57108),
            .I(N__57104));
    InMux I__11316 (
            .O(N__57107),
            .I(N__57101));
    LocalMux I__11315 (
            .O(N__57104),
            .I(N__57097));
    LocalMux I__11314 (
            .O(N__57101),
            .I(N__57094));
    InMux I__11313 (
            .O(N__57100),
            .I(N__57091));
    Span4Mux_h I__11312 (
            .O(N__57097),
            .I(N__57088));
    Span4Mux_h I__11311 (
            .O(N__57094),
            .I(N__57085));
    LocalMux I__11310 (
            .O(N__57091),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    Odrv4 I__11309 (
            .O(N__57088),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    Odrv4 I__11308 (
            .O(N__57085),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    InMux I__11307 (
            .O(N__57078),
            .I(N__57075));
    LocalMux I__11306 (
            .O(N__57075),
            .I(N__57072));
    Span4Mux_v I__11305 (
            .O(N__57072),
            .I(N__57069));
    Odrv4 I__11304 (
            .O(N__57069),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    InMux I__11303 (
            .O(N__57066),
            .I(N__57063));
    LocalMux I__11302 (
            .O(N__57063),
            .I(\ppm_encoder_1.N_287 ));
    InMux I__11301 (
            .O(N__57060),
            .I(N__57056));
    InMux I__11300 (
            .O(N__57059),
            .I(N__57053));
    LocalMux I__11299 (
            .O(N__57056),
            .I(N__57049));
    LocalMux I__11298 (
            .O(N__57053),
            .I(N__57046));
    InMux I__11297 (
            .O(N__57052),
            .I(N__57043));
    Span4Mux_v I__11296 (
            .O(N__57049),
            .I(N__57038));
    Span4Mux_v I__11295 (
            .O(N__57046),
            .I(N__57038));
    LocalMux I__11294 (
            .O(N__57043),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__11293 (
            .O(N__57038),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    CascadeMux I__11292 (
            .O(N__57033),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ));
    InMux I__11291 (
            .O(N__57030),
            .I(N__57027));
    LocalMux I__11290 (
            .O(N__57027),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13 ));
    CascadeMux I__11289 (
            .O(N__57024),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ));
    InMux I__11288 (
            .O(N__57021),
            .I(N__57018));
    LocalMux I__11287 (
            .O(N__57018),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4 ));
    CascadeMux I__11286 (
            .O(N__57015),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ));
    InMux I__11285 (
            .O(N__57012),
            .I(N__57009));
    LocalMux I__11284 (
            .O(N__57009),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5 ));
    CascadeMux I__11283 (
            .O(N__57006),
            .I(N__57002));
    InMux I__11282 (
            .O(N__57005),
            .I(N__56996));
    InMux I__11281 (
            .O(N__57002),
            .I(N__56996));
    CascadeMux I__11280 (
            .O(N__57001),
            .I(N__56993));
    LocalMux I__11279 (
            .O(N__56996),
            .I(N__56990));
    InMux I__11278 (
            .O(N__56993),
            .I(N__56987));
    Span4Mux_v I__11277 (
            .O(N__56990),
            .I(N__56984));
    LocalMux I__11276 (
            .O(N__56987),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__11275 (
            .O(N__56984),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__11274 (
            .O(N__56979),
            .I(\ppm_encoder_1.N_291_cascade_ ));
    InMux I__11273 (
            .O(N__56976),
            .I(N__56973));
    LocalMux I__11272 (
            .O(N__56973),
            .I(N__56970));
    Span4Mux_h I__11271 (
            .O(N__56970),
            .I(N__56967));
    Odrv4 I__11270 (
            .O(N__56967),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    InMux I__11269 (
            .O(N__56964),
            .I(N__56955));
    InMux I__11268 (
            .O(N__56963),
            .I(N__56955));
    InMux I__11267 (
            .O(N__56962),
            .I(N__56955));
    LocalMux I__11266 (
            .O(N__56955),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__11265 (
            .O(N__56952),
            .I(N__56948));
    CascadeMux I__11264 (
            .O(N__56951),
            .I(N__56945));
    LocalMux I__11263 (
            .O(N__56948),
            .I(N__56941));
    InMux I__11262 (
            .O(N__56945),
            .I(N__56938));
    InMux I__11261 (
            .O(N__56944),
            .I(N__56935));
    Span4Mux_h I__11260 (
            .O(N__56941),
            .I(N__56932));
    LocalMux I__11259 (
            .O(N__56938),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    LocalMux I__11258 (
            .O(N__56935),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__11257 (
            .O(N__56932),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    CascadeMux I__11256 (
            .O(N__56925),
            .I(N__56921));
    InMux I__11255 (
            .O(N__56924),
            .I(N__56918));
    InMux I__11254 (
            .O(N__56921),
            .I(N__56915));
    LocalMux I__11253 (
            .O(N__56918),
            .I(N__56911));
    LocalMux I__11252 (
            .O(N__56915),
            .I(N__56908));
    InMux I__11251 (
            .O(N__56914),
            .I(N__56905));
    Span4Mux_h I__11250 (
            .O(N__56911),
            .I(N__56902));
    Span4Mux_h I__11249 (
            .O(N__56908),
            .I(N__56899));
    LocalMux I__11248 (
            .O(N__56905),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__11247 (
            .O(N__56902),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__11246 (
            .O(N__56899),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    CascadeMux I__11245 (
            .O(N__56892),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ));
    InMux I__11244 (
            .O(N__56889),
            .I(N__56886));
    LocalMux I__11243 (
            .O(N__56886),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9 ));
    InMux I__11242 (
            .O(N__56883),
            .I(N__56879));
    InMux I__11241 (
            .O(N__56882),
            .I(N__56876));
    LocalMux I__11240 (
            .O(N__56879),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    LocalMux I__11239 (
            .O(N__56876),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    InMux I__11238 (
            .O(N__56871),
            .I(N__56868));
    LocalMux I__11237 (
            .O(N__56868),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    InMux I__11236 (
            .O(N__56865),
            .I(N__56861));
    InMux I__11235 (
            .O(N__56864),
            .I(N__56858));
    LocalMux I__11234 (
            .O(N__56861),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11233 (
            .O(N__56858),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    CascadeMux I__11232 (
            .O(N__56853),
            .I(\ppm_encoder_1.N_221_cascade_ ));
    InMux I__11231 (
            .O(N__56850),
            .I(N__56841));
    InMux I__11230 (
            .O(N__56849),
            .I(N__56841));
    InMux I__11229 (
            .O(N__56848),
            .I(N__56841));
    LocalMux I__11228 (
            .O(N__56841),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    CascadeMux I__11227 (
            .O(N__56838),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ));
    InMux I__11226 (
            .O(N__56835),
            .I(N__56832));
    LocalMux I__11225 (
            .O(N__56832),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    InMux I__11224 (
            .O(N__56829),
            .I(N__56826));
    LocalMux I__11223 (
            .O(N__56826),
            .I(N__56823));
    Odrv4 I__11222 (
            .O(N__56823),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    CascadeMux I__11221 (
            .O(N__56820),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ));
    InMux I__11220 (
            .O(N__56817),
            .I(N__56814));
    LocalMux I__11219 (
            .O(N__56814),
            .I(N__56811));
    Odrv4 I__11218 (
            .O(N__56811),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    InMux I__11217 (
            .O(N__56808),
            .I(N__56804));
    InMux I__11216 (
            .O(N__56807),
            .I(N__56799));
    LocalMux I__11215 (
            .O(N__56804),
            .I(N__56795));
    InMux I__11214 (
            .O(N__56803),
            .I(N__56790));
    InMux I__11213 (
            .O(N__56802),
            .I(N__56790));
    LocalMux I__11212 (
            .O(N__56799),
            .I(N__56787));
    InMux I__11211 (
            .O(N__56798),
            .I(N__56784));
    Span4Mux_v I__11210 (
            .O(N__56795),
            .I(N__56779));
    LocalMux I__11209 (
            .O(N__56790),
            .I(N__56779));
    Odrv4 I__11208 (
            .O(N__56787),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    LocalMux I__11207 (
            .O(N__56784),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__11206 (
            .O(N__56779),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    CascadeMux I__11205 (
            .O(N__56772),
            .I(\ppm_encoder_1.N_286_cascade_ ));
    InMux I__11204 (
            .O(N__56769),
            .I(N__56766));
    LocalMux I__11203 (
            .O(N__56766),
            .I(N__56763));
    Odrv12 I__11202 (
            .O(N__56763),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    InMux I__11201 (
            .O(N__56760),
            .I(N__56757));
    LocalMux I__11200 (
            .O(N__56757),
            .I(N__56754));
    Span4Mux_v I__11199 (
            .O(N__56754),
            .I(N__56751));
    Span4Mux_v I__11198 (
            .O(N__56751),
            .I(N__56748));
    Odrv4 I__11197 (
            .O(N__56748),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__11196 (
            .O(N__56745),
            .I(N__56742));
    LocalMux I__11195 (
            .O(N__56742),
            .I(N__56739));
    Span4Mux_h I__11194 (
            .O(N__56739),
            .I(N__56736));
    Odrv4 I__11193 (
            .O(N__56736),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    CascadeMux I__11192 (
            .O(N__56733),
            .I(N__56730));
    InMux I__11191 (
            .O(N__56730),
            .I(N__56727));
    LocalMux I__11190 (
            .O(N__56727),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__11189 (
            .O(N__56724),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__11188 (
            .O(N__56721),
            .I(N__56717));
    InMux I__11187 (
            .O(N__56720),
            .I(N__56714));
    LocalMux I__11186 (
            .O(N__56717),
            .I(N__56709));
    LocalMux I__11185 (
            .O(N__56714),
            .I(N__56706));
    InMux I__11184 (
            .O(N__56713),
            .I(N__56701));
    InMux I__11183 (
            .O(N__56712),
            .I(N__56701));
    Span4Mux_v I__11182 (
            .O(N__56709),
            .I(N__56698));
    Span4Mux_h I__11181 (
            .O(N__56706),
            .I(N__56695));
    LocalMux I__11180 (
            .O(N__56701),
            .I(N__56692));
    Odrv4 I__11179 (
            .O(N__56698),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__11178 (
            .O(N__56695),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__11177 (
            .O(N__56692),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__11176 (
            .O(N__56685),
            .I(N__56680));
    InMux I__11175 (
            .O(N__56684),
            .I(N__56677));
    InMux I__11174 (
            .O(N__56683),
            .I(N__56674));
    LocalMux I__11173 (
            .O(N__56680),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__11172 (
            .O(N__56677),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__11171 (
            .O(N__56674),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    CascadeMux I__11170 (
            .O(N__56667),
            .I(N__56664));
    InMux I__11169 (
            .O(N__56664),
            .I(N__56661));
    LocalMux I__11168 (
            .O(N__56661),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__11167 (
            .O(N__56658),
            .I(N__56655));
    LocalMux I__11166 (
            .O(N__56655),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CascadeMux I__11165 (
            .O(N__56652),
            .I(N__56649));
    InMux I__11164 (
            .O(N__56649),
            .I(N__56646));
    LocalMux I__11163 (
            .O(N__56646),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__11162 (
            .O(N__56643),
            .I(N__56640));
    LocalMux I__11161 (
            .O(N__56640),
            .I(N__56637));
    Span4Mux_v I__11160 (
            .O(N__56637),
            .I(N__56634));
    Odrv4 I__11159 (
            .O(N__56634),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__11158 (
            .O(N__56631),
            .I(N__56628));
    LocalMux I__11157 (
            .O(N__56628),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__11156 (
            .O(N__56625),
            .I(N__56619));
    InMux I__11155 (
            .O(N__56624),
            .I(N__56612));
    InMux I__11154 (
            .O(N__56623),
            .I(N__56612));
    InMux I__11153 (
            .O(N__56622),
            .I(N__56612));
    LocalMux I__11152 (
            .O(N__56619),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__11151 (
            .O(N__56612),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__11150 (
            .O(N__56607),
            .I(N__56602));
    InMux I__11149 (
            .O(N__56606),
            .I(N__56599));
    InMux I__11148 (
            .O(N__56605),
            .I(N__56596));
    LocalMux I__11147 (
            .O(N__56602),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__11146 (
            .O(N__56599),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__11145 (
            .O(N__56596),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__11144 (
            .O(N__56589),
            .I(N__56586));
    LocalMux I__11143 (
            .O(N__56586),
            .I(N__56583));
    Span4Mux_s3_v I__11142 (
            .O(N__56583),
            .I(N__56580));
    Odrv4 I__11141 (
            .O(N__56580),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    CascadeMux I__11140 (
            .O(N__56577),
            .I(N__56574));
    InMux I__11139 (
            .O(N__56574),
            .I(N__56571));
    LocalMux I__11138 (
            .O(N__56571),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__11137 (
            .O(N__56568),
            .I(N__56565));
    LocalMux I__11136 (
            .O(N__56565),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__11135 (
            .O(N__56562),
            .I(N__56559));
    LocalMux I__11134 (
            .O(N__56559),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__11133 (
            .O(N__56556),
            .I(N__56553));
    LocalMux I__11132 (
            .O(N__56553),
            .I(N__56550));
    Odrv4 I__11131 (
            .O(N__56550),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__11130 (
            .O(N__56547),
            .I(N__56544));
    LocalMux I__11129 (
            .O(N__56544),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__11128 (
            .O(N__56541),
            .I(N__56538));
    LocalMux I__11127 (
            .O(N__56538),
            .I(\pid_front.N_37_1 ));
    InMux I__11126 (
            .O(N__56535),
            .I(N__56531));
    InMux I__11125 (
            .O(N__56534),
            .I(N__56528));
    LocalMux I__11124 (
            .O(N__56531),
            .I(N__56524));
    LocalMux I__11123 (
            .O(N__56528),
            .I(N__56521));
    CascadeMux I__11122 (
            .O(N__56527),
            .I(N__56516));
    Span4Mux_h I__11121 (
            .O(N__56524),
            .I(N__56509));
    Span4Mux_s1_h I__11120 (
            .O(N__56521),
            .I(N__56506));
    InMux I__11119 (
            .O(N__56520),
            .I(N__56501));
    InMux I__11118 (
            .O(N__56519),
            .I(N__56498));
    InMux I__11117 (
            .O(N__56516),
            .I(N__56492));
    InMux I__11116 (
            .O(N__56515),
            .I(N__56489));
    InMux I__11115 (
            .O(N__56514),
            .I(N__56482));
    InMux I__11114 (
            .O(N__56513),
            .I(N__56482));
    InMux I__11113 (
            .O(N__56512),
            .I(N__56482));
    Span4Mux_v I__11112 (
            .O(N__56509),
            .I(N__56477));
    Span4Mux_h I__11111 (
            .O(N__56506),
            .I(N__56474));
    InMux I__11110 (
            .O(N__56505),
            .I(N__56468));
    InMux I__11109 (
            .O(N__56504),
            .I(N__56468));
    LocalMux I__11108 (
            .O(N__56501),
            .I(N__56462));
    LocalMux I__11107 (
            .O(N__56498),
            .I(N__56462));
    InMux I__11106 (
            .O(N__56497),
            .I(N__56455));
    InMux I__11105 (
            .O(N__56496),
            .I(N__56455));
    InMux I__11104 (
            .O(N__56495),
            .I(N__56455));
    LocalMux I__11103 (
            .O(N__56492),
            .I(N__56452));
    LocalMux I__11102 (
            .O(N__56489),
            .I(N__56447));
    LocalMux I__11101 (
            .O(N__56482),
            .I(N__56447));
    InMux I__11100 (
            .O(N__56481),
            .I(N__56442));
    InMux I__11099 (
            .O(N__56480),
            .I(N__56442));
    Span4Mux_h I__11098 (
            .O(N__56477),
            .I(N__56437));
    Span4Mux_h I__11097 (
            .O(N__56474),
            .I(N__56434));
    InMux I__11096 (
            .O(N__56473),
            .I(N__56431));
    LocalMux I__11095 (
            .O(N__56468),
            .I(N__56428));
    InMux I__11094 (
            .O(N__56467),
            .I(N__56425));
    Span4Mux_v I__11093 (
            .O(N__56462),
            .I(N__56420));
    LocalMux I__11092 (
            .O(N__56455),
            .I(N__56420));
    Span4Mux_v I__11091 (
            .O(N__56452),
            .I(N__56413));
    Span4Mux_v I__11090 (
            .O(N__56447),
            .I(N__56413));
    LocalMux I__11089 (
            .O(N__56442),
            .I(N__56413));
    InMux I__11088 (
            .O(N__56441),
            .I(N__56408));
    InMux I__11087 (
            .O(N__56440),
            .I(N__56408));
    Span4Mux_h I__11086 (
            .O(N__56437),
            .I(N__56403));
    Span4Mux_h I__11085 (
            .O(N__56434),
            .I(N__56403));
    LocalMux I__11084 (
            .O(N__56431),
            .I(\pid_front.error_15 ));
    Odrv4 I__11083 (
            .O(N__56428),
            .I(\pid_front.error_15 ));
    LocalMux I__11082 (
            .O(N__56425),
            .I(\pid_front.error_15 ));
    Odrv4 I__11081 (
            .O(N__56420),
            .I(\pid_front.error_15 ));
    Odrv4 I__11080 (
            .O(N__56413),
            .I(\pid_front.error_15 ));
    LocalMux I__11079 (
            .O(N__56408),
            .I(\pid_front.error_15 ));
    Odrv4 I__11078 (
            .O(N__56403),
            .I(\pid_front.error_15 ));
    InMux I__11077 (
            .O(N__56388),
            .I(N__56385));
    LocalMux I__11076 (
            .O(N__56385),
            .I(\pid_front.N_136 ));
    InMux I__11075 (
            .O(N__56382),
            .I(N__56379));
    LocalMux I__11074 (
            .O(N__56379),
            .I(N__56374));
    InMux I__11073 (
            .O(N__56378),
            .I(N__56371));
    InMux I__11072 (
            .O(N__56377),
            .I(N__56368));
    Span4Mux_h I__11071 (
            .O(N__56374),
            .I(N__56363));
    LocalMux I__11070 (
            .O(N__56371),
            .I(N__56363));
    LocalMux I__11069 (
            .O(N__56368),
            .I(\pid_front.N_63 ));
    Odrv4 I__11068 (
            .O(N__56363),
            .I(\pid_front.N_63 ));
    InMux I__11067 (
            .O(N__56358),
            .I(N__56355));
    LocalMux I__11066 (
            .O(N__56355),
            .I(\pid_front.error_cry_2_0_c_RNI1CZ0Z944 ));
    InMux I__11065 (
            .O(N__56352),
            .I(N__56349));
    LocalMux I__11064 (
            .O(N__56349),
            .I(\pid_front.error_cry_2_0_c_RNI1C944Z0Z_0 ));
    CascadeMux I__11063 (
            .O(N__56346),
            .I(\pid_front.N_110_cascade_ ));
    CascadeMux I__11062 (
            .O(N__56343),
            .I(\pid_front.m10_2_03_3_i_0_cascade_ ));
    InMux I__11061 (
            .O(N__56340),
            .I(N__56337));
    LocalMux I__11060 (
            .O(N__56337),
            .I(\pid_front.m26_2_03_0 ));
    CascadeMux I__11059 (
            .O(N__56334),
            .I(N__56331));
    InMux I__11058 (
            .O(N__56331),
            .I(N__56328));
    LocalMux I__11057 (
            .O(N__56328),
            .I(N__56325));
    Span4Mux_v I__11056 (
            .O(N__56325),
            .I(N__56322));
    Span4Mux_h I__11055 (
            .O(N__56322),
            .I(N__56319));
    Odrv4 I__11054 (
            .O(N__56319),
            .I(\pid_front.error_i_regZ0Z_22 ));
    CascadeMux I__11053 (
            .O(N__56316),
            .I(N__56312));
    CascadeMux I__11052 (
            .O(N__56315),
            .I(N__56309));
    InMux I__11051 (
            .O(N__56312),
            .I(N__56306));
    InMux I__11050 (
            .O(N__56309),
            .I(N__56303));
    LocalMux I__11049 (
            .O(N__56306),
            .I(N__56299));
    LocalMux I__11048 (
            .O(N__56303),
            .I(N__56296));
    CascadeMux I__11047 (
            .O(N__56302),
            .I(N__56293));
    Span4Mux_v I__11046 (
            .O(N__56299),
            .I(N__56289));
    Span4Mux_s2_v I__11045 (
            .O(N__56296),
            .I(N__56286));
    InMux I__11044 (
            .O(N__56293),
            .I(N__56281));
    InMux I__11043 (
            .O(N__56292),
            .I(N__56281));
    Odrv4 I__11042 (
            .O(N__56289),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv4 I__11041 (
            .O(N__56286),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__11040 (
            .O(N__56281),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__11039 (
            .O(N__56274),
            .I(N__56271));
    LocalMux I__11038 (
            .O(N__56271),
            .I(N__56268));
    Odrv4 I__11037 (
            .O(N__56268),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    InMux I__11036 (
            .O(N__56265),
            .I(N__56260));
    InMux I__11035 (
            .O(N__56264),
            .I(N__56257));
    InMux I__11034 (
            .O(N__56263),
            .I(N__56254));
    LocalMux I__11033 (
            .O(N__56260),
            .I(N__56251));
    LocalMux I__11032 (
            .O(N__56257),
            .I(N__56248));
    LocalMux I__11031 (
            .O(N__56254),
            .I(N__56245));
    Span4Mux_v I__11030 (
            .O(N__56251),
            .I(N__56236));
    Span4Mux_h I__11029 (
            .O(N__56248),
            .I(N__56236));
    Span4Mux_s2_v I__11028 (
            .O(N__56245),
            .I(N__56233));
    InMux I__11027 (
            .O(N__56244),
            .I(N__56224));
    InMux I__11026 (
            .O(N__56243),
            .I(N__56224));
    InMux I__11025 (
            .O(N__56242),
            .I(N__56224));
    InMux I__11024 (
            .O(N__56241),
            .I(N__56224));
    Odrv4 I__11023 (
            .O(N__56236),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__11022 (
            .O(N__56233),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__11021 (
            .O(N__56224),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    InMux I__11020 (
            .O(N__56217),
            .I(N__56214));
    LocalMux I__11019 (
            .O(N__56214),
            .I(N__56211));
    Odrv4 I__11018 (
            .O(N__56211),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    CascadeMux I__11017 (
            .O(N__56208),
            .I(N__56204));
    InMux I__11016 (
            .O(N__56207),
            .I(N__56199));
    InMux I__11015 (
            .O(N__56204),
            .I(N__56192));
    InMux I__11014 (
            .O(N__56203),
            .I(N__56192));
    InMux I__11013 (
            .O(N__56202),
            .I(N__56192));
    LocalMux I__11012 (
            .O(N__56199),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__11011 (
            .O(N__56192),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__11010 (
            .O(N__56187),
            .I(N__56181));
    InMux I__11009 (
            .O(N__56186),
            .I(N__56176));
    InMux I__11008 (
            .O(N__56185),
            .I(N__56176));
    InMux I__11007 (
            .O(N__56184),
            .I(N__56173));
    LocalMux I__11006 (
            .O(N__56181),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__11005 (
            .O(N__56176),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__11004 (
            .O(N__56173),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    CascadeMux I__11003 (
            .O(N__56166),
            .I(\pid_front.N_37_1_cascade_ ));
    InMux I__11002 (
            .O(N__56163),
            .I(N__56159));
    InMux I__11001 (
            .O(N__56162),
            .I(N__56153));
    LocalMux I__11000 (
            .O(N__56159),
            .I(N__56150));
    CascadeMux I__10999 (
            .O(N__56158),
            .I(N__56147));
    InMux I__10998 (
            .O(N__56157),
            .I(N__56144));
    InMux I__10997 (
            .O(N__56156),
            .I(N__56141));
    LocalMux I__10996 (
            .O(N__56153),
            .I(N__56138));
    Span4Mux_v I__10995 (
            .O(N__56150),
            .I(N__56135));
    InMux I__10994 (
            .O(N__56147),
            .I(N__56132));
    LocalMux I__10993 (
            .O(N__56144),
            .I(N__56129));
    LocalMux I__10992 (
            .O(N__56141),
            .I(N__56126));
    Span12Mux_h I__10991 (
            .O(N__56138),
            .I(N__56123));
    Sp12to4 I__10990 (
            .O(N__56135),
            .I(N__56120));
    LocalMux I__10989 (
            .O(N__56132),
            .I(N__56117));
    Span4Mux_v I__10988 (
            .O(N__56129),
            .I(N__56112));
    Span4Mux_v I__10987 (
            .O(N__56126),
            .I(N__56112));
    Odrv12 I__10986 (
            .O(N__56123),
            .I(\pid_front.error_13 ));
    Odrv12 I__10985 (
            .O(N__56120),
            .I(\pid_front.error_13 ));
    Odrv4 I__10984 (
            .O(N__56117),
            .I(\pid_front.error_13 ));
    Odrv4 I__10983 (
            .O(N__56112),
            .I(\pid_front.error_13 ));
    InMux I__10982 (
            .O(N__56103),
            .I(N__56099));
    InMux I__10981 (
            .O(N__56102),
            .I(N__56096));
    LocalMux I__10980 (
            .O(N__56099),
            .I(N__56093));
    LocalMux I__10979 (
            .O(N__56096),
            .I(N__56090));
    Span4Mux_h I__10978 (
            .O(N__56093),
            .I(N__56086));
    Span4Mux_s1_h I__10977 (
            .O(N__56090),
            .I(N__56083));
    InMux I__10976 (
            .O(N__56089),
            .I(N__56079));
    Span4Mux_v I__10975 (
            .O(N__56086),
            .I(N__56075));
    Span4Mux_h I__10974 (
            .O(N__56083),
            .I(N__56072));
    InMux I__10973 (
            .O(N__56082),
            .I(N__56069));
    LocalMux I__10972 (
            .O(N__56079),
            .I(N__56066));
    InMux I__10971 (
            .O(N__56078),
            .I(N__56063));
    Span4Mux_h I__10970 (
            .O(N__56075),
            .I(N__56059));
    Span4Mux_h I__10969 (
            .O(N__56072),
            .I(N__56054));
    LocalMux I__10968 (
            .O(N__56069),
            .I(N__56054));
    Span4Mux_v I__10967 (
            .O(N__56066),
            .I(N__56049));
    LocalMux I__10966 (
            .O(N__56063),
            .I(N__56049));
    InMux I__10965 (
            .O(N__56062),
            .I(N__56046));
    Span4Mux_h I__10964 (
            .O(N__56059),
            .I(N__56041));
    Span4Mux_h I__10963 (
            .O(N__56054),
            .I(N__56041));
    Odrv4 I__10962 (
            .O(N__56049),
            .I(\pid_front.error_14 ));
    LocalMux I__10961 (
            .O(N__56046),
            .I(\pid_front.error_14 ));
    Odrv4 I__10960 (
            .O(N__56041),
            .I(\pid_front.error_14 ));
    InMux I__10959 (
            .O(N__56034),
            .I(N__56030));
    InMux I__10958 (
            .O(N__56033),
            .I(N__56025));
    LocalMux I__10957 (
            .O(N__56030),
            .I(N__56022));
    InMux I__10956 (
            .O(N__56029),
            .I(N__56019));
    InMux I__10955 (
            .O(N__56028),
            .I(N__56016));
    LocalMux I__10954 (
            .O(N__56025),
            .I(\pid_front.N_36_0 ));
    Odrv12 I__10953 (
            .O(N__56022),
            .I(\pid_front.N_36_0 ));
    LocalMux I__10952 (
            .O(N__56019),
            .I(\pid_front.N_36_0 ));
    LocalMux I__10951 (
            .O(N__56016),
            .I(\pid_front.N_36_0 ));
    CascadeMux I__10950 (
            .O(N__56007),
            .I(\pid_side.m18_2_03_4_cascade_ ));
    InMux I__10949 (
            .O(N__56004),
            .I(N__56001));
    LocalMux I__10948 (
            .O(N__56001),
            .I(\pid_side.m2_2_03 ));
    InMux I__10947 (
            .O(N__55998),
            .I(N__55995));
    LocalMux I__10946 (
            .O(N__55995),
            .I(N__55991));
    InMux I__10945 (
            .O(N__55994),
            .I(N__55988));
    Span4Mux_v I__10944 (
            .O(N__55991),
            .I(N__55985));
    LocalMux I__10943 (
            .O(N__55988),
            .I(N__55982));
    Span4Mux_v I__10942 (
            .O(N__55985),
            .I(N__55977));
    Span4Mux_v I__10941 (
            .O(N__55982),
            .I(N__55977));
    Odrv4 I__10940 (
            .O(N__55977),
            .I(\pid_front.N_3 ));
    CascadeMux I__10939 (
            .O(N__55974),
            .I(\pid_front.m2_0_03_3_i_0_cascade_ ));
    CascadeMux I__10938 (
            .O(N__55971),
            .I(\pid_front.m2_2_03_cascade_ ));
    CascadeMux I__10937 (
            .O(N__55968),
            .I(\pid_front.error_i_reg_9_rn_1_14_cascade_ ));
    InMux I__10936 (
            .O(N__55965),
            .I(N__55962));
    LocalMux I__10935 (
            .O(N__55962),
            .I(N__55959));
    Span4Mux_h I__10934 (
            .O(N__55959),
            .I(N__55956));
    Span4Mux_v I__10933 (
            .O(N__55956),
            .I(N__55953));
    Odrv4 I__10932 (
            .O(N__55953),
            .I(\pid_front.error_i_regZ0Z_14 ));
    CascadeMux I__10931 (
            .O(N__55950),
            .I(\pid_front.m24_2_03_0_cascade_ ));
    InMux I__10930 (
            .O(N__55947),
            .I(N__55944));
    LocalMux I__10929 (
            .O(N__55944),
            .I(N__55941));
    Odrv12 I__10928 (
            .O(N__55941),
            .I(\pid_front.m8_2_03_3_i_0 ));
    CascadeMux I__10927 (
            .O(N__55938),
            .I(N__55935));
    InMux I__10926 (
            .O(N__55935),
            .I(N__55932));
    LocalMux I__10925 (
            .O(N__55932),
            .I(N__55929));
    Span4Mux_h I__10924 (
            .O(N__55929),
            .I(N__55926));
    Odrv4 I__10923 (
            .O(N__55926),
            .I(\pid_front.error_i_regZ0Z_20 ));
    CascadeMux I__10922 (
            .O(N__55923),
            .I(\pid_front.N_57_0_cascade_ ));
    InMux I__10921 (
            .O(N__55920),
            .I(N__55917));
    LocalMux I__10920 (
            .O(N__55917),
            .I(\pid_front.error_i_reg_esr_RNO_0_0_24 ));
    InMux I__10919 (
            .O(N__55914),
            .I(N__55911));
    LocalMux I__10918 (
            .O(N__55911),
            .I(\pid_front.m138_0_1 ));
    CascadeMux I__10917 (
            .O(N__55908),
            .I(N__55904));
    InMux I__10916 (
            .O(N__55907),
            .I(N__55900));
    InMux I__10915 (
            .O(N__55904),
            .I(N__55895));
    InMux I__10914 (
            .O(N__55903),
            .I(N__55895));
    LocalMux I__10913 (
            .O(N__55900),
            .I(N__55892));
    LocalMux I__10912 (
            .O(N__55895),
            .I(\pid_front.N_22_0 ));
    Odrv4 I__10911 (
            .O(N__55892),
            .I(\pid_front.N_22_0 ));
    InMux I__10910 (
            .O(N__55887),
            .I(N__55881));
    InMux I__10909 (
            .O(N__55886),
            .I(N__55881));
    LocalMux I__10908 (
            .O(N__55881),
            .I(\pid_front.N_57_0 ));
    CascadeMux I__10907 (
            .O(N__55878),
            .I(\pid_front.N_129_cascade_ ));
    CascadeMux I__10906 (
            .O(N__55875),
            .I(N__55872));
    InMux I__10905 (
            .O(N__55872),
            .I(N__55869));
    LocalMux I__10904 (
            .O(N__55869),
            .I(N__55866));
    Span4Mux_h I__10903 (
            .O(N__55866),
            .I(N__55863));
    Span4Mux_v I__10902 (
            .O(N__55863),
            .I(N__55860));
    Odrv4 I__10901 (
            .O(N__55860),
            .I(\pid_front.error_i_regZ0Z_12 ));
    InMux I__10900 (
            .O(N__55857),
            .I(N__55854));
    LocalMux I__10899 (
            .O(N__55854),
            .I(N__55850));
    InMux I__10898 (
            .O(N__55853),
            .I(N__55847));
    Span4Mux_h I__10897 (
            .O(N__55850),
            .I(N__55844));
    LocalMux I__10896 (
            .O(N__55847),
            .I(\pid_front.N_60_0 ));
    Odrv4 I__10895 (
            .O(N__55844),
            .I(\pid_front.N_60_0 ));
    InMux I__10894 (
            .O(N__55839),
            .I(N__55836));
    LocalMux I__10893 (
            .O(N__55836),
            .I(\pid_front.error_i_reg_9_1_12 ));
    InMux I__10892 (
            .O(N__55833),
            .I(N__55830));
    LocalMux I__10891 (
            .O(N__55830),
            .I(N__55826));
    InMux I__10890 (
            .O(N__55829),
            .I(N__55823));
    Span4Mux_s1_h I__10889 (
            .O(N__55826),
            .I(N__55819));
    LocalMux I__10888 (
            .O(N__55823),
            .I(N__55815));
    InMux I__10887 (
            .O(N__55822),
            .I(N__55812));
    Span4Mux_h I__10886 (
            .O(N__55819),
            .I(N__55809));
    InMux I__10885 (
            .O(N__55818),
            .I(N__55806));
    Span12Mux_v I__10884 (
            .O(N__55815),
            .I(N__55801));
    LocalMux I__10883 (
            .O(N__55812),
            .I(N__55798));
    Span4Mux_h I__10882 (
            .O(N__55809),
            .I(N__55792));
    LocalMux I__10881 (
            .O(N__55806),
            .I(N__55792));
    CascadeMux I__10880 (
            .O(N__55805),
            .I(N__55789));
    CascadeMux I__10879 (
            .O(N__55804),
            .I(N__55785));
    Span12Mux_h I__10878 (
            .O(N__55801),
            .I(N__55781));
    Span4Mux_v I__10877 (
            .O(N__55798),
            .I(N__55778));
    InMux I__10876 (
            .O(N__55797),
            .I(N__55775));
    Span4Mux_h I__10875 (
            .O(N__55792),
            .I(N__55772));
    InMux I__10874 (
            .O(N__55789),
            .I(N__55767));
    InMux I__10873 (
            .O(N__55788),
            .I(N__55767));
    InMux I__10872 (
            .O(N__55785),
            .I(N__55762));
    InMux I__10871 (
            .O(N__55784),
            .I(N__55762));
    Odrv12 I__10870 (
            .O(N__55781),
            .I(\pid_front.error_11 ));
    Odrv4 I__10869 (
            .O(N__55778),
            .I(\pid_front.error_11 ));
    LocalMux I__10868 (
            .O(N__55775),
            .I(\pid_front.error_11 ));
    Odrv4 I__10867 (
            .O(N__55772),
            .I(\pid_front.error_11 ));
    LocalMux I__10866 (
            .O(N__55767),
            .I(\pid_front.error_11 ));
    LocalMux I__10865 (
            .O(N__55762),
            .I(\pid_front.error_11 ));
    InMux I__10864 (
            .O(N__55749),
            .I(N__55746));
    LocalMux I__10863 (
            .O(N__55746),
            .I(N__55742));
    InMux I__10862 (
            .O(N__55745),
            .I(N__55737));
    Span4Mux_v I__10861 (
            .O(N__55742),
            .I(N__55734));
    InMux I__10860 (
            .O(N__55741),
            .I(N__55731));
    InMux I__10859 (
            .O(N__55740),
            .I(N__55728));
    LocalMux I__10858 (
            .O(N__55737),
            .I(N__55724));
    Span4Mux_h I__10857 (
            .O(N__55734),
            .I(N__55720));
    LocalMux I__10856 (
            .O(N__55731),
            .I(N__55717));
    LocalMux I__10855 (
            .O(N__55728),
            .I(N__55714));
    CascadeMux I__10854 (
            .O(N__55727),
            .I(N__55711));
    Span4Mux_v I__10853 (
            .O(N__55724),
            .I(N__55707));
    InMux I__10852 (
            .O(N__55723),
            .I(N__55704));
    Span4Mux_h I__10851 (
            .O(N__55720),
            .I(N__55701));
    Span4Mux_v I__10850 (
            .O(N__55717),
            .I(N__55696));
    Span4Mux_v I__10849 (
            .O(N__55714),
            .I(N__55696));
    InMux I__10848 (
            .O(N__55711),
            .I(N__55691));
    InMux I__10847 (
            .O(N__55710),
            .I(N__55691));
    Sp12to4 I__10846 (
            .O(N__55707),
            .I(N__55688));
    LocalMux I__10845 (
            .O(N__55704),
            .I(N__55683));
    Span4Mux_h I__10844 (
            .O(N__55701),
            .I(N__55683));
    Odrv4 I__10843 (
            .O(N__55696),
            .I(\pid_front.error_12 ));
    LocalMux I__10842 (
            .O(N__55691),
            .I(\pid_front.error_12 ));
    Odrv12 I__10841 (
            .O(N__55688),
            .I(\pid_front.error_12 ));
    Odrv4 I__10840 (
            .O(N__55683),
            .I(\pid_front.error_12 ));
    InMux I__10839 (
            .O(N__55674),
            .I(N__55671));
    LocalMux I__10838 (
            .O(N__55671),
            .I(\pid_front.N_18_1 ));
    CascadeMux I__10837 (
            .O(N__55668),
            .I(\pid_front.N_18_1_cascade_ ));
    CascadeMux I__10836 (
            .O(N__55665),
            .I(\pid_side.N_11_0_cascade_ ));
    InMux I__10835 (
            .O(N__55662),
            .I(N__55653));
    InMux I__10834 (
            .O(N__55661),
            .I(N__55653));
    InMux I__10833 (
            .O(N__55660),
            .I(N__55653));
    LocalMux I__10832 (
            .O(N__55653),
            .I(\pid_side.N_14_1 ));
    InMux I__10831 (
            .O(N__55650),
            .I(N__55644));
    InMux I__10830 (
            .O(N__55649),
            .I(N__55644));
    LocalMux I__10829 (
            .O(N__55644),
            .I(\pid_side.N_11_0 ));
    CascadeMux I__10828 (
            .O(N__55641),
            .I(\pid_side.N_104_cascade_ ));
    CascadeMux I__10827 (
            .O(N__55638),
            .I(\pid_side.error_i_reg_9_1_15_cascade_ ));
    InMux I__10826 (
            .O(N__55635),
            .I(N__55632));
    LocalMux I__10825 (
            .O(N__55632),
            .I(\pid_side.m19_2_03_0 ));
    CascadeMux I__10824 (
            .O(N__55629),
            .I(\pid_side.N_41_0_cascade_ ));
    InMux I__10823 (
            .O(N__55626),
            .I(N__55623));
    LocalMux I__10822 (
            .O(N__55623),
            .I(\pid_side.error_i_reg_9_rn_0_26 ));
    CascadeMux I__10821 (
            .O(N__55620),
            .I(\pid_front.m8_2_03_3_i_0_cascade_ ));
    CascadeMux I__10820 (
            .O(N__55617),
            .I(N__55613));
    InMux I__10819 (
            .O(N__55616),
            .I(N__55610));
    InMux I__10818 (
            .O(N__55613),
            .I(N__55607));
    LocalMux I__10817 (
            .O(N__55610),
            .I(N__55604));
    LocalMux I__10816 (
            .O(N__55607),
            .I(N__55601));
    Span4Mux_h I__10815 (
            .O(N__55604),
            .I(N__55596));
    Span4Mux_h I__10814 (
            .O(N__55601),
            .I(N__55596));
    Odrv4 I__10813 (
            .O(N__55596),
            .I(\pid_front.error_i_regZ0Z_4 ));
    CascadeMux I__10812 (
            .O(N__55593),
            .I(N__55589));
    InMux I__10811 (
            .O(N__55592),
            .I(N__55584));
    InMux I__10810 (
            .O(N__55589),
            .I(N__55584));
    LocalMux I__10809 (
            .O(N__55584),
            .I(N__55580));
    InMux I__10808 (
            .O(N__55583),
            .I(N__55577));
    Span4Mux_h I__10807 (
            .O(N__55580),
            .I(N__55574));
    LocalMux I__10806 (
            .O(N__55577),
            .I(N__55571));
    Span4Mux_v I__10805 (
            .O(N__55574),
            .I(N__55568));
    Span4Mux_v I__10804 (
            .O(N__55571),
            .I(N__55565));
    Span4Mux_v I__10803 (
            .O(N__55568),
            .I(N__55562));
    Span4Mux_v I__10802 (
            .O(N__55565),
            .I(N__55559));
    Odrv4 I__10801 (
            .O(N__55562),
            .I(\pid_front.state_ns_0 ));
    Odrv4 I__10800 (
            .O(N__55559),
            .I(\pid_front.state_ns_0 ));
    InMux I__10799 (
            .O(N__55554),
            .I(N__55551));
    LocalMux I__10798 (
            .O(N__55551),
            .I(N__55547));
    InMux I__10797 (
            .O(N__55550),
            .I(N__55544));
    Odrv12 I__10796 (
            .O(N__55547),
            .I(\pid_front.N_54_0 ));
    LocalMux I__10795 (
            .O(N__55544),
            .I(\pid_front.N_54_0 ));
    CascadeMux I__10794 (
            .O(N__55539),
            .I(N__55536));
    InMux I__10793 (
            .O(N__55536),
            .I(N__55533));
    LocalMux I__10792 (
            .O(N__55533),
            .I(N__55529));
    InMux I__10791 (
            .O(N__55532),
            .I(N__55526));
    Span4Mux_h I__10790 (
            .O(N__55529),
            .I(N__55523));
    LocalMux I__10789 (
            .O(N__55526),
            .I(\pid_front.error_i_regZ0Z_11 ));
    Odrv4 I__10788 (
            .O(N__55523),
            .I(\pid_front.error_i_regZ0Z_11 ));
    InMux I__10787 (
            .O(N__55518),
            .I(N__55515));
    LocalMux I__10786 (
            .O(N__55515),
            .I(N__55511));
    InMux I__10785 (
            .O(N__55514),
            .I(N__55508));
    Span4Mux_v I__10784 (
            .O(N__55511),
            .I(N__55501));
    LocalMux I__10783 (
            .O(N__55508),
            .I(N__55501));
    InMux I__10782 (
            .O(N__55507),
            .I(N__55498));
    InMux I__10781 (
            .O(N__55506),
            .I(N__55495));
    Odrv4 I__10780 (
            .O(N__55501),
            .I(\pid_front.N_15_1 ));
    LocalMux I__10779 (
            .O(N__55498),
            .I(\pid_front.N_15_1 ));
    LocalMux I__10778 (
            .O(N__55495),
            .I(\pid_front.N_15_1 ));
    InMux I__10777 (
            .O(N__55488),
            .I(N__55485));
    LocalMux I__10776 (
            .O(N__55485),
            .I(\pid_front.m3_2_03 ));
    InMux I__10775 (
            .O(N__55482),
            .I(N__55479));
    LocalMux I__10774 (
            .O(N__55479),
            .I(N__55476));
    Odrv4 I__10773 (
            .O(N__55476),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_7 ));
    CascadeMux I__10772 (
            .O(N__55473),
            .I(\pid_side.N_49_0_cascade_ ));
    CascadeMux I__10771 (
            .O(N__55470),
            .I(\pid_side.m134_0_ns_1_cascade_ ));
    CascadeMux I__10770 (
            .O(N__55467),
            .I(N__55463));
    InMux I__10769 (
            .O(N__55466),
            .I(N__55460));
    InMux I__10768 (
            .O(N__55463),
            .I(N__55457));
    LocalMux I__10767 (
            .O(N__55460),
            .I(N__55452));
    LocalMux I__10766 (
            .O(N__55457),
            .I(N__55452));
    Span12Mux_v I__10765 (
            .O(N__55452),
            .I(N__55449));
    Odrv12 I__10764 (
            .O(N__55449),
            .I(\ppm_encoder_1.N_2569_i ));
    CascadeMux I__10763 (
            .O(N__55446),
            .I(pid_front_N_331_cascade_));
    CascadeMux I__10762 (
            .O(N__55443),
            .I(pid_side_N_166_mux_cascade_));
    InMux I__10761 (
            .O(N__55440),
            .I(N__55437));
    LocalMux I__10760 (
            .O(N__55437),
            .I(N__55433));
    InMux I__10759 (
            .O(N__55436),
            .I(N__55430));
    Span4Mux_v I__10758 (
            .O(N__55433),
            .I(N__55423));
    LocalMux I__10757 (
            .O(N__55430),
            .I(N__55423));
    InMux I__10756 (
            .O(N__55429),
            .I(N__55418));
    InMux I__10755 (
            .O(N__55428),
            .I(N__55418));
    Odrv4 I__10754 (
            .O(N__55423),
            .I(\pid_front.N_39_0 ));
    LocalMux I__10753 (
            .O(N__55418),
            .I(\pid_front.N_39_0 ));
    CascadeMux I__10752 (
            .O(N__55413),
            .I(N__55410));
    InMux I__10751 (
            .O(N__55410),
            .I(N__55407));
    LocalMux I__10750 (
            .O(N__55407),
            .I(N__55404));
    Span4Mux_h I__10749 (
            .O(N__55404),
            .I(N__55401));
    Odrv4 I__10748 (
            .O(N__55401),
            .I(\pid_front.error_i_regZ0Z_3 ));
    InMux I__10747 (
            .O(N__55398),
            .I(N__55395));
    LocalMux I__10746 (
            .O(N__55395),
            .I(N__55391));
    InMux I__10745 (
            .O(N__55394),
            .I(N__55388));
    Span4Mux_h I__10744 (
            .O(N__55391),
            .I(N__55382));
    LocalMux I__10743 (
            .O(N__55388),
            .I(N__55382));
    InMux I__10742 (
            .O(N__55387),
            .I(N__55379));
    Odrv4 I__10741 (
            .O(N__55382),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__10740 (
            .O(N__55379),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    InMux I__10739 (
            .O(N__55374),
            .I(N__55370));
    InMux I__10738 (
            .O(N__55373),
            .I(N__55367));
    LocalMux I__10737 (
            .O(N__55370),
            .I(N__55361));
    LocalMux I__10736 (
            .O(N__55367),
            .I(N__55361));
    InMux I__10735 (
            .O(N__55366),
            .I(N__55358));
    Odrv12 I__10734 (
            .O(N__55361),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__10733 (
            .O(N__55358),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    InMux I__10732 (
            .O(N__55353),
            .I(N__55350));
    LocalMux I__10731 (
            .O(N__55350),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ));
    InMux I__10730 (
            .O(N__55347),
            .I(N__55344));
    LocalMux I__10729 (
            .O(N__55344),
            .I(N__55339));
    InMux I__10728 (
            .O(N__55343),
            .I(N__55336));
    InMux I__10727 (
            .O(N__55342),
            .I(N__55333));
    Span4Mux_v I__10726 (
            .O(N__55339),
            .I(N__55330));
    LocalMux I__10725 (
            .O(N__55336),
            .I(\pid_side.un10lto12 ));
    LocalMux I__10724 (
            .O(N__55333),
            .I(\pid_side.un10lto12 ));
    Odrv4 I__10723 (
            .O(N__55330),
            .I(\pid_side.un10lto12 ));
    CascadeMux I__10722 (
            .O(N__55323),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ));
    InMux I__10721 (
            .O(N__55320),
            .I(N__55317));
    LocalMux I__10720 (
            .O(N__55317),
            .I(N__55314));
    Odrv12 I__10719 (
            .O(N__55314),
            .I(\pid_side.error_i_acumm16lt9_0 ));
    InMux I__10718 (
            .O(N__55311),
            .I(N__55308));
    LocalMux I__10717 (
            .O(N__55308),
            .I(N__55305));
    Odrv4 I__10716 (
            .O(N__55305),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ));
    InMux I__10715 (
            .O(N__55302),
            .I(N__55299));
    LocalMux I__10714 (
            .O(N__55299),
            .I(N__55294));
    InMux I__10713 (
            .O(N__55298),
            .I(N__55289));
    InMux I__10712 (
            .O(N__55297),
            .I(N__55289));
    Odrv4 I__10711 (
            .O(N__55294),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__10710 (
            .O(N__55289),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    InMux I__10709 (
            .O(N__55284),
            .I(N__55281));
    LocalMux I__10708 (
            .O(N__55281),
            .I(N__55278));
    Odrv12 I__10707 (
            .O(N__55278),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ));
    InMux I__10706 (
            .O(N__55275),
            .I(N__55272));
    LocalMux I__10705 (
            .O(N__55272),
            .I(N__55269));
    Span4Mux_v I__10704 (
            .O(N__55269),
            .I(N__55264));
    InMux I__10703 (
            .O(N__55268),
            .I(N__55259));
    InMux I__10702 (
            .O(N__55267),
            .I(N__55259));
    Odrv4 I__10701 (
            .O(N__55264),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__10700 (
            .O(N__55259),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    InMux I__10699 (
            .O(N__55254),
            .I(N__55250));
    InMux I__10698 (
            .O(N__55253),
            .I(N__55247));
    LocalMux I__10697 (
            .O(N__55250),
            .I(N__55242));
    LocalMux I__10696 (
            .O(N__55247),
            .I(N__55242));
    Span4Mux_v I__10695 (
            .O(N__55242),
            .I(N__55238));
    InMux I__10694 (
            .O(N__55241),
            .I(N__55235));
    Odrv4 I__10693 (
            .O(N__55238),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__10692 (
            .O(N__55235),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    InMux I__10691 (
            .O(N__55230),
            .I(N__55227));
    LocalMux I__10690 (
            .O(N__55227),
            .I(N__55223));
    InMux I__10689 (
            .O(N__55226),
            .I(N__55220));
    Span4Mux_h I__10688 (
            .O(N__55223),
            .I(N__55215));
    LocalMux I__10687 (
            .O(N__55220),
            .I(N__55215));
    Odrv4 I__10686 (
            .O(N__55215),
            .I(\pid_side.error_i_acumm_preregZ0Z_0 ));
    InMux I__10685 (
            .O(N__55212),
            .I(N__55209));
    LocalMux I__10684 (
            .O(N__55209),
            .I(N__55204));
    InMux I__10683 (
            .O(N__55208),
            .I(N__55199));
    InMux I__10682 (
            .O(N__55207),
            .I(N__55199));
    Odrv4 I__10681 (
            .O(N__55204),
            .I(\pid_side.error_i_acumm_preregZ0Z_13 ));
    LocalMux I__10680 (
            .O(N__55199),
            .I(\pid_side.error_i_acumm_preregZ0Z_13 ));
    CascadeMux I__10679 (
            .O(N__55194),
            .I(N__55191));
    InMux I__10678 (
            .O(N__55191),
            .I(N__55185));
    InMux I__10677 (
            .O(N__55190),
            .I(N__55185));
    LocalMux I__10676 (
            .O(N__55185),
            .I(\pid_side.error_i_acumm_preregZ0Z_23 ));
    InMux I__10675 (
            .O(N__55182),
            .I(N__55176));
    InMux I__10674 (
            .O(N__55181),
            .I(N__55176));
    LocalMux I__10673 (
            .O(N__55176),
            .I(\pid_side.error_i_acumm_preregZ0Z_22 ));
    InMux I__10672 (
            .O(N__55173),
            .I(N__55167));
    InMux I__10671 (
            .O(N__55172),
            .I(N__55167));
    LocalMux I__10670 (
            .O(N__55167),
            .I(\pid_side.error_i_acumm_preregZ0Z_24 ));
    InMux I__10669 (
            .O(N__55164),
            .I(N__55146));
    InMux I__10668 (
            .O(N__55163),
            .I(N__55146));
    InMux I__10667 (
            .O(N__55162),
            .I(N__55146));
    InMux I__10666 (
            .O(N__55161),
            .I(N__55146));
    InMux I__10665 (
            .O(N__55160),
            .I(N__55146));
    InMux I__10664 (
            .O(N__55159),
            .I(N__55146));
    LocalMux I__10663 (
            .O(N__55146),
            .I(\pid_side.error_i_acumm_2_sqmuxa_1 ));
    InMux I__10662 (
            .O(N__55143),
            .I(N__55128));
    InMux I__10661 (
            .O(N__55142),
            .I(N__55128));
    InMux I__10660 (
            .O(N__55141),
            .I(N__55128));
    InMux I__10659 (
            .O(N__55140),
            .I(N__55128));
    InMux I__10658 (
            .O(N__55139),
            .I(N__55128));
    LocalMux I__10657 (
            .O(N__55128),
            .I(N__55117));
    InMux I__10656 (
            .O(N__55127),
            .I(N__55110));
    InMux I__10655 (
            .O(N__55126),
            .I(N__55110));
    InMux I__10654 (
            .O(N__55125),
            .I(N__55110));
    InMux I__10653 (
            .O(N__55124),
            .I(N__55099));
    InMux I__10652 (
            .O(N__55123),
            .I(N__55099));
    InMux I__10651 (
            .O(N__55122),
            .I(N__55099));
    InMux I__10650 (
            .O(N__55121),
            .I(N__55099));
    InMux I__10649 (
            .O(N__55120),
            .I(N__55099));
    Odrv4 I__10648 (
            .O(N__55117),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    LocalMux I__10647 (
            .O(N__55110),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    LocalMux I__10646 (
            .O(N__55099),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    CEMux I__10645 (
            .O(N__55092),
            .I(N__55088));
    CEMux I__10644 (
            .O(N__55091),
            .I(N__55085));
    LocalMux I__10643 (
            .O(N__55088),
            .I(N__55081));
    LocalMux I__10642 (
            .O(N__55085),
            .I(N__55078));
    CEMux I__10641 (
            .O(N__55084),
            .I(N__55075));
    Span4Mux_v I__10640 (
            .O(N__55081),
            .I(N__55072));
    Span4Mux_v I__10639 (
            .O(N__55078),
            .I(N__55067));
    LocalMux I__10638 (
            .O(N__55075),
            .I(N__55067));
    Odrv4 I__10637 (
            .O(N__55072),
            .I(\pid_side.error_i_acumm_1_sqmuxa_1_i ));
    Odrv4 I__10636 (
            .O(N__55067),
            .I(\pid_side.error_i_acumm_1_sqmuxa_1_i ));
    InMux I__10635 (
            .O(N__55062),
            .I(N__55059));
    LocalMux I__10634 (
            .O(N__55059),
            .I(\pid_side.error_i_acumm16lto27_10 ));
    InMux I__10633 (
            .O(N__55056),
            .I(N__55053));
    LocalMux I__10632 (
            .O(N__55053),
            .I(\pid_side.error_i_acumm16lto27_8 ));
    CascadeMux I__10631 (
            .O(N__55050),
            .I(\pid_side.error_i_acumm16lto27_9_cascade_ ));
    InMux I__10630 (
            .O(N__55047),
            .I(N__55044));
    LocalMux I__10629 (
            .O(N__55044),
            .I(\pid_side.error_i_acumm16lto27_7 ));
    InMux I__10628 (
            .O(N__55041),
            .I(N__55038));
    LocalMux I__10627 (
            .O(N__55038),
            .I(\pid_side.error_i_acumm16lto27_13 ));
    CascadeMux I__10626 (
            .O(N__55035),
            .I(\pid_side.un10lto27_8_cascade_ ));
    CascadeMux I__10625 (
            .O(N__55032),
            .I(N__55029));
    InMux I__10624 (
            .O(N__55029),
            .I(N__55023));
    InMux I__10623 (
            .O(N__55028),
            .I(N__55023));
    LocalMux I__10622 (
            .O(N__55023),
            .I(\pid_side.error_i_acumm_preregZ0Z_26 ));
    CascadeMux I__10621 (
            .O(N__55020),
            .I(\pid_side.un10lt9_1_cascade_ ));
    CascadeMux I__10620 (
            .O(N__55017),
            .I(\pid_side.un10lt9_cascade_ ));
    CascadeMux I__10619 (
            .O(N__55014),
            .I(\pid_side.un10lt11_0_cascade_ ));
    CascadeMux I__10618 (
            .O(N__55011),
            .I(N__55008));
    InMux I__10617 (
            .O(N__55008),
            .I(N__55004));
    InMux I__10616 (
            .O(N__55007),
            .I(N__55000));
    LocalMux I__10615 (
            .O(N__55004),
            .I(N__54996));
    InMux I__10614 (
            .O(N__55003),
            .I(N__54993));
    LocalMux I__10613 (
            .O(N__55000),
            .I(N__54990));
    InMux I__10612 (
            .O(N__54999),
            .I(N__54987));
    Span4Mux_v I__10611 (
            .O(N__54996),
            .I(N__54984));
    LocalMux I__10610 (
            .O(N__54993),
            .I(N__54979));
    Span4Mux_h I__10609 (
            .O(N__54990),
            .I(N__54974));
    LocalMux I__10608 (
            .O(N__54987),
            .I(N__54974));
    Span4Mux_h I__10607 (
            .O(N__54984),
            .I(N__54969));
    InMux I__10606 (
            .O(N__54983),
            .I(N__54964));
    InMux I__10605 (
            .O(N__54982),
            .I(N__54961));
    Span4Mux_v I__10604 (
            .O(N__54979),
            .I(N__54958));
    Span4Mux_v I__10603 (
            .O(N__54974),
            .I(N__54955));
    InMux I__10602 (
            .O(N__54973),
            .I(N__54952));
    InMux I__10601 (
            .O(N__54972),
            .I(N__54949));
    Span4Mux_h I__10600 (
            .O(N__54969),
            .I(N__54946));
    InMux I__10599 (
            .O(N__54968),
            .I(N__54941));
    InMux I__10598 (
            .O(N__54967),
            .I(N__54941));
    LocalMux I__10597 (
            .O(N__54964),
            .I(N__54938));
    LocalMux I__10596 (
            .O(N__54961),
            .I(N__54933));
    Span4Mux_h I__10595 (
            .O(N__54958),
            .I(N__54933));
    Span4Mux_h I__10594 (
            .O(N__54955),
            .I(N__54928));
    LocalMux I__10593 (
            .O(N__54952),
            .I(N__54928));
    LocalMux I__10592 (
            .O(N__54949),
            .I(N__54925));
    Sp12to4 I__10591 (
            .O(N__54946),
            .I(N__54922));
    LocalMux I__10590 (
            .O(N__54941),
            .I(N__54919));
    Span4Mux_h I__10589 (
            .O(N__54938),
            .I(N__54912));
    Span4Mux_h I__10588 (
            .O(N__54933),
            .I(N__54912));
    Span4Mux_h I__10587 (
            .O(N__54928),
            .I(N__54912));
    Span4Mux_v I__10586 (
            .O(N__54925),
            .I(N__54909));
    Span12Mux_v I__10585 (
            .O(N__54922),
            .I(N__54904));
    Sp12to4 I__10584 (
            .O(N__54919),
            .I(N__54904));
    Sp12to4 I__10583 (
            .O(N__54912),
            .I(N__54901));
    Sp12to4 I__10582 (
            .O(N__54909),
            .I(N__54895));
    Span12Mux_v I__10581 (
            .O(N__54904),
            .I(N__54895));
    Span12Mux_v I__10580 (
            .O(N__54901),
            .I(N__54892));
    IoInMux I__10579 (
            .O(N__54900),
            .I(N__54889));
    Odrv12 I__10578 (
            .O(N__54895),
            .I(reset_system));
    Odrv12 I__10577 (
            .O(N__54892),
            .I(reset_system));
    LocalMux I__10576 (
            .O(N__54889),
            .I(reset_system));
    CascadeMux I__10575 (
            .O(N__54882),
            .I(\pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ));
    InMux I__10574 (
            .O(N__54879),
            .I(N__54876));
    LocalMux I__10573 (
            .O(N__54876),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ));
    CascadeMux I__10572 (
            .O(N__54873),
            .I(\pid_side.error_i_acumm_2_sqmuxa_cascade_ ));
    InMux I__10571 (
            .O(N__54870),
            .I(N__54865));
    InMux I__10570 (
            .O(N__54869),
            .I(N__54860));
    InMux I__10569 (
            .O(N__54868),
            .I(N__54860));
    LocalMux I__10568 (
            .O(N__54865),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    LocalMux I__10567 (
            .O(N__54860),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    CascadeMux I__10566 (
            .O(N__54855),
            .I(N__54852));
    InMux I__10565 (
            .O(N__54852),
            .I(N__54849));
    LocalMux I__10564 (
            .O(N__54849),
            .I(N__54844));
    InMux I__10563 (
            .O(N__54848),
            .I(N__54839));
    InMux I__10562 (
            .O(N__54847),
            .I(N__54839));
    Odrv4 I__10561 (
            .O(N__54844),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    LocalMux I__10560 (
            .O(N__54839),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    CascadeMux I__10559 (
            .O(N__54834),
            .I(N__54831));
    InMux I__10558 (
            .O(N__54831),
            .I(N__54827));
    CascadeMux I__10557 (
            .O(N__54830),
            .I(N__54823));
    LocalMux I__10556 (
            .O(N__54827),
            .I(N__54820));
    InMux I__10555 (
            .O(N__54826),
            .I(N__54817));
    InMux I__10554 (
            .O(N__54823),
            .I(N__54814));
    Odrv4 I__10553 (
            .O(N__54820),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__10552 (
            .O(N__54817),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__10551 (
            .O(N__54814),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    InMux I__10550 (
            .O(N__54807),
            .I(N__54801));
    InMux I__10549 (
            .O(N__54806),
            .I(N__54801));
    LocalMux I__10548 (
            .O(N__54801),
            .I(N__54798));
    Odrv4 I__10547 (
            .O(N__54798),
            .I(\pid_side.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__10546 (
            .O(N__54795),
            .I(N__54792));
    InMux I__10545 (
            .O(N__54792),
            .I(N__54788));
    InMux I__10544 (
            .O(N__54791),
            .I(N__54785));
    LocalMux I__10543 (
            .O(N__54788),
            .I(N__54782));
    LocalMux I__10542 (
            .O(N__54785),
            .I(\pid_side.error_i_acumm16lto3 ));
    Odrv4 I__10541 (
            .O(N__54782),
            .I(\pid_side.error_i_acumm16lto3 ));
    InMux I__10540 (
            .O(N__54777),
            .I(N__54771));
    InMux I__10539 (
            .O(N__54776),
            .I(N__54771));
    LocalMux I__10538 (
            .O(N__54771),
            .I(\pid_side.error_i_acumm_preregZ0Z_2 ));
    InMux I__10537 (
            .O(N__54768),
            .I(N__54765));
    LocalMux I__10536 (
            .O(N__54765),
            .I(\pid_side.un10lt9_1 ));
    CascadeMux I__10535 (
            .O(N__54762),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    InMux I__10534 (
            .O(N__54759),
            .I(N__54756));
    LocalMux I__10533 (
            .O(N__54756),
            .I(N__54753));
    Span4Mux_v I__10532 (
            .O(N__54753),
            .I(N__54750));
    Odrv4 I__10531 (
            .O(N__54750),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__10530 (
            .O(N__54747),
            .I(N__54738));
    InMux I__10529 (
            .O(N__54746),
            .I(N__54738));
    InMux I__10528 (
            .O(N__54745),
            .I(N__54738));
    LocalMux I__10527 (
            .O(N__54738),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    CascadeMux I__10526 (
            .O(N__54735),
            .I(N__54732));
    InMux I__10525 (
            .O(N__54732),
            .I(N__54729));
    LocalMux I__10524 (
            .O(N__54729),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__10523 (
            .O(N__54726),
            .I(N__54723));
    LocalMux I__10522 (
            .O(N__54723),
            .I(N__54720));
    Span4Mux_v I__10521 (
            .O(N__54720),
            .I(N__54716));
    InMux I__10520 (
            .O(N__54719),
            .I(N__54713));
    Span4Mux_h I__10519 (
            .O(N__54716),
            .I(N__54708));
    LocalMux I__10518 (
            .O(N__54713),
            .I(N__54708));
    Odrv4 I__10517 (
            .O(N__54708),
            .I(front_order_12));
    CascadeMux I__10516 (
            .O(N__54705),
            .I(N__54700));
    InMux I__10515 (
            .O(N__54704),
            .I(N__54693));
    InMux I__10514 (
            .O(N__54703),
            .I(N__54693));
    InMux I__10513 (
            .O(N__54700),
            .I(N__54693));
    LocalMux I__10512 (
            .O(N__54693),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__10511 (
            .O(N__54690),
            .I(N__54687));
    LocalMux I__10510 (
            .O(N__54687),
            .I(N__54683));
    InMux I__10509 (
            .O(N__54686),
            .I(N__54680));
    Span4Mux_v I__10508 (
            .O(N__54683),
            .I(N__54675));
    LocalMux I__10507 (
            .O(N__54680),
            .I(N__54675));
    Span4Mux_h I__10506 (
            .O(N__54675),
            .I(N__54672));
    Span4Mux_h I__10505 (
            .O(N__54672),
            .I(N__54669));
    Odrv4 I__10504 (
            .O(N__54669),
            .I(throttle_order_12));
    InMux I__10503 (
            .O(N__54666),
            .I(N__54663));
    LocalMux I__10502 (
            .O(N__54663),
            .I(N__54660));
    Span4Mux_v I__10501 (
            .O(N__54660),
            .I(N__54657));
    Odrv4 I__10500 (
            .O(N__54657),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    CascadeMux I__10499 (
            .O(N__54654),
            .I(N__54649));
    InMux I__10498 (
            .O(N__54653),
            .I(N__54642));
    InMux I__10497 (
            .O(N__54652),
            .I(N__54642));
    InMux I__10496 (
            .O(N__54649),
            .I(N__54642));
    LocalMux I__10495 (
            .O(N__54642),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    CascadeMux I__10494 (
            .O(N__54639),
            .I(\pid_side.un1_reset_0_i_cascade_ ));
    CascadeMux I__10493 (
            .O(N__54636),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ));
    InMux I__10492 (
            .O(N__54633),
            .I(N__54628));
    InMux I__10491 (
            .O(N__54632),
            .I(N__54625));
    InMux I__10490 (
            .O(N__54631),
            .I(N__54622));
    LocalMux I__10489 (
            .O(N__54628),
            .I(N__54619));
    LocalMux I__10488 (
            .O(N__54625),
            .I(N__54616));
    LocalMux I__10487 (
            .O(N__54622),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv12 I__10486 (
            .O(N__54619),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv12 I__10485 (
            .O(N__54616),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__10484 (
            .O(N__54609),
            .I(N__54606));
    LocalMux I__10483 (
            .O(N__54606),
            .I(N__54603));
    Span4Mux_v I__10482 (
            .O(N__54603),
            .I(N__54600));
    Odrv4 I__10481 (
            .O(N__54600),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__10480 (
            .O(N__54597),
            .I(N__54594));
    InMux I__10479 (
            .O(N__54594),
            .I(N__54591));
    LocalMux I__10478 (
            .O(N__54591),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__10477 (
            .O(N__54588),
            .I(N__54583));
    InMux I__10476 (
            .O(N__54587),
            .I(N__54580));
    InMux I__10475 (
            .O(N__54586),
            .I(N__54577));
    LocalMux I__10474 (
            .O(N__54583),
            .I(N__54574));
    LocalMux I__10473 (
            .O(N__54580),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__10472 (
            .O(N__54577),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv12 I__10471 (
            .O(N__54574),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    CascadeMux I__10470 (
            .O(N__54567),
            .I(\ppm_encoder_1.N_295_cascade_ ));
    InMux I__10469 (
            .O(N__54564),
            .I(N__54561));
    LocalMux I__10468 (
            .O(N__54561),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ));
    CascadeMux I__10467 (
            .O(N__54558),
            .I(N__54554));
    CascadeMux I__10466 (
            .O(N__54557),
            .I(N__54550));
    InMux I__10465 (
            .O(N__54554),
            .I(N__54547));
    InMux I__10464 (
            .O(N__54553),
            .I(N__54542));
    InMux I__10463 (
            .O(N__54550),
            .I(N__54542));
    LocalMux I__10462 (
            .O(N__54547),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__10461 (
            .O(N__54542),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__10460 (
            .O(N__54537),
            .I(N__54534));
    LocalMux I__10459 (
            .O(N__54534),
            .I(N__54530));
    InMux I__10458 (
            .O(N__54533),
            .I(N__54526));
    Span4Mux_h I__10457 (
            .O(N__54530),
            .I(N__54523));
    InMux I__10456 (
            .O(N__54529),
            .I(N__54520));
    LocalMux I__10455 (
            .O(N__54526),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__10454 (
            .O(N__54523),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    LocalMux I__10453 (
            .O(N__54520),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__10452 (
            .O(N__54513),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    InMux I__10451 (
            .O(N__54510),
            .I(N__54507));
    LocalMux I__10450 (
            .O(N__54507),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    CascadeMux I__10449 (
            .O(N__54504),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ));
    InMux I__10448 (
            .O(N__54501),
            .I(N__54498));
    LocalMux I__10447 (
            .O(N__54498),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8 ));
    CascadeMux I__10446 (
            .O(N__54495),
            .I(\ppm_encoder_1.N_294_cascade_ ));
    InMux I__10445 (
            .O(N__54492),
            .I(N__54489));
    LocalMux I__10444 (
            .O(N__54489),
            .I(N__54486));
    Span4Mux_h I__10443 (
            .O(N__54486),
            .I(N__54483));
    Odrv4 I__10442 (
            .O(N__54483),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ));
    InMux I__10441 (
            .O(N__54480),
            .I(N__54471));
    InMux I__10440 (
            .O(N__54479),
            .I(N__54471));
    InMux I__10439 (
            .O(N__54478),
            .I(N__54471));
    LocalMux I__10438 (
            .O(N__54471),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__10437 (
            .O(N__54468),
            .I(N__54465));
    InMux I__10436 (
            .O(N__54465),
            .I(N__54462));
    LocalMux I__10435 (
            .O(N__54462),
            .I(N__54459));
    Odrv4 I__10434 (
            .O(N__54459),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__10433 (
            .O(N__54456),
            .I(N__54453));
    LocalMux I__10432 (
            .O(N__54453),
            .I(N__54449));
    InMux I__10431 (
            .O(N__54452),
            .I(N__54446));
    Span4Mux_v I__10430 (
            .O(N__54449),
            .I(N__54441));
    LocalMux I__10429 (
            .O(N__54446),
            .I(N__54441));
    Odrv4 I__10428 (
            .O(N__54441),
            .I(front_order_8));
    CascadeMux I__10427 (
            .O(N__54438),
            .I(N__54433));
    InMux I__10426 (
            .O(N__54437),
            .I(N__54426));
    InMux I__10425 (
            .O(N__54436),
            .I(N__54426));
    InMux I__10424 (
            .O(N__54433),
            .I(N__54426));
    LocalMux I__10423 (
            .O(N__54426),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__10422 (
            .O(N__54423),
            .I(N__54420));
    LocalMux I__10421 (
            .O(N__54420),
            .I(N__54417));
    Span4Mux_v I__10420 (
            .O(N__54417),
            .I(N__54414));
    Odrv4 I__10419 (
            .O(N__54414),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__10418 (
            .O(N__54411),
            .I(N__54408));
    LocalMux I__10417 (
            .O(N__54408),
            .I(N__54404));
    CascadeMux I__10416 (
            .O(N__54407),
            .I(N__54400));
    Span4Mux_v I__10415 (
            .O(N__54404),
            .I(N__54397));
    InMux I__10414 (
            .O(N__54403),
            .I(N__54394));
    InMux I__10413 (
            .O(N__54400),
            .I(N__54391));
    Sp12to4 I__10412 (
            .O(N__54397),
            .I(N__54386));
    LocalMux I__10411 (
            .O(N__54394),
            .I(N__54386));
    LocalMux I__10410 (
            .O(N__54391),
            .I(throttle_order_8));
    Odrv12 I__10409 (
            .O(N__54386),
            .I(throttle_order_8));
    CascadeMux I__10408 (
            .O(N__54381),
            .I(N__54376));
    InMux I__10407 (
            .O(N__54380),
            .I(N__54369));
    InMux I__10406 (
            .O(N__54379),
            .I(N__54369));
    InMux I__10405 (
            .O(N__54376),
            .I(N__54369));
    LocalMux I__10404 (
            .O(N__54369),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    CascadeMux I__10403 (
            .O(N__54366),
            .I(\ppm_encoder_1.PPM_STATE_53_d_cascade_ ));
    CascadeMux I__10402 (
            .O(N__54363),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6_cascade_ ));
    CascadeMux I__10401 (
            .O(N__54360),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ));
    CascadeMux I__10400 (
            .O(N__54357),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ));
    CascadeMux I__10399 (
            .O(N__54354),
            .I(N__54351));
    InMux I__10398 (
            .O(N__54351),
            .I(N__54345));
    InMux I__10397 (
            .O(N__54350),
            .I(N__54345));
    LocalMux I__10396 (
            .O(N__54345),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    InMux I__10395 (
            .O(N__54342),
            .I(N__54338));
    InMux I__10394 (
            .O(N__54341),
            .I(N__54335));
    LocalMux I__10393 (
            .O(N__54338),
            .I(N__54332));
    LocalMux I__10392 (
            .O(N__54335),
            .I(N__54329));
    Span4Mux_v I__10391 (
            .O(N__54332),
            .I(N__54326));
    Span4Mux_h I__10390 (
            .O(N__54329),
            .I(N__54323));
    Odrv4 I__10389 (
            .O(N__54326),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv4 I__10388 (
            .O(N__54323),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    CascadeMux I__10387 (
            .O(N__54318),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    CascadeMux I__10386 (
            .O(N__54315),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ));
    CascadeMux I__10385 (
            .O(N__54312),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ));
    CascadeMux I__10384 (
            .O(N__54309),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ));
    InMux I__10383 (
            .O(N__54306),
            .I(N__54300));
    InMux I__10382 (
            .O(N__54305),
            .I(N__54300));
    LocalMux I__10381 (
            .O(N__54300),
            .I(N__54297));
    Span4Mux_v I__10380 (
            .O(N__54297),
            .I(N__54294));
    Odrv4 I__10379 (
            .O(N__54294),
            .I(\ppm_encoder_1.N_232 ));
    InMux I__10378 (
            .O(N__54291),
            .I(N__54288));
    LocalMux I__10377 (
            .O(N__54288),
            .I(N__54285));
    Span4Mux_h I__10376 (
            .O(N__54285),
            .I(N__54282));
    Odrv4 I__10375 (
            .O(N__54282),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__10374 (
            .O(N__54279),
            .I(N__54276));
    LocalMux I__10373 (
            .O(N__54276),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__10372 (
            .O(N__54273),
            .I(N__54270));
    LocalMux I__10371 (
            .O(N__54270),
            .I(N__54267));
    Span4Mux_v I__10370 (
            .O(N__54267),
            .I(N__54264));
    Odrv4 I__10369 (
            .O(N__54264),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__10368 (
            .O(N__54261),
            .I(N__54258));
    LocalMux I__10367 (
            .O(N__54258),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    CascadeMux I__10366 (
            .O(N__54255),
            .I(N__54252));
    InMux I__10365 (
            .O(N__54252),
            .I(N__54249));
    LocalMux I__10364 (
            .O(N__54249),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__10363 (
            .O(N__54246),
            .I(N__54241));
    InMux I__10362 (
            .O(N__54245),
            .I(N__54238));
    InMux I__10361 (
            .O(N__54244),
            .I(N__54235));
    LocalMux I__10360 (
            .O(N__54241),
            .I(N__54232));
    LocalMux I__10359 (
            .O(N__54238),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__10358 (
            .O(N__54235),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__10357 (
            .O(N__54232),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__10356 (
            .O(N__54225),
            .I(N__54222));
    LocalMux I__10355 (
            .O(N__54222),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    CascadeMux I__10354 (
            .O(N__54219),
            .I(N__54216));
    InMux I__10353 (
            .O(N__54216),
            .I(N__54213));
    LocalMux I__10352 (
            .O(N__54213),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__10351 (
            .O(N__54210),
            .I(N__54205));
    InMux I__10350 (
            .O(N__54209),
            .I(N__54202));
    InMux I__10349 (
            .O(N__54208),
            .I(N__54199));
    LocalMux I__10348 (
            .O(N__54205),
            .I(N__54196));
    LocalMux I__10347 (
            .O(N__54202),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__10346 (
            .O(N__54199),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__10345 (
            .O(N__54196),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    CascadeMux I__10344 (
            .O(N__54189),
            .I(N__54184));
    InMux I__10343 (
            .O(N__54188),
            .I(N__54181));
    CascadeMux I__10342 (
            .O(N__54187),
            .I(N__54178));
    InMux I__10341 (
            .O(N__54184),
            .I(N__54175));
    LocalMux I__10340 (
            .O(N__54181),
            .I(N__54172));
    InMux I__10339 (
            .O(N__54178),
            .I(N__54169));
    LocalMux I__10338 (
            .O(N__54175),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv4 I__10337 (
            .O(N__54172),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    LocalMux I__10336 (
            .O(N__54169),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__10335 (
            .O(N__54162),
            .I(N__54157));
    InMux I__10334 (
            .O(N__54161),
            .I(N__54154));
    CascadeMux I__10333 (
            .O(N__54160),
            .I(N__54151));
    LocalMux I__10332 (
            .O(N__54157),
            .I(N__54148));
    LocalMux I__10331 (
            .O(N__54154),
            .I(N__54145));
    InMux I__10330 (
            .O(N__54151),
            .I(N__54142));
    Odrv4 I__10329 (
            .O(N__54148),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    Odrv4 I__10328 (
            .O(N__54145),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    LocalMux I__10327 (
            .O(N__54142),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__10326 (
            .O(N__54135),
            .I(N__54132));
    LocalMux I__10325 (
            .O(N__54132),
            .I(N__54129));
    Span4Mux_v I__10324 (
            .O(N__54129),
            .I(N__54126));
    Odrv4 I__10323 (
            .O(N__54126),
            .I(\ppm_encoder_1.N_293 ));
    InMux I__10322 (
            .O(N__54123),
            .I(N__54120));
    LocalMux I__10321 (
            .O(N__54120),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    CascadeMux I__10320 (
            .O(N__54117),
            .I(\ppm_encoder_1.N_314_cascade_ ));
    InMux I__10319 (
            .O(N__54114),
            .I(N__54111));
    LocalMux I__10318 (
            .O(N__54111),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    CascadeMux I__10317 (
            .O(N__54108),
            .I(N__54104));
    CascadeMux I__10316 (
            .O(N__54107),
            .I(N__54100));
    InMux I__10315 (
            .O(N__54104),
            .I(N__54097));
    InMux I__10314 (
            .O(N__54103),
            .I(N__54094));
    InMux I__10313 (
            .O(N__54100),
            .I(N__54091));
    LocalMux I__10312 (
            .O(N__54097),
            .I(N__54088));
    LocalMux I__10311 (
            .O(N__54094),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__10310 (
            .O(N__54091),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__10309 (
            .O(N__54088),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__10308 (
            .O(N__54081),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__10307 (
            .O(N__54078),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__10306 (
            .O(N__54075),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__10305 (
            .O(N__54072),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__10304 (
            .O(N__54069),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__10303 (
            .O(N__54066),
            .I(bfn_14_4_0_));
    InMux I__10302 (
            .O(N__54063),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__10301 (
            .O(N__54060),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__10300 (
            .O(N__54057),
            .I(N__54054));
    LocalMux I__10299 (
            .O(N__54054),
            .I(N__54050));
    SRMux I__10298 (
            .O(N__54053),
            .I(N__54047));
    Span4Mux_v I__10297 (
            .O(N__54050),
            .I(N__54042));
    LocalMux I__10296 (
            .O(N__54047),
            .I(N__54042));
    Span4Mux_s2_v I__10295 (
            .O(N__54042),
            .I(N__54038));
    SRMux I__10294 (
            .O(N__54041),
            .I(N__54035));
    Sp12to4 I__10293 (
            .O(N__54038),
            .I(N__54030));
    LocalMux I__10292 (
            .O(N__54035),
            .I(N__54030));
    Odrv12 I__10291 (
            .O(N__54030),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__10290 (
            .O(N__54027),
            .I(N__54022));
    InMux I__10289 (
            .O(N__54026),
            .I(N__54019));
    InMux I__10288 (
            .O(N__54025),
            .I(N__54016));
    LocalMux I__10287 (
            .O(N__54022),
            .I(N__54013));
    LocalMux I__10286 (
            .O(N__54019),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__10285 (
            .O(N__54016),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__10284 (
            .O(N__54013),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    CascadeMux I__10283 (
            .O(N__54006),
            .I(N__54001));
    InMux I__10282 (
            .O(N__54005),
            .I(N__53998));
    InMux I__10281 (
            .O(N__54004),
            .I(N__53995));
    InMux I__10280 (
            .O(N__54001),
            .I(N__53992));
    LocalMux I__10279 (
            .O(N__53998),
            .I(N__53989));
    LocalMux I__10278 (
            .O(N__53995),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__10277 (
            .O(N__53992),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__10276 (
            .O(N__53989),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__10275 (
            .O(N__53982),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__10274 (
            .O(N__53979),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__10273 (
            .O(N__53976),
            .I(N__53971));
    InMux I__10272 (
            .O(N__53975),
            .I(N__53968));
    InMux I__10271 (
            .O(N__53974),
            .I(N__53965));
    LocalMux I__10270 (
            .O(N__53971),
            .I(N__53962));
    LocalMux I__10269 (
            .O(N__53968),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__10268 (
            .O(N__53965),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__10267 (
            .O(N__53962),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__10266 (
            .O(N__53955),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__10265 (
            .O(N__53952),
            .I(N__53949));
    LocalMux I__10264 (
            .O(N__53949),
            .I(N__53944));
    InMux I__10263 (
            .O(N__53948),
            .I(N__53941));
    InMux I__10262 (
            .O(N__53947),
            .I(N__53938));
    Span4Mux_h I__10261 (
            .O(N__53944),
            .I(N__53935));
    LocalMux I__10260 (
            .O(N__53941),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__10259 (
            .O(N__53938),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    Odrv4 I__10258 (
            .O(N__53935),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__10257 (
            .O(N__53928),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__10256 (
            .O(N__53925),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__10255 (
            .O(N__53922),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__10254 (
            .O(N__53919),
            .I(bfn_14_3_0_));
    InMux I__10253 (
            .O(N__53916),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__10252 (
            .O(N__53913),
            .I(N__53908));
    InMux I__10251 (
            .O(N__53912),
            .I(N__53905));
    InMux I__10250 (
            .O(N__53911),
            .I(N__53902));
    LocalMux I__10249 (
            .O(N__53908),
            .I(N__53899));
    LocalMux I__10248 (
            .O(N__53905),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__10247 (
            .O(N__53902),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__10246 (
            .O(N__53899),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__10245 (
            .O(N__53892),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__10244 (
            .O(N__53889),
            .I(N__53886));
    LocalMux I__10243 (
            .O(N__53886),
            .I(N__53882));
    InMux I__10242 (
            .O(N__53885),
            .I(N__53879));
    Span12Mux_v I__10241 (
            .O(N__53882),
            .I(N__53876));
    LocalMux I__10240 (
            .O(N__53879),
            .I(N__53873));
    Span12Mux_h I__10239 (
            .O(N__53876),
            .I(N__53867));
    Span12Mux_s1_h I__10238 (
            .O(N__53873),
            .I(N__53867));
    InMux I__10237 (
            .O(N__53872),
            .I(N__53861));
    Span12Mux_h I__10236 (
            .O(N__53867),
            .I(N__53858));
    InMux I__10235 (
            .O(N__53866),
            .I(N__53855));
    InMux I__10234 (
            .O(N__53865),
            .I(N__53852));
    InMux I__10233 (
            .O(N__53864),
            .I(N__53849));
    LocalMux I__10232 (
            .O(N__53861),
            .I(N__53846));
    Odrv12 I__10231 (
            .O(N__53858),
            .I(\pid_front.error_9 ));
    LocalMux I__10230 (
            .O(N__53855),
            .I(\pid_front.error_9 ));
    LocalMux I__10229 (
            .O(N__53852),
            .I(\pid_front.error_9 ));
    LocalMux I__10228 (
            .O(N__53849),
            .I(\pid_front.error_9 ));
    Odrv4 I__10227 (
            .O(N__53846),
            .I(\pid_front.error_9 ));
    InMux I__10226 (
            .O(N__53835),
            .I(N__53832));
    LocalMux I__10225 (
            .O(N__53832),
            .I(N__53828));
    InMux I__10224 (
            .O(N__53831),
            .I(N__53825));
    Span4Mux_v I__10223 (
            .O(N__53828),
            .I(N__53821));
    LocalMux I__10222 (
            .O(N__53825),
            .I(N__53818));
    InMux I__10221 (
            .O(N__53824),
            .I(N__53815));
    Span4Mux_h I__10220 (
            .O(N__53821),
            .I(N__53812));
    Span12Mux_v I__10219 (
            .O(N__53818),
            .I(N__53808));
    LocalMux I__10218 (
            .O(N__53815),
            .I(N__53805));
    Span4Mux_h I__10217 (
            .O(N__53812),
            .I(N__53799));
    InMux I__10216 (
            .O(N__53811),
            .I(N__53796));
    Span12Mux_h I__10215 (
            .O(N__53808),
            .I(N__53793));
    Span4Mux_v I__10214 (
            .O(N__53805),
            .I(N__53790));
    InMux I__10213 (
            .O(N__53804),
            .I(N__53787));
    InMux I__10212 (
            .O(N__53803),
            .I(N__53782));
    InMux I__10211 (
            .O(N__53802),
            .I(N__53782));
    Span4Mux_h I__10210 (
            .O(N__53799),
            .I(N__53777));
    LocalMux I__10209 (
            .O(N__53796),
            .I(N__53777));
    Odrv12 I__10208 (
            .O(N__53793),
            .I(\pid_front.error_10 ));
    Odrv4 I__10207 (
            .O(N__53790),
            .I(\pid_front.error_10 ));
    LocalMux I__10206 (
            .O(N__53787),
            .I(\pid_front.error_10 ));
    LocalMux I__10205 (
            .O(N__53782),
            .I(\pid_front.error_10 ));
    Odrv4 I__10204 (
            .O(N__53777),
            .I(\pid_front.error_10 ));
    CascadeMux I__10203 (
            .O(N__53766),
            .I(\pid_front.N_21_1_cascade_ ));
    InMux I__10202 (
            .O(N__53763),
            .I(N__53758));
    InMux I__10201 (
            .O(N__53762),
            .I(N__53753));
    InMux I__10200 (
            .O(N__53761),
            .I(N__53753));
    LocalMux I__10199 (
            .O(N__53758),
            .I(\pid_front.N_21_1 ));
    LocalMux I__10198 (
            .O(N__53753),
            .I(\pid_front.N_21_1 ));
    InMux I__10197 (
            .O(N__53748),
            .I(N__53742));
    InMux I__10196 (
            .O(N__53747),
            .I(N__53742));
    LocalMux I__10195 (
            .O(N__53742),
            .I(\pid_front.N_25_0 ));
    InMux I__10194 (
            .O(N__53739),
            .I(N__53736));
    LocalMux I__10193 (
            .O(N__53736),
            .I(\pid_front.m38_1_ns_1 ));
    CascadeMux I__10192 (
            .O(N__53733),
            .I(\pid_front.N_39_1_cascade_ ));
    InMux I__10191 (
            .O(N__53730),
            .I(N__53727));
    LocalMux I__10190 (
            .O(N__53727),
            .I(N__53724));
    Odrv4 I__10189 (
            .O(N__53724),
            .I(\pid_front.error_i_reg_9_rn_1_18 ));
    CascadeMux I__10188 (
            .O(N__53721),
            .I(N__53718));
    InMux I__10187 (
            .O(N__53718),
            .I(N__53715));
    LocalMux I__10186 (
            .O(N__53715),
            .I(N__53712));
    Span4Mux_h I__10185 (
            .O(N__53712),
            .I(N__53709));
    Span4Mux_v I__10184 (
            .O(N__53709),
            .I(N__53706));
    Odrv4 I__10183 (
            .O(N__53706),
            .I(\pid_front.error_i_regZ0Z_18 ));
    InMux I__10182 (
            .O(N__53703),
            .I(N__53700));
    LocalMux I__10181 (
            .O(N__53700),
            .I(\pid_front.error_i_reg_9_rn_1_26 ));
    InMux I__10180 (
            .O(N__53697),
            .I(N__53693));
    InMux I__10179 (
            .O(N__53696),
            .I(N__53690));
    LocalMux I__10178 (
            .O(N__53693),
            .I(\pid_front.N_39_1 ));
    LocalMux I__10177 (
            .O(N__53690),
            .I(\pid_front.N_39_1 ));
    CascadeMux I__10176 (
            .O(N__53685),
            .I(N__53682));
    InMux I__10175 (
            .O(N__53682),
            .I(N__53679));
    LocalMux I__10174 (
            .O(N__53679),
            .I(N__53676));
    Span4Mux_h I__10173 (
            .O(N__53676),
            .I(N__53673));
    Span4Mux_v I__10172 (
            .O(N__53673),
            .I(N__53670));
    Odrv4 I__10171 (
            .O(N__53670),
            .I(\pid_front.error_i_regZ0Z_26 ));
    InMux I__10170 (
            .O(N__53667),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    CascadeMux I__10169 (
            .O(N__53664),
            .I(\pid_front.error_i_reg_esr_RNO_1_0_24_cascade_ ));
    CascadeMux I__10168 (
            .O(N__53661),
            .I(N__53658));
    InMux I__10167 (
            .O(N__53658),
            .I(N__53655));
    LocalMux I__10166 (
            .O(N__53655),
            .I(N__53652));
    Span4Mux_h I__10165 (
            .O(N__53652),
            .I(N__53649));
    Odrv4 I__10164 (
            .O(N__53649),
            .I(\pid_front.error_i_regZ0Z_24 ));
    InMux I__10163 (
            .O(N__53646),
            .I(N__53643));
    LocalMux I__10162 (
            .O(N__53643),
            .I(\pid_front.error_cry_7_c_RNI1ADUZ0Z1 ));
    InMux I__10161 (
            .O(N__53640),
            .I(N__53637));
    LocalMux I__10160 (
            .O(N__53637),
            .I(\pid_front.error_cry_7_c_RNI1ADU1Z0Z_0 ));
    CascadeMux I__10159 (
            .O(N__53634),
            .I(\pid_front.N_22_0_cascade_ ));
    InMux I__10158 (
            .O(N__53631),
            .I(N__53628));
    LocalMux I__10157 (
            .O(N__53628),
            .I(\pid_front.N_27_1 ));
    CascadeMux I__10156 (
            .O(N__53625),
            .I(\pid_front.error_cry_2_0_c_RNI198HZ0Z2_cascade_ ));
    InMux I__10155 (
            .O(N__53622),
            .I(N__53619));
    LocalMux I__10154 (
            .O(N__53619),
            .I(\pid_front.error_cry_2_0_c_RNI198H2Z0Z_0 ));
    InMux I__10153 (
            .O(N__53616),
            .I(N__53613));
    LocalMux I__10152 (
            .O(N__53613),
            .I(N__53609));
    InMux I__10151 (
            .O(N__53612),
            .I(N__53606));
    Odrv4 I__10150 (
            .O(N__53609),
            .I(\pid_front.N_28_1 ));
    LocalMux I__10149 (
            .O(N__53606),
            .I(\pid_front.N_28_1 ));
    CascadeMux I__10148 (
            .O(N__53601),
            .I(\pid_front.N_28_1_cascade_ ));
    InMux I__10147 (
            .O(N__53598),
            .I(N__53594));
    InMux I__10146 (
            .O(N__53597),
            .I(N__53591));
    LocalMux I__10145 (
            .O(N__53594),
            .I(N__53588));
    LocalMux I__10144 (
            .O(N__53591),
            .I(N__53585));
    Span4Mux_h I__10143 (
            .O(N__53588),
            .I(N__53582));
    Span4Mux_v I__10142 (
            .O(N__53585),
            .I(N__53579));
    Span4Mux_v I__10141 (
            .O(N__53582),
            .I(N__53576));
    Span4Mux_h I__10140 (
            .O(N__53579),
            .I(N__53573));
    Span4Mux_h I__10139 (
            .O(N__53576),
            .I(N__53569));
    Span4Mux_h I__10138 (
            .O(N__53573),
            .I(N__53563));
    InMux I__10137 (
            .O(N__53572),
            .I(N__53560));
    Span4Mux_h I__10136 (
            .O(N__53569),
            .I(N__53555));
    InMux I__10135 (
            .O(N__53568),
            .I(N__53552));
    InMux I__10134 (
            .O(N__53567),
            .I(N__53549));
    InMux I__10133 (
            .O(N__53566),
            .I(N__53546));
    Span4Mux_h I__10132 (
            .O(N__53563),
            .I(N__53541));
    LocalMux I__10131 (
            .O(N__53560),
            .I(N__53541));
    InMux I__10130 (
            .O(N__53559),
            .I(N__53536));
    InMux I__10129 (
            .O(N__53558),
            .I(N__53536));
    Odrv4 I__10128 (
            .O(N__53555),
            .I(\pid_front.error_8 ));
    LocalMux I__10127 (
            .O(N__53552),
            .I(\pid_front.error_8 ));
    LocalMux I__10126 (
            .O(N__53549),
            .I(\pid_front.error_8 ));
    LocalMux I__10125 (
            .O(N__53546),
            .I(\pid_front.error_8 ));
    Odrv4 I__10124 (
            .O(N__53541),
            .I(\pid_front.error_8 ));
    LocalMux I__10123 (
            .O(N__53536),
            .I(\pid_front.error_8 ));
    InMux I__10122 (
            .O(N__53523),
            .I(N__53520));
    LocalMux I__10121 (
            .O(N__53520),
            .I(N__53516));
    InMux I__10120 (
            .O(N__53519),
            .I(N__53512));
    Span4Mux_v I__10119 (
            .O(N__53516),
            .I(N__53509));
    CascadeMux I__10118 (
            .O(N__53515),
            .I(N__53504));
    LocalMux I__10117 (
            .O(N__53512),
            .I(N__53500));
    Span4Mux_h I__10116 (
            .O(N__53509),
            .I(N__53497));
    InMux I__10115 (
            .O(N__53508),
            .I(N__53494));
    InMux I__10114 (
            .O(N__53507),
            .I(N__53489));
    InMux I__10113 (
            .O(N__53504),
            .I(N__53484));
    InMux I__10112 (
            .O(N__53503),
            .I(N__53484));
    Span12Mux_s7_v I__10111 (
            .O(N__53500),
            .I(N__53481));
    Span4Mux_h I__10110 (
            .O(N__53497),
            .I(N__53478));
    LocalMux I__10109 (
            .O(N__53494),
            .I(N__53475));
    InMux I__10108 (
            .O(N__53493),
            .I(N__53470));
    InMux I__10107 (
            .O(N__53492),
            .I(N__53470));
    LocalMux I__10106 (
            .O(N__53489),
            .I(N__53465));
    LocalMux I__10105 (
            .O(N__53484),
            .I(N__53465));
    Span12Mux_h I__10104 (
            .O(N__53481),
            .I(N__53462));
    Span4Mux_h I__10103 (
            .O(N__53478),
            .I(N__53459));
    Odrv4 I__10102 (
            .O(N__53475),
            .I(\pid_front.error_7 ));
    LocalMux I__10101 (
            .O(N__53470),
            .I(\pid_front.error_7 ));
    Odrv4 I__10100 (
            .O(N__53465),
            .I(\pid_front.error_7 ));
    Odrv12 I__10099 (
            .O(N__53462),
            .I(\pid_front.error_7 ));
    Odrv4 I__10098 (
            .O(N__53459),
            .I(\pid_front.error_7 ));
    CascadeMux I__10097 (
            .O(N__53448),
            .I(\pid_front.N_25_0_cascade_ ));
    CascadeMux I__10096 (
            .O(N__53445),
            .I(N__53442));
    InMux I__10095 (
            .O(N__53442),
            .I(N__53439));
    LocalMux I__10094 (
            .O(N__53439),
            .I(N__53434));
    InMux I__10093 (
            .O(N__53438),
            .I(N__53429));
    InMux I__10092 (
            .O(N__53437),
            .I(N__53429));
    Odrv4 I__10091 (
            .O(N__53434),
            .I(drone_H_disp_front_13));
    LocalMux I__10090 (
            .O(N__53429),
            .I(drone_H_disp_front_13));
    InMux I__10089 (
            .O(N__53424),
            .I(N__53421));
    LocalMux I__10088 (
            .O(N__53421),
            .I(drone_H_disp_front_i_13));
    InMux I__10087 (
            .O(N__53418),
            .I(N__53412));
    InMux I__10086 (
            .O(N__53417),
            .I(N__53412));
    LocalMux I__10085 (
            .O(N__53412),
            .I(\dron_frame_decoder_1.drone_H_disp_front_5 ));
    InMux I__10084 (
            .O(N__53409),
            .I(N__53406));
    LocalMux I__10083 (
            .O(N__53406),
            .I(drone_H_disp_front_i_5));
    InMux I__10082 (
            .O(N__53403),
            .I(N__53397));
    InMux I__10081 (
            .O(N__53402),
            .I(N__53397));
    LocalMux I__10080 (
            .O(N__53397),
            .I(\dron_frame_decoder_1.drone_H_disp_front_6 ));
    InMux I__10079 (
            .O(N__53394),
            .I(N__53391));
    LocalMux I__10078 (
            .O(N__53391),
            .I(drone_H_disp_front_i_6));
    CascadeMux I__10077 (
            .O(N__53388),
            .I(N__53384));
    InMux I__10076 (
            .O(N__53387),
            .I(N__53378));
    InMux I__10075 (
            .O(N__53384),
            .I(N__53378));
    InMux I__10074 (
            .O(N__53383),
            .I(N__53375));
    LocalMux I__10073 (
            .O(N__53378),
            .I(N__53372));
    LocalMux I__10072 (
            .O(N__53375),
            .I(drone_H_disp_front_14));
    Odrv4 I__10071 (
            .O(N__53372),
            .I(drone_H_disp_front_14));
    InMux I__10070 (
            .O(N__53367),
            .I(N__53364));
    LocalMux I__10069 (
            .O(N__53364),
            .I(N__53361));
    Span4Mux_h I__10068 (
            .O(N__53361),
            .I(N__53356));
    CascadeMux I__10067 (
            .O(N__53360),
            .I(N__53352));
    InMux I__10066 (
            .O(N__53359),
            .I(N__53349));
    Sp12to4 I__10065 (
            .O(N__53356),
            .I(N__53346));
    InMux I__10064 (
            .O(N__53355),
            .I(N__53341));
    InMux I__10063 (
            .O(N__53352),
            .I(N__53341));
    LocalMux I__10062 (
            .O(N__53349),
            .I(N__53338));
    Span12Mux_v I__10061 (
            .O(N__53346),
            .I(N__53335));
    LocalMux I__10060 (
            .O(N__53341),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    Odrv4 I__10059 (
            .O(N__53338),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    Odrv12 I__10058 (
            .O(N__53335),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    CascadeMux I__10057 (
            .O(N__53328),
            .I(N__53322));
    CascadeMux I__10056 (
            .O(N__53327),
            .I(N__53319));
    CascadeMux I__10055 (
            .O(N__53326),
            .I(N__53316));
    CascadeMux I__10054 (
            .O(N__53325),
            .I(N__53312));
    InMux I__10053 (
            .O(N__53322),
            .I(N__53295));
    InMux I__10052 (
            .O(N__53319),
            .I(N__53295));
    InMux I__10051 (
            .O(N__53316),
            .I(N__53295));
    InMux I__10050 (
            .O(N__53315),
            .I(N__53292));
    InMux I__10049 (
            .O(N__53312),
            .I(N__53285));
    InMux I__10048 (
            .O(N__53311),
            .I(N__53285));
    InMux I__10047 (
            .O(N__53310),
            .I(N__53285));
    InMux I__10046 (
            .O(N__53309),
            .I(N__53278));
    InMux I__10045 (
            .O(N__53308),
            .I(N__53278));
    InMux I__10044 (
            .O(N__53307),
            .I(N__53278));
    InMux I__10043 (
            .O(N__53306),
            .I(N__53271));
    InMux I__10042 (
            .O(N__53305),
            .I(N__53271));
    InMux I__10041 (
            .O(N__53304),
            .I(N__53271));
    InMux I__10040 (
            .O(N__53303),
            .I(N__53266));
    InMux I__10039 (
            .O(N__53302),
            .I(N__53266));
    LocalMux I__10038 (
            .O(N__53295),
            .I(N__53262));
    LocalMux I__10037 (
            .O(N__53292),
            .I(N__53257));
    LocalMux I__10036 (
            .O(N__53285),
            .I(N__53257));
    LocalMux I__10035 (
            .O(N__53278),
            .I(N__53252));
    LocalMux I__10034 (
            .O(N__53271),
            .I(N__53252));
    LocalMux I__10033 (
            .O(N__53266),
            .I(N__53249));
    CascadeMux I__10032 (
            .O(N__53265),
            .I(N__53246));
    Span4Mux_v I__10031 (
            .O(N__53262),
            .I(N__53241));
    Span4Mux_v I__10030 (
            .O(N__53257),
            .I(N__53241));
    Span4Mux_v I__10029 (
            .O(N__53252),
            .I(N__53236));
    Span4Mux_v I__10028 (
            .O(N__53249),
            .I(N__53236));
    InMux I__10027 (
            .O(N__53246),
            .I(N__53231));
    Sp12to4 I__10026 (
            .O(N__53241),
            .I(N__53226));
    Sp12to4 I__10025 (
            .O(N__53236),
            .I(N__53226));
    InMux I__10024 (
            .O(N__53235),
            .I(N__53221));
    InMux I__10023 (
            .O(N__53234),
            .I(N__53221));
    LocalMux I__10022 (
            .O(N__53231),
            .I(N__53216));
    Span12Mux_h I__10021 (
            .O(N__53226),
            .I(N__53216));
    LocalMux I__10020 (
            .O(N__53221),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    Odrv12 I__10019 (
            .O(N__53216),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__10018 (
            .O(N__53211),
            .I(N__53205));
    CascadeMux I__10017 (
            .O(N__53210),
            .I(N__53202));
    CascadeMux I__10016 (
            .O(N__53209),
            .I(N__53197));
    CascadeMux I__10015 (
            .O(N__53208),
            .I(N__53193));
    InMux I__10014 (
            .O(N__53205),
            .I(N__53184));
    InMux I__10013 (
            .O(N__53202),
            .I(N__53184));
    InMux I__10012 (
            .O(N__53201),
            .I(N__53184));
    InMux I__10011 (
            .O(N__53200),
            .I(N__53184));
    InMux I__10010 (
            .O(N__53197),
            .I(N__53177));
    InMux I__10009 (
            .O(N__53196),
            .I(N__53177));
    InMux I__10008 (
            .O(N__53193),
            .I(N__53177));
    LocalMux I__10007 (
            .O(N__53184),
            .I(N__53168));
    LocalMux I__10006 (
            .O(N__53177),
            .I(N__53168));
    CascadeMux I__10005 (
            .O(N__53176),
            .I(N__53165));
    CascadeMux I__10004 (
            .O(N__53175),
            .I(N__53162));
    CascadeMux I__10003 (
            .O(N__53174),
            .I(N__53159));
    CascadeMux I__10002 (
            .O(N__53173),
            .I(N__53156));
    Span4Mux_v I__10001 (
            .O(N__53168),
            .I(N__53153));
    InMux I__10000 (
            .O(N__53165),
            .I(N__53144));
    InMux I__9999 (
            .O(N__53162),
            .I(N__53144));
    InMux I__9998 (
            .O(N__53159),
            .I(N__53144));
    InMux I__9997 (
            .O(N__53156),
            .I(N__53144));
    Odrv4 I__9996 (
            .O(N__53153),
            .I(\dron_frame_decoder_1.N_122_mux_i ));
    LocalMux I__9995 (
            .O(N__53144),
            .I(\dron_frame_decoder_1.N_122_mux_i ));
    InMux I__9994 (
            .O(N__53139),
            .I(N__53133));
    InMux I__9993 (
            .O(N__53138),
            .I(N__53133));
    LocalMux I__9992 (
            .O(N__53133),
            .I(\dron_frame_decoder_1.drone_H_disp_front_10 ));
    InMux I__9991 (
            .O(N__53130),
            .I(N__53127));
    LocalMux I__9990 (
            .O(N__53127),
            .I(N__53124));
    Odrv4 I__9989 (
            .O(N__53124),
            .I(drone_H_disp_front_i_10));
    CascadeMux I__9988 (
            .O(N__53121),
            .I(\pid_front.error_cry_5_c_RNIUOTVZ0Z1_cascade_ ));
    InMux I__9987 (
            .O(N__53118),
            .I(N__53115));
    LocalMux I__9986 (
            .O(N__53115),
            .I(\pid_front.error_cry_5_c_RNIUOTV1Z0Z_0 ));
    InMux I__9985 (
            .O(N__53112),
            .I(N__53105));
    InMux I__9984 (
            .O(N__53111),
            .I(N__53105));
    InMux I__9983 (
            .O(N__53110),
            .I(N__53102));
    LocalMux I__9982 (
            .O(N__53105),
            .I(N__53099));
    LocalMux I__9981 (
            .O(N__53102),
            .I(N__53096));
    Span4Mux_h I__9980 (
            .O(N__53099),
            .I(N__53093));
    Odrv4 I__9979 (
            .O(N__53096),
            .I(\pid_front.N_49_0 ));
    Odrv4 I__9978 (
            .O(N__53093),
            .I(\pid_front.N_49_0 ));
    CascadeMux I__9977 (
            .O(N__53088),
            .I(\pid_front.N_49_0_cascade_ ));
    InMux I__9976 (
            .O(N__53085),
            .I(N__53082));
    LocalMux I__9975 (
            .O(N__53082),
            .I(N__53077));
    InMux I__9974 (
            .O(N__53081),
            .I(N__53074));
    InMux I__9973 (
            .O(N__53080),
            .I(N__53071));
    Odrv4 I__9972 (
            .O(N__53077),
            .I(\pid_front.N_46_1 ));
    LocalMux I__9971 (
            .O(N__53074),
            .I(\pid_front.N_46_1 ));
    LocalMux I__9970 (
            .O(N__53071),
            .I(\pid_front.N_46_1 ));
    CascadeMux I__9969 (
            .O(N__53064),
            .I(\pid_front.m134_0_ns_1_cascade_ ));
    CascadeMux I__9968 (
            .O(N__53061),
            .I(\pid_front.m19_2_03_0_cascade_ ));
    CascadeMux I__9967 (
            .O(N__53058),
            .I(N__53055));
    InMux I__9966 (
            .O(N__53055),
            .I(N__53052));
    LocalMux I__9965 (
            .O(N__53052),
            .I(N__53049));
    Span4Mux_h I__9964 (
            .O(N__53049),
            .I(N__53046));
    Odrv4 I__9963 (
            .O(N__53046),
            .I(\pid_front.error_i_regZ0Z_15 ));
    InMux I__9962 (
            .O(N__53043),
            .I(N__53040));
    LocalMux I__9961 (
            .O(N__53040),
            .I(N__53037));
    Span4Mux_h I__9960 (
            .O(N__53037),
            .I(N__53033));
    InMux I__9959 (
            .O(N__53036),
            .I(N__53030));
    Odrv4 I__9958 (
            .O(N__53033),
            .I(\pid_front.N_48_1 ));
    LocalMux I__9957 (
            .O(N__53030),
            .I(\pid_front.N_48_1 ));
    InMux I__9956 (
            .O(N__53025),
            .I(N__53022));
    LocalMux I__9955 (
            .O(N__53022),
            .I(N__53019));
    Span4Mux_v I__9954 (
            .O(N__53019),
            .I(N__53016));
    Span4Mux_h I__9953 (
            .O(N__53016),
            .I(N__53013));
    Span4Mux_h I__9952 (
            .O(N__53013),
            .I(N__53010));
    Odrv4 I__9951 (
            .O(N__53010),
            .I(\pid_front.O_3 ));
    InMux I__9950 (
            .O(N__53007),
            .I(N__53001));
    InMux I__9949 (
            .O(N__53006),
            .I(N__53001));
    LocalMux I__9948 (
            .O(N__53001),
            .I(N__52994));
    InMux I__9947 (
            .O(N__53000),
            .I(N__52991));
    InMux I__9946 (
            .O(N__52999),
            .I(N__52984));
    InMux I__9945 (
            .O(N__52998),
            .I(N__52984));
    InMux I__9944 (
            .O(N__52997),
            .I(N__52984));
    Odrv4 I__9943 (
            .O(N__52994),
            .I(\pid_front.error_d_regZ0Z_1 ));
    LocalMux I__9942 (
            .O(N__52991),
            .I(\pid_front.error_d_regZ0Z_1 ));
    LocalMux I__9941 (
            .O(N__52984),
            .I(\pid_front.error_d_regZ0Z_1 ));
    InMux I__9940 (
            .O(N__52977),
            .I(N__52973));
    CascadeMux I__9939 (
            .O(N__52976),
            .I(N__52970));
    LocalMux I__9938 (
            .O(N__52973),
            .I(N__52967));
    InMux I__9937 (
            .O(N__52970),
            .I(N__52964));
    Span4Mux_v I__9936 (
            .O(N__52967),
            .I(N__52961));
    LocalMux I__9935 (
            .O(N__52964),
            .I(N__52958));
    Span4Mux_h I__9934 (
            .O(N__52961),
            .I(N__52955));
    Span4Mux_h I__9933 (
            .O(N__52958),
            .I(N__52952));
    Odrv4 I__9932 (
            .O(N__52955),
            .I(\pid_front.un1_pid_prereg_0 ));
    Odrv4 I__9931 (
            .O(N__52952),
            .I(\pid_front.un1_pid_prereg_0 ));
    InMux I__9930 (
            .O(N__52947),
            .I(N__52939));
    InMux I__9929 (
            .O(N__52946),
            .I(N__52939));
    InMux I__9928 (
            .O(N__52945),
            .I(N__52934));
    InMux I__9927 (
            .O(N__52944),
            .I(N__52934));
    LocalMux I__9926 (
            .O(N__52939),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    LocalMux I__9925 (
            .O(N__52934),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    InMux I__9924 (
            .O(N__52929),
            .I(N__52926));
    LocalMux I__9923 (
            .O(N__52926),
            .I(N__52923));
    Span4Mux_h I__9922 (
            .O(N__52923),
            .I(N__52920));
    Span4Mux_v I__9921 (
            .O(N__52920),
            .I(N__52917));
    Odrv4 I__9920 (
            .O(N__52917),
            .I(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ));
    InMux I__9919 (
            .O(N__52914),
            .I(N__52911));
    LocalMux I__9918 (
            .O(N__52911),
            .I(N__52908));
    Span12Mux_h I__9917 (
            .O(N__52908),
            .I(N__52905));
    Odrv12 I__9916 (
            .O(N__52905),
            .I(\pid_front.O_2 ));
    InMux I__9915 (
            .O(N__52902),
            .I(N__52893));
    InMux I__9914 (
            .O(N__52901),
            .I(N__52893));
    InMux I__9913 (
            .O(N__52900),
            .I(N__52886));
    InMux I__9912 (
            .O(N__52899),
            .I(N__52886));
    InMux I__9911 (
            .O(N__52898),
            .I(N__52886));
    LocalMux I__9910 (
            .O(N__52893),
            .I(\pid_front.error_d_regZ0Z_0 ));
    LocalMux I__9909 (
            .O(N__52886),
            .I(\pid_front.error_d_regZ0Z_0 ));
    InMux I__9908 (
            .O(N__52881),
            .I(N__52877));
    InMux I__9907 (
            .O(N__52880),
            .I(N__52874));
    LocalMux I__9906 (
            .O(N__52877),
            .I(N__52868));
    LocalMux I__9905 (
            .O(N__52874),
            .I(N__52868));
    InMux I__9904 (
            .O(N__52873),
            .I(N__52865));
    Span12Mux_h I__9903 (
            .O(N__52868),
            .I(N__52862));
    LocalMux I__9902 (
            .O(N__52865),
            .I(drone_altitude_15));
    Odrv12 I__9901 (
            .O(N__52862),
            .I(drone_altitude_15));
    InMux I__9900 (
            .O(N__52857),
            .I(N__52841));
    InMux I__9899 (
            .O(N__52856),
            .I(N__52841));
    InMux I__9898 (
            .O(N__52855),
            .I(N__52841));
    InMux I__9897 (
            .O(N__52854),
            .I(N__52841));
    InMux I__9896 (
            .O(N__52853),
            .I(N__52830));
    InMux I__9895 (
            .O(N__52852),
            .I(N__52830));
    InMux I__9894 (
            .O(N__52851),
            .I(N__52830));
    InMux I__9893 (
            .O(N__52850),
            .I(N__52830));
    LocalMux I__9892 (
            .O(N__52841),
            .I(N__52827));
    InMux I__9891 (
            .O(N__52840),
            .I(N__52819));
    InMux I__9890 (
            .O(N__52839),
            .I(N__52819));
    LocalMux I__9889 (
            .O(N__52830),
            .I(N__52814));
    Span4Mux_v I__9888 (
            .O(N__52827),
            .I(N__52814));
    InMux I__9887 (
            .O(N__52826),
            .I(N__52809));
    InMux I__9886 (
            .O(N__52825),
            .I(N__52809));
    CascadeMux I__9885 (
            .O(N__52824),
            .I(N__52806));
    LocalMux I__9884 (
            .O(N__52819),
            .I(N__52800));
    Span4Mux_s3_h I__9883 (
            .O(N__52814),
            .I(N__52795));
    LocalMux I__9882 (
            .O(N__52809),
            .I(N__52795));
    InMux I__9881 (
            .O(N__52806),
            .I(N__52786));
    InMux I__9880 (
            .O(N__52805),
            .I(N__52786));
    InMux I__9879 (
            .O(N__52804),
            .I(N__52786));
    InMux I__9878 (
            .O(N__52803),
            .I(N__52786));
    Span12Mux_h I__9877 (
            .O(N__52800),
            .I(N__52783));
    Span4Mux_h I__9876 (
            .O(N__52795),
            .I(N__52780));
    LocalMux I__9875 (
            .O(N__52786),
            .I(N__52777));
    Odrv12 I__9874 (
            .O(N__52783),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_0 ));
    Odrv4 I__9873 (
            .O(N__52780),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_0 ));
    Odrv12 I__9872 (
            .O(N__52777),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_0 ));
    InMux I__9871 (
            .O(N__52770),
            .I(N__52767));
    LocalMux I__9870 (
            .O(N__52767),
            .I(N__52764));
    Span4Mux_v I__9869 (
            .O(N__52764),
            .I(N__52761));
    Sp12to4 I__9868 (
            .O(N__52761),
            .I(N__52758));
    Span12Mux_h I__9867 (
            .O(N__52758),
            .I(N__52753));
    InMux I__9866 (
            .O(N__52757),
            .I(N__52748));
    InMux I__9865 (
            .O(N__52756),
            .I(N__52748));
    Odrv12 I__9864 (
            .O(N__52753),
            .I(drone_altitude_7));
    LocalMux I__9863 (
            .O(N__52748),
            .I(drone_altitude_7));
    InMux I__9862 (
            .O(N__52743),
            .I(N__52740));
    LocalMux I__9861 (
            .O(N__52740),
            .I(N__52737));
    Span12Mux_v I__9860 (
            .O(N__52737),
            .I(N__52734));
    Span12Mux_h I__9859 (
            .O(N__52734),
            .I(N__52731));
    Odrv12 I__9858 (
            .O(N__52731),
            .I(drone_altitude_i_7));
    InMux I__9857 (
            .O(N__52728),
            .I(N__52724));
    CascadeMux I__9856 (
            .O(N__52727),
            .I(N__52721));
    LocalMux I__9855 (
            .O(N__52724),
            .I(N__52718));
    InMux I__9854 (
            .O(N__52721),
            .I(N__52715));
    Span4Mux_v I__9853 (
            .O(N__52718),
            .I(N__52712));
    LocalMux I__9852 (
            .O(N__52715),
            .I(drone_H_disp_front_15));
    Odrv4 I__9851 (
            .O(N__52712),
            .I(drone_H_disp_front_15));
    InMux I__9850 (
            .O(N__52707),
            .I(N__52701));
    InMux I__9849 (
            .O(N__52706),
            .I(N__52701));
    LocalMux I__9848 (
            .O(N__52701),
            .I(\dron_frame_decoder_1.drone_H_disp_front_7 ));
    InMux I__9847 (
            .O(N__52698),
            .I(N__52695));
    LocalMux I__9846 (
            .O(N__52695),
            .I(drone_H_disp_front_i_7));
    InMux I__9845 (
            .O(N__52692),
            .I(N__52689));
    LocalMux I__9844 (
            .O(N__52689),
            .I(N__52686));
    Span4Mux_v I__9843 (
            .O(N__52686),
            .I(N__52682));
    InMux I__9842 (
            .O(N__52685),
            .I(N__52679));
    Span4Mux_h I__9841 (
            .O(N__52682),
            .I(N__52676));
    LocalMux I__9840 (
            .O(N__52679),
            .I(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ));
    Odrv4 I__9839 (
            .O(N__52676),
            .I(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ));
    InMux I__9838 (
            .O(N__52671),
            .I(N__52665));
    InMux I__9837 (
            .O(N__52670),
            .I(N__52665));
    LocalMux I__9836 (
            .O(N__52665),
            .I(N__52662));
    Span4Mux_h I__9835 (
            .O(N__52662),
            .I(N__52659));
    Span4Mux_h I__9834 (
            .O(N__52659),
            .I(N__52656));
    Span4Mux_h I__9833 (
            .O(N__52656),
            .I(N__52653));
    Odrv4 I__9832 (
            .O(N__52653),
            .I(\pid_front.error_p_regZ0Z_16 ));
    InMux I__9831 (
            .O(N__52650),
            .I(N__52644));
    InMux I__9830 (
            .O(N__52649),
            .I(N__52644));
    LocalMux I__9829 (
            .O(N__52644),
            .I(\pid_front.error_d_reg_prevZ0Z_16 ));
    InMux I__9828 (
            .O(N__52641),
            .I(N__52635));
    InMux I__9827 (
            .O(N__52640),
            .I(N__52635));
    LocalMux I__9826 (
            .O(N__52635),
            .I(N__52632));
    Span4Mux_h I__9825 (
            .O(N__52632),
            .I(N__52629));
    Odrv4 I__9824 (
            .O(N__52629),
            .I(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ));
    InMux I__9823 (
            .O(N__52626),
            .I(N__52623));
    LocalMux I__9822 (
            .O(N__52623),
            .I(N__52619));
    InMux I__9821 (
            .O(N__52622),
            .I(N__52616));
    Span4Mux_v I__9820 (
            .O(N__52619),
            .I(N__52611));
    LocalMux I__9819 (
            .O(N__52616),
            .I(N__52611));
    Span4Mux_h I__9818 (
            .O(N__52611),
            .I(N__52608));
    Span4Mux_h I__9817 (
            .O(N__52608),
            .I(N__52605));
    Span4Mux_v I__9816 (
            .O(N__52605),
            .I(N__52602));
    Odrv4 I__9815 (
            .O(N__52602),
            .I(\pid_front.error_p_regZ0Z_18 ));
    InMux I__9814 (
            .O(N__52599),
            .I(N__52596));
    LocalMux I__9813 (
            .O(N__52596),
            .I(N__52592));
    InMux I__9812 (
            .O(N__52595),
            .I(N__52589));
    Odrv4 I__9811 (
            .O(N__52592),
            .I(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ));
    LocalMux I__9810 (
            .O(N__52589),
            .I(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ));
    InMux I__9809 (
            .O(N__52584),
            .I(N__52580));
    InMux I__9808 (
            .O(N__52583),
            .I(N__52577));
    LocalMux I__9807 (
            .O(N__52580),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    LocalMux I__9806 (
            .O(N__52577),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    CEMux I__9805 (
            .O(N__52572),
            .I(N__52566));
    CEMux I__9804 (
            .O(N__52571),
            .I(N__52563));
    CEMux I__9803 (
            .O(N__52570),
            .I(N__52560));
    CEMux I__9802 (
            .O(N__52569),
            .I(N__52555));
    LocalMux I__9801 (
            .O(N__52566),
            .I(N__52552));
    LocalMux I__9800 (
            .O(N__52563),
            .I(N__52547));
    LocalMux I__9799 (
            .O(N__52560),
            .I(N__52547));
    CEMux I__9798 (
            .O(N__52559),
            .I(N__52544));
    CEMux I__9797 (
            .O(N__52558),
            .I(N__52537));
    LocalMux I__9796 (
            .O(N__52555),
            .I(N__52528));
    Span4Mux_v I__9795 (
            .O(N__52552),
            .I(N__52528));
    Span4Mux_v I__9794 (
            .O(N__52547),
            .I(N__52528));
    LocalMux I__9793 (
            .O(N__52544),
            .I(N__52528));
    CEMux I__9792 (
            .O(N__52543),
            .I(N__52524));
    CEMux I__9791 (
            .O(N__52542),
            .I(N__52521));
    CEMux I__9790 (
            .O(N__52541),
            .I(N__52518));
    CEMux I__9789 (
            .O(N__52540),
            .I(N__52515));
    LocalMux I__9788 (
            .O(N__52537),
            .I(N__52510));
    Span4Mux_v I__9787 (
            .O(N__52528),
            .I(N__52510));
    CEMux I__9786 (
            .O(N__52527),
            .I(N__52507));
    LocalMux I__9785 (
            .O(N__52524),
            .I(N__52504));
    LocalMux I__9784 (
            .O(N__52521),
            .I(N__52501));
    LocalMux I__9783 (
            .O(N__52518),
            .I(N__52498));
    LocalMux I__9782 (
            .O(N__52515),
            .I(N__52495));
    Span4Mux_v I__9781 (
            .O(N__52510),
            .I(N__52492));
    LocalMux I__9780 (
            .O(N__52507),
            .I(N__52489));
    Span4Mux_h I__9779 (
            .O(N__52504),
            .I(N__52486));
    Span4Mux_v I__9778 (
            .O(N__52501),
            .I(N__52483));
    Span4Mux_h I__9777 (
            .O(N__52498),
            .I(N__52476));
    Span4Mux_v I__9776 (
            .O(N__52495),
            .I(N__52476));
    Span4Mux_h I__9775 (
            .O(N__52492),
            .I(N__52476));
    Odrv12 I__9774 (
            .O(N__52489),
            .I(\pid_front.N_404_0 ));
    Odrv4 I__9773 (
            .O(N__52486),
            .I(\pid_front.N_404_0 ));
    Odrv4 I__9772 (
            .O(N__52483),
            .I(\pid_front.N_404_0 ));
    Odrv4 I__9771 (
            .O(N__52476),
            .I(\pid_front.N_404_0 ));
    SRMux I__9770 (
            .O(N__52467),
            .I(N__52462));
    SRMux I__9769 (
            .O(N__52466),
            .I(N__52458));
    SRMux I__9768 (
            .O(N__52465),
            .I(N__52455));
    LocalMux I__9767 (
            .O(N__52462),
            .I(N__52452));
    SRMux I__9766 (
            .O(N__52461),
            .I(N__52449));
    LocalMux I__9765 (
            .O(N__52458),
            .I(N__52441));
    LocalMux I__9764 (
            .O(N__52455),
            .I(N__52438));
    Span4Mux_v I__9763 (
            .O(N__52452),
            .I(N__52433));
    LocalMux I__9762 (
            .O(N__52449),
            .I(N__52433));
    SRMux I__9761 (
            .O(N__52448),
            .I(N__52430));
    SRMux I__9760 (
            .O(N__52447),
            .I(N__52425));
    SRMux I__9759 (
            .O(N__52446),
            .I(N__52422));
    SRMux I__9758 (
            .O(N__52445),
            .I(N__52419));
    SRMux I__9757 (
            .O(N__52444),
            .I(N__52416));
    Span4Mux_v I__9756 (
            .O(N__52441),
            .I(N__52411));
    Span4Mux_h I__9755 (
            .O(N__52438),
            .I(N__52411));
    Span4Mux_h I__9754 (
            .O(N__52433),
            .I(N__52406));
    LocalMux I__9753 (
            .O(N__52430),
            .I(N__52406));
    SRMux I__9752 (
            .O(N__52429),
            .I(N__52403));
    SRMux I__9751 (
            .O(N__52428),
            .I(N__52400));
    LocalMux I__9750 (
            .O(N__52425),
            .I(N__52397));
    LocalMux I__9749 (
            .O(N__52422),
            .I(N__52394));
    LocalMux I__9748 (
            .O(N__52419),
            .I(N__52391));
    LocalMux I__9747 (
            .O(N__52416),
            .I(N__52388));
    Span4Mux_h I__9746 (
            .O(N__52411),
            .I(N__52379));
    Span4Mux_h I__9745 (
            .O(N__52406),
            .I(N__52379));
    LocalMux I__9744 (
            .O(N__52403),
            .I(N__52379));
    LocalMux I__9743 (
            .O(N__52400),
            .I(N__52379));
    Span4Mux_h I__9742 (
            .O(N__52397),
            .I(N__52375));
    Span4Mux_v I__9741 (
            .O(N__52394),
            .I(N__52370));
    Span4Mux_h I__9740 (
            .O(N__52391),
            .I(N__52370));
    Span4Mux_h I__9739 (
            .O(N__52388),
            .I(N__52367));
    Span4Mux_v I__9738 (
            .O(N__52379),
            .I(N__52364));
    InMux I__9737 (
            .O(N__52378),
            .I(N__52361));
    Span4Mux_h I__9736 (
            .O(N__52375),
            .I(N__52358));
    Span4Mux_h I__9735 (
            .O(N__52370),
            .I(N__52355));
    Span4Mux_h I__9734 (
            .O(N__52367),
            .I(N__52352));
    Span4Mux_h I__9733 (
            .O(N__52364),
            .I(N__52347));
    LocalMux I__9732 (
            .O(N__52361),
            .I(N__52347));
    Odrv4 I__9731 (
            .O(N__52358),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    Odrv4 I__9730 (
            .O(N__52355),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    Odrv4 I__9729 (
            .O(N__52352),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    Odrv4 I__9728 (
            .O(N__52347),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    InMux I__9727 (
            .O(N__52338),
            .I(N__52335));
    LocalMux I__9726 (
            .O(N__52335),
            .I(N__52332));
    Span4Mux_v I__9725 (
            .O(N__52332),
            .I(N__52329));
    Sp12to4 I__9724 (
            .O(N__52329),
            .I(N__52326));
    Span12Mux_h I__9723 (
            .O(N__52326),
            .I(N__52323));
    Odrv12 I__9722 (
            .O(N__52323),
            .I(\pid_front.O_0_4 ));
    CascadeMux I__9721 (
            .O(N__52320),
            .I(N__52316));
    InMux I__9720 (
            .O(N__52319),
            .I(N__52311));
    InMux I__9719 (
            .O(N__52316),
            .I(N__52304));
    InMux I__9718 (
            .O(N__52315),
            .I(N__52304));
    InMux I__9717 (
            .O(N__52314),
            .I(N__52304));
    LocalMux I__9716 (
            .O(N__52311),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    LocalMux I__9715 (
            .O(N__52304),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__9714 (
            .O(N__52299),
            .I(N__52294));
    CascadeMux I__9713 (
            .O(N__52298),
            .I(N__52291));
    InMux I__9712 (
            .O(N__52297),
            .I(N__52288));
    InMux I__9711 (
            .O(N__52294),
            .I(N__52283));
    InMux I__9710 (
            .O(N__52291),
            .I(N__52283));
    LocalMux I__9709 (
            .O(N__52288),
            .I(\pid_front.error_p_regZ0Z_1 ));
    LocalMux I__9708 (
            .O(N__52283),
            .I(\pid_front.error_p_regZ0Z_1 ));
    InMux I__9707 (
            .O(N__52278),
            .I(N__52274));
    CascadeMux I__9706 (
            .O(N__52277),
            .I(N__52270));
    LocalMux I__9705 (
            .O(N__52274),
            .I(N__52267));
    InMux I__9704 (
            .O(N__52273),
            .I(N__52264));
    InMux I__9703 (
            .O(N__52270),
            .I(N__52261));
    Span4Mux_v I__9702 (
            .O(N__52267),
            .I(N__52258));
    LocalMux I__9701 (
            .O(N__52264),
            .I(N__52255));
    LocalMux I__9700 (
            .O(N__52261),
            .I(N__52252));
    Span4Mux_h I__9699 (
            .O(N__52258),
            .I(N__52247));
    Span4Mux_h I__9698 (
            .O(N__52255),
            .I(N__52247));
    Span4Mux_h I__9697 (
            .O(N__52252),
            .I(N__52244));
    Odrv4 I__9696 (
            .O(N__52247),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    Odrv4 I__9695 (
            .O(N__52244),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    CascadeMux I__9694 (
            .O(N__52239),
            .I(\pid_front.un1_pid_prereg_9_0_cascade_ ));
    InMux I__9693 (
            .O(N__52236),
            .I(N__52233));
    LocalMux I__9692 (
            .O(N__52233),
            .I(N__52230));
    Span4Mux_v I__9691 (
            .O(N__52230),
            .I(N__52227));
    Span4Mux_v I__9690 (
            .O(N__52227),
            .I(N__52224));
    Odrv4 I__9689 (
            .O(N__52224),
            .I(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ));
    InMux I__9688 (
            .O(N__52221),
            .I(N__52218));
    LocalMux I__9687 (
            .O(N__52218),
            .I(pid_side_m153_e_5));
    CascadeMux I__9686 (
            .O(N__52215),
            .I(pid_side_m153_e_5_cascade_));
    CascadeMux I__9685 (
            .O(N__52212),
            .I(\pid_side.N_196_mux_cascade_ ));
    CascadeMux I__9684 (
            .O(N__52209),
            .I(N__52206));
    InMux I__9683 (
            .O(N__52206),
            .I(N__52200));
    InMux I__9682 (
            .O(N__52205),
            .I(N__52200));
    LocalMux I__9681 (
            .O(N__52200),
            .I(pid_side_m153_e_4));
    InMux I__9680 (
            .O(N__52197),
            .I(N__52186));
    InMux I__9679 (
            .O(N__52196),
            .I(N__52186));
    InMux I__9678 (
            .O(N__52195),
            .I(N__52186));
    InMux I__9677 (
            .O(N__52194),
            .I(N__52179));
    InMux I__9676 (
            .O(N__52193),
            .I(N__52179));
    LocalMux I__9675 (
            .O(N__52186),
            .I(N__52176));
    InMux I__9674 (
            .O(N__52185),
            .I(N__52173));
    CascadeMux I__9673 (
            .O(N__52184),
            .I(N__52170));
    LocalMux I__9672 (
            .O(N__52179),
            .I(N__52166));
    Span4Mux_v I__9671 (
            .O(N__52176),
            .I(N__52163));
    LocalMux I__9670 (
            .O(N__52173),
            .I(N__52160));
    InMux I__9669 (
            .O(N__52170),
            .I(N__52155));
    InMux I__9668 (
            .O(N__52169),
            .I(N__52155));
    Span4Mux_h I__9667 (
            .O(N__52166),
            .I(N__52152));
    Span4Mux_h I__9666 (
            .O(N__52163),
            .I(N__52149));
    Span12Mux_s8_v I__9665 (
            .O(N__52160),
            .I(N__52146));
    LocalMux I__9664 (
            .O(N__52155),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__9663 (
            .O(N__52152),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__9662 (
            .O(N__52149),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv12 I__9661 (
            .O(N__52146),
            .I(\pid_front.stateZ0Z_0 ));
    InMux I__9660 (
            .O(N__52137),
            .I(N__52127));
    InMux I__9659 (
            .O(N__52136),
            .I(N__52111));
    InMux I__9658 (
            .O(N__52135),
            .I(N__52111));
    InMux I__9657 (
            .O(N__52134),
            .I(N__52111));
    InMux I__9656 (
            .O(N__52133),
            .I(N__52111));
    InMux I__9655 (
            .O(N__52132),
            .I(N__52111));
    InMux I__9654 (
            .O(N__52131),
            .I(N__52111));
    InMux I__9653 (
            .O(N__52130),
            .I(N__52111));
    LocalMux I__9652 (
            .O(N__52127),
            .I(N__52106));
    CascadeMux I__9651 (
            .O(N__52126),
            .I(N__52101));
    LocalMux I__9650 (
            .O(N__52111),
            .I(N__52098));
    InMux I__9649 (
            .O(N__52110),
            .I(N__52095));
    InMux I__9648 (
            .O(N__52109),
            .I(N__52092));
    Span4Mux_v I__9647 (
            .O(N__52106),
            .I(N__52089));
    InMux I__9646 (
            .O(N__52105),
            .I(N__52082));
    InMux I__9645 (
            .O(N__52104),
            .I(N__52082));
    InMux I__9644 (
            .O(N__52101),
            .I(N__52082));
    Span4Mux_h I__9643 (
            .O(N__52098),
            .I(N__52077));
    LocalMux I__9642 (
            .O(N__52095),
            .I(N__52072));
    LocalMux I__9641 (
            .O(N__52092),
            .I(N__52072));
    Span4Mux_h I__9640 (
            .O(N__52089),
            .I(N__52067));
    LocalMux I__9639 (
            .O(N__52082),
            .I(N__52067));
    InMux I__9638 (
            .O(N__52081),
            .I(N__52062));
    InMux I__9637 (
            .O(N__52080),
            .I(N__52062));
    Span4Mux_v I__9636 (
            .O(N__52077),
            .I(N__52057));
    Span4Mux_h I__9635 (
            .O(N__52072),
            .I(N__52057));
    Span4Mux_v I__9634 (
            .O(N__52067),
            .I(N__52054));
    LocalMux I__9633 (
            .O(N__52062),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__9632 (
            .O(N__52057),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__9631 (
            .O(N__52054),
            .I(\pid_front.stateZ0Z_1 ));
    InMux I__9630 (
            .O(N__52047),
            .I(N__52044));
    LocalMux I__9629 (
            .O(N__52044),
            .I(N__52041));
    Span4Mux_h I__9628 (
            .O(N__52041),
            .I(N__52038));
    Span4Mux_h I__9627 (
            .O(N__52038),
            .I(N__52035));
    Odrv4 I__9626 (
            .O(N__52035),
            .I(\pid_front.state_RNIVIRQZ0Z_0 ));
    InMux I__9625 (
            .O(N__52032),
            .I(N__52026));
    InMux I__9624 (
            .O(N__52031),
            .I(N__52026));
    LocalMux I__9623 (
            .O(N__52026),
            .I(N__52023));
    Odrv4 I__9622 (
            .O(N__52023),
            .I(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ));
    InMux I__9621 (
            .O(N__52020),
            .I(N__52014));
    InMux I__9620 (
            .O(N__52019),
            .I(N__52014));
    LocalMux I__9619 (
            .O(N__52014),
            .I(N__52011));
    Span4Mux_h I__9618 (
            .O(N__52011),
            .I(N__52008));
    Span4Mux_h I__9617 (
            .O(N__52008),
            .I(N__52005));
    Span4Mux_h I__9616 (
            .O(N__52005),
            .I(N__52002));
    Odrv4 I__9615 (
            .O(N__52002),
            .I(\pid_front.error_p_regZ0Z_15 ));
    InMux I__9614 (
            .O(N__51999),
            .I(N__51993));
    InMux I__9613 (
            .O(N__51998),
            .I(N__51993));
    LocalMux I__9612 (
            .O(N__51993),
            .I(\pid_front.error_d_reg_prevZ0Z_15 ));
    InMux I__9611 (
            .O(N__51990),
            .I(N__51987));
    LocalMux I__9610 (
            .O(N__51987),
            .I(N__51983));
    InMux I__9609 (
            .O(N__51986),
            .I(N__51980));
    Span4Mux_v I__9608 (
            .O(N__51983),
            .I(N__51977));
    LocalMux I__9607 (
            .O(N__51980),
            .I(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ));
    Odrv4 I__9606 (
            .O(N__51977),
            .I(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ));
    CascadeMux I__9605 (
            .O(N__51972),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ));
    InMux I__9604 (
            .O(N__51969),
            .I(N__51965));
    InMux I__9603 (
            .O(N__51968),
            .I(N__51962));
    LocalMux I__9602 (
            .O(N__51965),
            .I(\pid_front.error_d_reg_prev_esr_RNIKI4D7Z0Z_12 ));
    LocalMux I__9601 (
            .O(N__51962),
            .I(\pid_front.error_d_reg_prev_esr_RNIKI4D7Z0Z_12 ));
    CascadeMux I__9600 (
            .O(N__51957),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ));
    CascadeMux I__9599 (
            .O(N__51954),
            .I(N__51951));
    InMux I__9598 (
            .O(N__51951),
            .I(N__51948));
    LocalMux I__9597 (
            .O(N__51948),
            .I(N__51945));
    Span4Mux_h I__9596 (
            .O(N__51945),
            .I(N__51942));
    Odrv4 I__9595 (
            .O(N__51942),
            .I(\pid_front.error_p_reg_esr_RNIJ35VFZ0Z_12 ));
    InMux I__9594 (
            .O(N__51939),
            .I(N__51933));
    InMux I__9593 (
            .O(N__51938),
            .I(N__51933));
    LocalMux I__9592 (
            .O(N__51933),
            .I(N__51930));
    Odrv12 I__9591 (
            .O(N__51930),
            .I(\pid_front.error_p_reg_esr_RNIROQ33_0Z0Z_12 ));
    InMux I__9590 (
            .O(N__51927),
            .I(N__51922));
    InMux I__9589 (
            .O(N__51926),
            .I(N__51919));
    InMux I__9588 (
            .O(N__51925),
            .I(N__51916));
    LocalMux I__9587 (
            .O(N__51922),
            .I(N__51911));
    LocalMux I__9586 (
            .O(N__51919),
            .I(N__51911));
    LocalMux I__9585 (
            .O(N__51916),
            .I(N__51908));
    Span4Mux_h I__9584 (
            .O(N__51911),
            .I(N__51905));
    Odrv4 I__9583 (
            .O(N__51908),
            .I(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ));
    Odrv4 I__9582 (
            .O(N__51905),
            .I(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ));
    InMux I__9581 (
            .O(N__51900),
            .I(N__51896));
    CascadeMux I__9580 (
            .O(N__51899),
            .I(N__51893));
    LocalMux I__9579 (
            .O(N__51896),
            .I(N__51888));
    InMux I__9578 (
            .O(N__51893),
            .I(N__51883));
    InMux I__9577 (
            .O(N__51892),
            .I(N__51883));
    InMux I__9576 (
            .O(N__51891),
            .I(N__51880));
    Span4Mux_v I__9575 (
            .O(N__51888),
            .I(N__51875));
    LocalMux I__9574 (
            .O(N__51883),
            .I(N__51875));
    LocalMux I__9573 (
            .O(N__51880),
            .I(N__51872));
    Span4Mux_h I__9572 (
            .O(N__51875),
            .I(N__51869));
    Odrv4 I__9571 (
            .O(N__51872),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ));
    Odrv4 I__9570 (
            .O(N__51869),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ));
    CascadeMux I__9569 (
            .O(N__51864),
            .I(\pid_front.un1_pid_prereg_153_0_cascade_ ));
    InMux I__9568 (
            .O(N__51861),
            .I(N__51858));
    LocalMux I__9567 (
            .O(N__51858),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ));
    InMux I__9566 (
            .O(N__51855),
            .I(N__51852));
    LocalMux I__9565 (
            .O(N__51852),
            .I(N__51849));
    Span4Mux_h I__9564 (
            .O(N__51849),
            .I(N__51846));
    Odrv4 I__9563 (
            .O(N__51846),
            .I(\pid_front.error_d_reg_prev_esr_RNINH0UDZ0Z_10 ));
    InMux I__9562 (
            .O(N__51843),
            .I(N__51837));
    InMux I__9561 (
            .O(N__51842),
            .I(N__51837));
    LocalMux I__9560 (
            .O(N__51837),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ));
    CascadeMux I__9559 (
            .O(N__51834),
            .I(N__51829));
    InMux I__9558 (
            .O(N__51833),
            .I(N__51825));
    InMux I__9557 (
            .O(N__51832),
            .I(N__51818));
    InMux I__9556 (
            .O(N__51829),
            .I(N__51818));
    InMux I__9555 (
            .O(N__51828),
            .I(N__51818));
    LocalMux I__9554 (
            .O(N__51825),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    LocalMux I__9553 (
            .O(N__51818),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    InMux I__9552 (
            .O(N__51813),
            .I(N__51810));
    LocalMux I__9551 (
            .O(N__51810),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ));
    InMux I__9550 (
            .O(N__51807),
            .I(N__51802));
    InMux I__9549 (
            .O(N__51806),
            .I(N__51797));
    InMux I__9548 (
            .O(N__51805),
            .I(N__51797));
    LocalMux I__9547 (
            .O(N__51802),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    LocalMux I__9546 (
            .O(N__51797),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    CascadeMux I__9545 (
            .O(N__51792),
            .I(N__51789));
    InMux I__9544 (
            .O(N__51789),
            .I(N__51781));
    InMux I__9543 (
            .O(N__51788),
            .I(N__51781));
    InMux I__9542 (
            .O(N__51787),
            .I(N__51776));
    InMux I__9541 (
            .O(N__51786),
            .I(N__51776));
    LocalMux I__9540 (
            .O(N__51781),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    LocalMux I__9539 (
            .O(N__51776),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    InMux I__9538 (
            .O(N__51771),
            .I(N__51767));
    CascadeMux I__9537 (
            .O(N__51770),
            .I(N__51763));
    LocalMux I__9536 (
            .O(N__51767),
            .I(N__51760));
    InMux I__9535 (
            .O(N__51766),
            .I(N__51755));
    InMux I__9534 (
            .O(N__51763),
            .I(N__51755));
    Span4Mux_h I__9533 (
            .O(N__51760),
            .I(N__51752));
    LocalMux I__9532 (
            .O(N__51755),
            .I(N__51749));
    Odrv4 I__9531 (
            .O(N__51752),
            .I(\pid_front.error_p_regZ0Z_10 ));
    Odrv12 I__9530 (
            .O(N__51749),
            .I(\pid_front.error_p_regZ0Z_10 ));
    InMux I__9529 (
            .O(N__51744),
            .I(N__51741));
    LocalMux I__9528 (
            .O(N__51741),
            .I(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ));
    CascadeMux I__9527 (
            .O(N__51738),
            .I(\pid_front.N_196_mux_cascade_ ));
    InMux I__9526 (
            .O(N__51735),
            .I(N__51732));
    LocalMux I__9525 (
            .O(N__51732),
            .I(N__51729));
    Span4Mux_h I__9524 (
            .O(N__51729),
            .I(N__51726));
    Span4Mux_h I__9523 (
            .O(N__51726),
            .I(N__51722));
    InMux I__9522 (
            .O(N__51725),
            .I(N__51719));
    Odrv4 I__9521 (
            .O(N__51722),
            .I(\pid_front.error_i_acumm16lto3 ));
    LocalMux I__9520 (
            .O(N__51719),
            .I(\pid_front.error_i_acumm16lto3 ));
    InMux I__9519 (
            .O(N__51714),
            .I(N__51711));
    LocalMux I__9518 (
            .O(N__51711),
            .I(N__51708));
    Span4Mux_v I__9517 (
            .O(N__51708),
            .I(N__51693));
    InMux I__9516 (
            .O(N__51707),
            .I(N__51678));
    InMux I__9515 (
            .O(N__51706),
            .I(N__51678));
    InMux I__9514 (
            .O(N__51705),
            .I(N__51678));
    InMux I__9513 (
            .O(N__51704),
            .I(N__51678));
    InMux I__9512 (
            .O(N__51703),
            .I(N__51678));
    InMux I__9511 (
            .O(N__51702),
            .I(N__51678));
    InMux I__9510 (
            .O(N__51701),
            .I(N__51678));
    InMux I__9509 (
            .O(N__51700),
            .I(N__51667));
    InMux I__9508 (
            .O(N__51699),
            .I(N__51667));
    InMux I__9507 (
            .O(N__51698),
            .I(N__51667));
    InMux I__9506 (
            .O(N__51697),
            .I(N__51667));
    InMux I__9505 (
            .O(N__51696),
            .I(N__51667));
    Odrv4 I__9504 (
            .O(N__51693),
            .I(\pid_front.error_i_acumm_2_sqmuxa ));
    LocalMux I__9503 (
            .O(N__51678),
            .I(\pid_front.error_i_acumm_2_sqmuxa ));
    LocalMux I__9502 (
            .O(N__51667),
            .I(\pid_front.error_i_acumm_2_sqmuxa ));
    InMux I__9501 (
            .O(N__51660),
            .I(N__51657));
    LocalMux I__9500 (
            .O(N__51657),
            .I(N__51654));
    Odrv4 I__9499 (
            .O(N__51654),
            .I(\pid_front.error_i_acummZ0Z_3 ));
    CEMux I__9498 (
            .O(N__51651),
            .I(N__51648));
    LocalMux I__9497 (
            .O(N__51648),
            .I(N__51644));
    CEMux I__9496 (
            .O(N__51647),
            .I(N__51641));
    Span4Mux_h I__9495 (
            .O(N__51644),
            .I(N__51637));
    LocalMux I__9494 (
            .O(N__51641),
            .I(N__51634));
    CEMux I__9493 (
            .O(N__51640),
            .I(N__51631));
    Span4Mux_h I__9492 (
            .O(N__51637),
            .I(N__51628));
    Span4Mux_h I__9491 (
            .O(N__51634),
            .I(N__51623));
    LocalMux I__9490 (
            .O(N__51631),
            .I(N__51623));
    Odrv4 I__9489 (
            .O(N__51628),
            .I(\pid_front.error_i_acumm_1_sqmuxa_1_i ));
    Odrv4 I__9488 (
            .O(N__51623),
            .I(\pid_front.error_i_acumm_1_sqmuxa_1_i ));
    InMux I__9487 (
            .O(N__51618),
            .I(N__51614));
    InMux I__9486 (
            .O(N__51617),
            .I(N__51606));
    LocalMux I__9485 (
            .O(N__51614),
            .I(N__51603));
    InMux I__9484 (
            .O(N__51613),
            .I(N__51596));
    InMux I__9483 (
            .O(N__51612),
            .I(N__51596));
    InMux I__9482 (
            .O(N__51611),
            .I(N__51596));
    InMux I__9481 (
            .O(N__51610),
            .I(N__51593));
    InMux I__9480 (
            .O(N__51609),
            .I(N__51590));
    LocalMux I__9479 (
            .O(N__51606),
            .I(N__51581));
    Span12Mux_v I__9478 (
            .O(N__51603),
            .I(N__51581));
    LocalMux I__9477 (
            .O(N__51596),
            .I(N__51581));
    LocalMux I__9476 (
            .O(N__51593),
            .I(N__51581));
    LocalMux I__9475 (
            .O(N__51590),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    Odrv12 I__9474 (
            .O(N__51581),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    InMux I__9473 (
            .O(N__51576),
            .I(N__51570));
    InMux I__9472 (
            .O(N__51575),
            .I(N__51570));
    LocalMux I__9471 (
            .O(N__51570),
            .I(N__51567));
    Span4Mux_h I__9470 (
            .O(N__51567),
            .I(N__51564));
    Span4Mux_v I__9469 (
            .O(N__51564),
            .I(N__51561));
    Odrv4 I__9468 (
            .O(N__51561),
            .I(\pid_front.error_d_reg_prevZ0Z_20 ));
    CascadeMux I__9467 (
            .O(N__51558),
            .I(N__51555));
    InMux I__9466 (
            .O(N__51555),
            .I(N__51549));
    InMux I__9465 (
            .O(N__51554),
            .I(N__51549));
    LocalMux I__9464 (
            .O(N__51549),
            .I(N__51546));
    Span4Mux_h I__9463 (
            .O(N__51546),
            .I(N__51543));
    Span4Mux_v I__9462 (
            .O(N__51543),
            .I(N__51540));
    Odrv4 I__9461 (
            .O(N__51540),
            .I(\pid_front.error_d_reg_prevZ0Z_21 ));
    CascadeMux I__9460 (
            .O(N__51537),
            .I(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ));
    InMux I__9459 (
            .O(N__51534),
            .I(N__51531));
    LocalMux I__9458 (
            .O(N__51531),
            .I(N__51527));
    InMux I__9457 (
            .O(N__51530),
            .I(N__51524));
    Span4Mux_v I__9456 (
            .O(N__51527),
            .I(N__51521));
    LocalMux I__9455 (
            .O(N__51524),
            .I(N__51518));
    Sp12to4 I__9454 (
            .O(N__51521),
            .I(N__51515));
    Span12Mux_v I__9453 (
            .O(N__51518),
            .I(N__51510));
    Span12Mux_h I__9452 (
            .O(N__51515),
            .I(N__51510));
    Odrv12 I__9451 (
            .O(N__51510),
            .I(xy_kp_5));
    InMux I__9450 (
            .O(N__51507),
            .I(N__51503));
    InMux I__9449 (
            .O(N__51506),
            .I(N__51500));
    LocalMux I__9448 (
            .O(N__51503),
            .I(N__51497));
    LocalMux I__9447 (
            .O(N__51500),
            .I(N__51494));
    Span4Mux_s3_h I__9446 (
            .O(N__51497),
            .I(N__51491));
    Span4Mux_v I__9445 (
            .O(N__51494),
            .I(N__51488));
    Span4Mux_h I__9444 (
            .O(N__51491),
            .I(N__51485));
    Span4Mux_h I__9443 (
            .O(N__51488),
            .I(N__51482));
    Span4Mux_h I__9442 (
            .O(N__51485),
            .I(N__51479));
    Sp12to4 I__9441 (
            .O(N__51482),
            .I(N__51476));
    Odrv4 I__9440 (
            .O(N__51479),
            .I(xy_kp_6));
    Odrv12 I__9439 (
            .O(N__51476),
            .I(xy_kp_6));
    InMux I__9438 (
            .O(N__51471),
            .I(N__51467));
    InMux I__9437 (
            .O(N__51470),
            .I(N__51464));
    LocalMux I__9436 (
            .O(N__51467),
            .I(N__51461));
    LocalMux I__9435 (
            .O(N__51464),
            .I(N__51458));
    Span4Mux_v I__9434 (
            .O(N__51461),
            .I(N__51455));
    Span12Mux_v I__9433 (
            .O(N__51458),
            .I(N__51452));
    Sp12to4 I__9432 (
            .O(N__51455),
            .I(N__51449));
    Span12Mux_h I__9431 (
            .O(N__51452),
            .I(N__51446));
    Span12Mux_s3_h I__9430 (
            .O(N__51449),
            .I(N__51443));
    Odrv12 I__9429 (
            .O(N__51446),
            .I(xy_kp_7));
    Odrv12 I__9428 (
            .O(N__51443),
            .I(xy_kp_7));
    CEMux I__9427 (
            .O(N__51438),
            .I(N__51435));
    LocalMux I__9426 (
            .O(N__51435),
            .I(N__51432));
    Span4Mux_h I__9425 (
            .O(N__51432),
            .I(N__51429));
    Odrv4 I__9424 (
            .O(N__51429),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    InMux I__9423 (
            .O(N__51426),
            .I(N__51423));
    LocalMux I__9422 (
            .O(N__51423),
            .I(N__51420));
    Odrv12 I__9421 (
            .O(N__51420),
            .I(\dron_frame_decoder_1.N_186 ));
    InMux I__9420 (
            .O(N__51417),
            .I(N__51414));
    LocalMux I__9419 (
            .O(N__51414),
            .I(N__51411));
    Span4Mux_v I__9418 (
            .O(N__51411),
            .I(N__51408));
    Span4Mux_h I__9417 (
            .O(N__51408),
            .I(N__51399));
    InMux I__9416 (
            .O(N__51407),
            .I(N__51386));
    InMux I__9415 (
            .O(N__51406),
            .I(N__51386));
    InMux I__9414 (
            .O(N__51405),
            .I(N__51386));
    InMux I__9413 (
            .O(N__51404),
            .I(N__51386));
    InMux I__9412 (
            .O(N__51403),
            .I(N__51386));
    InMux I__9411 (
            .O(N__51402),
            .I(N__51386));
    Odrv4 I__9410 (
            .O(N__51399),
            .I(\dron_frame_decoder_1.WDT10_0 ));
    LocalMux I__9409 (
            .O(N__51386),
            .I(\dron_frame_decoder_1.WDT10_0 ));
    CascadeMux I__9408 (
            .O(N__51381),
            .I(N__51376));
    CascadeMux I__9407 (
            .O(N__51380),
            .I(N__51373));
    InMux I__9406 (
            .O(N__51379),
            .I(N__51368));
    InMux I__9405 (
            .O(N__51376),
            .I(N__51368));
    InMux I__9404 (
            .O(N__51373),
            .I(N__51365));
    LocalMux I__9403 (
            .O(N__51368),
            .I(N__51362));
    LocalMux I__9402 (
            .O(N__51365),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv12 I__9401 (
            .O(N__51362),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__9400 (
            .O(N__51357),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__9399 (
            .O(N__51354),
            .I(N__51351));
    LocalMux I__9398 (
            .O(N__51351),
            .I(N__51347));
    InMux I__9397 (
            .O(N__51350),
            .I(N__51344));
    Span4Mux_h I__9396 (
            .O(N__51347),
            .I(N__51341));
    LocalMux I__9395 (
            .O(N__51344),
            .I(N__51338));
    Odrv4 I__9394 (
            .O(N__51341),
            .I(front_order_11));
    Odrv12 I__9393 (
            .O(N__51338),
            .I(front_order_11));
    InMux I__9392 (
            .O(N__51333),
            .I(N__51330));
    LocalMux I__9391 (
            .O(N__51330),
            .I(N__51327));
    Odrv4 I__9390 (
            .O(N__51327),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__9389 (
            .O(N__51324),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__9388 (
            .O(N__51321),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__9387 (
            .O(N__51318),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__9386 (
            .O(N__51315),
            .I(\ppm_encoder_1.un1_elevator_cry_13 ));
    InMux I__9385 (
            .O(N__51312),
            .I(N__51308));
    InMux I__9384 (
            .O(N__51311),
            .I(N__51305));
    LocalMux I__9383 (
            .O(N__51308),
            .I(N__51302));
    LocalMux I__9382 (
            .O(N__51305),
            .I(N__51299));
    Span4Mux_s3_h I__9381 (
            .O(N__51302),
            .I(N__51296));
    Span4Mux_v I__9380 (
            .O(N__51299),
            .I(N__51293));
    Span4Mux_h I__9379 (
            .O(N__51296),
            .I(N__51290));
    Sp12to4 I__9378 (
            .O(N__51293),
            .I(N__51287));
    Span4Mux_h I__9377 (
            .O(N__51290),
            .I(N__51284));
    Span12Mux_s9_h I__9376 (
            .O(N__51287),
            .I(N__51281));
    Odrv4 I__9375 (
            .O(N__51284),
            .I(xy_kp_0));
    Odrv12 I__9374 (
            .O(N__51281),
            .I(xy_kp_0));
    InMux I__9373 (
            .O(N__51276),
            .I(N__51273));
    LocalMux I__9372 (
            .O(N__51273),
            .I(N__51269));
    InMux I__9371 (
            .O(N__51272),
            .I(N__51266));
    Span4Mux_v I__9370 (
            .O(N__51269),
            .I(N__51263));
    LocalMux I__9369 (
            .O(N__51266),
            .I(N__51260));
    Span4Mux_h I__9368 (
            .O(N__51263),
            .I(N__51257));
    Span12Mux_v I__9367 (
            .O(N__51260),
            .I(N__51254));
    Span4Mux_h I__9366 (
            .O(N__51257),
            .I(N__51251));
    Span12Mux_h I__9365 (
            .O(N__51254),
            .I(N__51248));
    Span4Mux_h I__9364 (
            .O(N__51251),
            .I(N__51245));
    Odrv12 I__9363 (
            .O(N__51248),
            .I(xy_kp_1));
    Odrv4 I__9362 (
            .O(N__51245),
            .I(xy_kp_1));
    InMux I__9361 (
            .O(N__51240),
            .I(N__51237));
    LocalMux I__9360 (
            .O(N__51237),
            .I(N__51233));
    InMux I__9359 (
            .O(N__51236),
            .I(N__51230));
    Span4Mux_s2_h I__9358 (
            .O(N__51233),
            .I(N__51227));
    LocalMux I__9357 (
            .O(N__51230),
            .I(N__51224));
    Span4Mux_h I__9356 (
            .O(N__51227),
            .I(N__51221));
    Span12Mux_s0_h I__9355 (
            .O(N__51224),
            .I(N__51218));
    Span4Mux_h I__9354 (
            .O(N__51221),
            .I(N__51215));
    Span12Mux_h I__9353 (
            .O(N__51218),
            .I(N__51212));
    Span4Mux_h I__9352 (
            .O(N__51215),
            .I(N__51209));
    Odrv12 I__9351 (
            .O(N__51212),
            .I(xy_kp_2));
    Odrv4 I__9350 (
            .O(N__51209),
            .I(xy_kp_2));
    InMux I__9349 (
            .O(N__51204),
            .I(N__51200));
    InMux I__9348 (
            .O(N__51203),
            .I(N__51197));
    LocalMux I__9347 (
            .O(N__51200),
            .I(N__51194));
    LocalMux I__9346 (
            .O(N__51197),
            .I(N__51191));
    Span4Mux_v I__9345 (
            .O(N__51194),
            .I(N__51188));
    Span12Mux_v I__9344 (
            .O(N__51191),
            .I(N__51185));
    Sp12to4 I__9343 (
            .O(N__51188),
            .I(N__51182));
    Span12Mux_h I__9342 (
            .O(N__51185),
            .I(N__51179));
    Span12Mux_s6_h I__9341 (
            .O(N__51182),
            .I(N__51176));
    Odrv12 I__9340 (
            .O(N__51179),
            .I(xy_kp_3));
    Odrv12 I__9339 (
            .O(N__51176),
            .I(xy_kp_3));
    InMux I__9338 (
            .O(N__51171),
            .I(\ppm_encoder_1.un1_elevator_cry_1 ));
    InMux I__9337 (
            .O(N__51168),
            .I(\ppm_encoder_1.un1_elevator_cry_2 ));
    InMux I__9336 (
            .O(N__51165),
            .I(\ppm_encoder_1.un1_elevator_cry_3 ));
    InMux I__9335 (
            .O(N__51162),
            .I(\ppm_encoder_1.un1_elevator_cry_4 ));
    InMux I__9334 (
            .O(N__51159),
            .I(N__51156));
    LocalMux I__9333 (
            .O(N__51156),
            .I(N__51152));
    InMux I__9332 (
            .O(N__51155),
            .I(N__51149));
    Span4Mux_h I__9331 (
            .O(N__51152),
            .I(N__51146));
    LocalMux I__9330 (
            .O(N__51149),
            .I(N__51143));
    Span4Mux_v I__9329 (
            .O(N__51146),
            .I(N__51138));
    Span4Mux_h I__9328 (
            .O(N__51143),
            .I(N__51138));
    Odrv4 I__9327 (
            .O(N__51138),
            .I(front_order_6));
    InMux I__9326 (
            .O(N__51135),
            .I(N__51132));
    LocalMux I__9325 (
            .O(N__51132),
            .I(N__51129));
    Odrv12 I__9324 (
            .O(N__51129),
            .I(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ));
    InMux I__9323 (
            .O(N__51126),
            .I(\ppm_encoder_1.un1_elevator_cry_5 ));
    InMux I__9322 (
            .O(N__51123),
            .I(N__51119));
    InMux I__9321 (
            .O(N__51122),
            .I(N__51116));
    LocalMux I__9320 (
            .O(N__51119),
            .I(N__51113));
    LocalMux I__9319 (
            .O(N__51116),
            .I(N__51110));
    Span4Mux_h I__9318 (
            .O(N__51113),
            .I(N__51107));
    Span4Mux_h I__9317 (
            .O(N__51110),
            .I(N__51104));
    Odrv4 I__9316 (
            .O(N__51107),
            .I(front_order_7));
    Odrv4 I__9315 (
            .O(N__51104),
            .I(front_order_7));
    CascadeMux I__9314 (
            .O(N__51099),
            .I(N__51096));
    InMux I__9313 (
            .O(N__51096),
            .I(N__51093));
    LocalMux I__9312 (
            .O(N__51093),
            .I(N__51090));
    Odrv12 I__9311 (
            .O(N__51090),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__9310 (
            .O(N__51087),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__9309 (
            .O(N__51084),
            .I(bfn_13_12_0_));
    InMux I__9308 (
            .O(N__51081),
            .I(N__51078));
    LocalMux I__9307 (
            .O(N__51078),
            .I(N__51075));
    Span4Mux_h I__9306 (
            .O(N__51075),
            .I(N__51071));
    InMux I__9305 (
            .O(N__51074),
            .I(N__51068));
    Span4Mux_h I__9304 (
            .O(N__51071),
            .I(N__51065));
    LocalMux I__9303 (
            .O(N__51068),
            .I(N__51062));
    Odrv4 I__9302 (
            .O(N__51065),
            .I(front_order_9));
    Odrv4 I__9301 (
            .O(N__51062),
            .I(front_order_9));
    InMux I__9300 (
            .O(N__51057),
            .I(N__51054));
    LocalMux I__9299 (
            .O(N__51054),
            .I(N__51051));
    Odrv4 I__9298 (
            .O(N__51051),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__9297 (
            .O(N__51048),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__9296 (
            .O(N__51045),
            .I(N__51042));
    LocalMux I__9295 (
            .O(N__51042),
            .I(N__51039));
    Span4Mux_h I__9294 (
            .O(N__51039),
            .I(N__51035));
    InMux I__9293 (
            .O(N__51038),
            .I(N__51032));
    Odrv4 I__9292 (
            .O(N__51035),
            .I(scaler_4_data_11));
    LocalMux I__9291 (
            .O(N__51032),
            .I(scaler_4_data_11));
    InMux I__9290 (
            .O(N__51027),
            .I(N__51024));
    LocalMux I__9289 (
            .O(N__51024),
            .I(N__51021));
    Odrv4 I__9288 (
            .O(N__51021),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__9287 (
            .O(N__51018),
            .I(N__51014));
    InMux I__9286 (
            .O(N__51017),
            .I(N__51010));
    LocalMux I__9285 (
            .O(N__51014),
            .I(N__51007));
    InMux I__9284 (
            .O(N__51013),
            .I(N__51004));
    LocalMux I__9283 (
            .O(N__51010),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv12 I__9282 (
            .O(N__51007),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    LocalMux I__9281 (
            .O(N__51004),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__9280 (
            .O(N__50997),
            .I(N__50994));
    LocalMux I__9279 (
            .O(N__50994),
            .I(N__50991));
    Odrv4 I__9278 (
            .O(N__50991),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    CascadeMux I__9277 (
            .O(N__50988),
            .I(N__50985));
    InMux I__9276 (
            .O(N__50985),
            .I(N__50982));
    LocalMux I__9275 (
            .O(N__50982),
            .I(N__50979));
    Span4Mux_h I__9274 (
            .O(N__50979),
            .I(N__50975));
    InMux I__9273 (
            .O(N__50978),
            .I(N__50972));
    Odrv4 I__9272 (
            .O(N__50975),
            .I(scaler_4_data_12));
    LocalMux I__9271 (
            .O(N__50972),
            .I(scaler_4_data_12));
    InMux I__9270 (
            .O(N__50967),
            .I(N__50964));
    LocalMux I__9269 (
            .O(N__50964),
            .I(N__50961));
    Span4Mux_v I__9268 (
            .O(N__50961),
            .I(N__50957));
    InMux I__9267 (
            .O(N__50960),
            .I(N__50954));
    Odrv4 I__9266 (
            .O(N__50957),
            .I(scaler_4_data_8));
    LocalMux I__9265 (
            .O(N__50954),
            .I(scaler_4_data_8));
    InMux I__9264 (
            .O(N__50949),
            .I(N__50946));
    LocalMux I__9263 (
            .O(N__50946),
            .I(N__50943));
    Span4Mux_v I__9262 (
            .O(N__50943),
            .I(N__50940));
    Odrv4 I__9261 (
            .O(N__50940),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__9260 (
            .O(N__50937),
            .I(N__50934));
    LocalMux I__9259 (
            .O(N__50934),
            .I(N__50931));
    Odrv4 I__9258 (
            .O(N__50931),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__9257 (
            .O(N__50928),
            .I(N__50925));
    LocalMux I__9256 (
            .O(N__50925),
            .I(N__50922));
    Span4Mux_h I__9255 (
            .O(N__50922),
            .I(N__50918));
    InMux I__9254 (
            .O(N__50921),
            .I(N__50915));
    Odrv4 I__9253 (
            .O(N__50918),
            .I(scaler_4_data_9));
    LocalMux I__9252 (
            .O(N__50915),
            .I(scaler_4_data_9));
    InMux I__9251 (
            .O(N__50910),
            .I(N__50907));
    LocalMux I__9250 (
            .O(N__50907),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__9249 (
            .O(N__50904),
            .I(N__50900));
    InMux I__9248 (
            .O(N__50903),
            .I(N__50897));
    LocalMux I__9247 (
            .O(N__50900),
            .I(N__50894));
    LocalMux I__9246 (
            .O(N__50897),
            .I(N__50891));
    Span4Mux_v I__9245 (
            .O(N__50894),
            .I(N__50888));
    Span12Mux_h I__9244 (
            .O(N__50891),
            .I(N__50885));
    Sp12to4 I__9243 (
            .O(N__50888),
            .I(N__50882));
    Odrv12 I__9242 (
            .O(N__50885),
            .I(throttle_order_1));
    Odrv12 I__9241 (
            .O(N__50882),
            .I(throttle_order_1));
    InMux I__9240 (
            .O(N__50877),
            .I(N__50873));
    InMux I__9239 (
            .O(N__50876),
            .I(N__50870));
    LocalMux I__9238 (
            .O(N__50873),
            .I(N__50864));
    LocalMux I__9237 (
            .O(N__50870),
            .I(N__50864));
    CascadeMux I__9236 (
            .O(N__50869),
            .I(N__50861));
    Span4Mux_v I__9235 (
            .O(N__50864),
            .I(N__50858));
    InMux I__9234 (
            .O(N__50861),
            .I(N__50855));
    Span4Mux_h I__9233 (
            .O(N__50858),
            .I(N__50852));
    LocalMux I__9232 (
            .O(N__50855),
            .I(throttle_order_10));
    Odrv4 I__9231 (
            .O(N__50852),
            .I(throttle_order_10));
    InMux I__9230 (
            .O(N__50847),
            .I(N__50844));
    LocalMux I__9229 (
            .O(N__50844),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__9228 (
            .O(N__50841),
            .I(\ppm_encoder_1.un1_elevator_cry_0 ));
    InMux I__9227 (
            .O(N__50838),
            .I(N__50835));
    LocalMux I__9226 (
            .O(N__50835),
            .I(N__50831));
    InMux I__9225 (
            .O(N__50834),
            .I(N__50828));
    Span4Mux_v I__9224 (
            .O(N__50831),
            .I(N__50822));
    LocalMux I__9223 (
            .O(N__50828),
            .I(N__50822));
    CascadeMux I__9222 (
            .O(N__50827),
            .I(N__50819));
    Span4Mux_h I__9221 (
            .O(N__50822),
            .I(N__50816));
    InMux I__9220 (
            .O(N__50819),
            .I(N__50813));
    Span4Mux_h I__9219 (
            .O(N__50816),
            .I(N__50810));
    LocalMux I__9218 (
            .O(N__50813),
            .I(throttle_order_7));
    Odrv4 I__9217 (
            .O(N__50810),
            .I(throttle_order_7));
    InMux I__9216 (
            .O(N__50805),
            .I(N__50802));
    LocalMux I__9215 (
            .O(N__50802),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    CascadeMux I__9214 (
            .O(N__50799),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11_cascade_ ));
    InMux I__9213 (
            .O(N__50796),
            .I(N__50793));
    LocalMux I__9212 (
            .O(N__50793),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11 ));
    CascadeMux I__9211 (
            .O(N__50790),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    InMux I__9210 (
            .O(N__50787),
            .I(N__50784));
    LocalMux I__9209 (
            .O(N__50784),
            .I(N__50781));
    Odrv12 I__9208 (
            .O(N__50781),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    CascadeMux I__9207 (
            .O(N__50778),
            .I(N__50775));
    InMux I__9206 (
            .O(N__50775),
            .I(N__50770));
    InMux I__9205 (
            .O(N__50774),
            .I(N__50765));
    InMux I__9204 (
            .O(N__50773),
            .I(N__50765));
    LocalMux I__9203 (
            .O(N__50770),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    LocalMux I__9202 (
            .O(N__50765),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    CascadeMux I__9201 (
            .O(N__50760),
            .I(N__50755));
    InMux I__9200 (
            .O(N__50759),
            .I(N__50748));
    InMux I__9199 (
            .O(N__50758),
            .I(N__50748));
    InMux I__9198 (
            .O(N__50755),
            .I(N__50748));
    LocalMux I__9197 (
            .O(N__50748),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__9196 (
            .O(N__50745),
            .I(N__50742));
    LocalMux I__9195 (
            .O(N__50742),
            .I(N__50738));
    InMux I__9194 (
            .O(N__50741),
            .I(N__50735));
    Span4Mux_v I__9193 (
            .O(N__50738),
            .I(N__50731));
    LocalMux I__9192 (
            .O(N__50735),
            .I(N__50728));
    InMux I__9191 (
            .O(N__50734),
            .I(N__50725));
    Span4Mux_h I__9190 (
            .O(N__50731),
            .I(N__50720));
    Span4Mux_h I__9189 (
            .O(N__50728),
            .I(N__50720));
    LocalMux I__9188 (
            .O(N__50725),
            .I(throttle_order_11));
    Odrv4 I__9187 (
            .O(N__50720),
            .I(throttle_order_11));
    InMux I__9186 (
            .O(N__50715),
            .I(N__50712));
    LocalMux I__9185 (
            .O(N__50712),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    CascadeMux I__9184 (
            .O(N__50709),
            .I(N__50705));
    CascadeMux I__9183 (
            .O(N__50708),
            .I(N__50701));
    InMux I__9182 (
            .O(N__50705),
            .I(N__50698));
    InMux I__9181 (
            .O(N__50704),
            .I(N__50693));
    InMux I__9180 (
            .O(N__50701),
            .I(N__50693));
    LocalMux I__9179 (
            .O(N__50698),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__9178 (
            .O(N__50693),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    InMux I__9177 (
            .O(N__50688),
            .I(N__50679));
    InMux I__9176 (
            .O(N__50687),
            .I(N__50679));
    InMux I__9175 (
            .O(N__50686),
            .I(N__50679));
    LocalMux I__9174 (
            .O(N__50679),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    CascadeMux I__9173 (
            .O(N__50676),
            .I(N__50671));
    InMux I__9172 (
            .O(N__50675),
            .I(N__50664));
    InMux I__9171 (
            .O(N__50674),
            .I(N__50664));
    InMux I__9170 (
            .O(N__50671),
            .I(N__50664));
    LocalMux I__9169 (
            .O(N__50664),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__9168 (
            .O(N__50661),
            .I(N__50658));
    LocalMux I__9167 (
            .O(N__50658),
            .I(N__50655));
    Odrv4 I__9166 (
            .O(N__50655),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    CascadeMux I__9165 (
            .O(N__50652),
            .I(N__50649));
    InMux I__9164 (
            .O(N__50649),
            .I(N__50645));
    CascadeMux I__9163 (
            .O(N__50648),
            .I(N__50642));
    LocalMux I__9162 (
            .O(N__50645),
            .I(N__50639));
    InMux I__9161 (
            .O(N__50642),
            .I(N__50636));
    Span4Mux_v I__9160 (
            .O(N__50639),
            .I(N__50632));
    LocalMux I__9159 (
            .O(N__50636),
            .I(N__50629));
    CascadeMux I__9158 (
            .O(N__50635),
            .I(N__50626));
    Span4Mux_h I__9157 (
            .O(N__50632),
            .I(N__50621));
    Span4Mux_h I__9156 (
            .O(N__50629),
            .I(N__50621));
    InMux I__9155 (
            .O(N__50626),
            .I(N__50618));
    Span4Mux_h I__9154 (
            .O(N__50621),
            .I(N__50615));
    LocalMux I__9153 (
            .O(N__50618),
            .I(throttle_order_6));
    Odrv4 I__9152 (
            .O(N__50615),
            .I(throttle_order_6));
    CascadeMux I__9151 (
            .O(N__50610),
            .I(N__50605));
    InMux I__9150 (
            .O(N__50609),
            .I(N__50598));
    InMux I__9149 (
            .O(N__50608),
            .I(N__50598));
    InMux I__9148 (
            .O(N__50605),
            .I(N__50598));
    LocalMux I__9147 (
            .O(N__50598),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    CascadeMux I__9146 (
            .O(N__50595),
            .I(N__50590));
    InMux I__9145 (
            .O(N__50594),
            .I(N__50587));
    InMux I__9144 (
            .O(N__50593),
            .I(N__50584));
    InMux I__9143 (
            .O(N__50590),
            .I(N__50581));
    LocalMux I__9142 (
            .O(N__50587),
            .I(N__50578));
    LocalMux I__9141 (
            .O(N__50584),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    LocalMux I__9140 (
            .O(N__50581),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__9139 (
            .O(N__50578),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    CascadeMux I__9138 (
            .O(N__50571),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    InMux I__9137 (
            .O(N__50568),
            .I(N__50565));
    LocalMux I__9136 (
            .O(N__50565),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    InMux I__9135 (
            .O(N__50562),
            .I(N__50553));
    InMux I__9134 (
            .O(N__50561),
            .I(N__50553));
    InMux I__9133 (
            .O(N__50560),
            .I(N__50553));
    LocalMux I__9132 (
            .O(N__50553),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__9131 (
            .O(N__50550),
            .I(N__50547));
    LocalMux I__9130 (
            .O(N__50547),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__9129 (
            .O(N__50544),
            .I(N__50541));
    LocalMux I__9128 (
            .O(N__50541),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__9127 (
            .O(N__50538),
            .I(N__50535));
    LocalMux I__9126 (
            .O(N__50535),
            .I(N__50532));
    Span4Mux_v I__9125 (
            .O(N__50532),
            .I(N__50528));
    InMux I__9124 (
            .O(N__50531),
            .I(N__50525));
    Odrv4 I__9123 (
            .O(N__50528),
            .I(scaler_4_data_7));
    LocalMux I__9122 (
            .O(N__50525),
            .I(scaler_4_data_7));
    CascadeMux I__9121 (
            .O(N__50520),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    InMux I__9120 (
            .O(N__50517),
            .I(N__50514));
    LocalMux I__9119 (
            .O(N__50514),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    CascadeMux I__9118 (
            .O(N__50511),
            .I(\ppm_encoder_1.N_292_cascade_ ));
    CascadeMux I__9117 (
            .O(N__50508),
            .I(\ppm_encoder_1.N_313_cascade_ ));
    InMux I__9116 (
            .O(N__50505),
            .I(N__50502));
    LocalMux I__9115 (
            .O(N__50502),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    CascadeMux I__9114 (
            .O(N__50499),
            .I(N__50496));
    InMux I__9113 (
            .O(N__50496),
            .I(N__50493));
    LocalMux I__9112 (
            .O(N__50493),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__9111 (
            .O(N__50490),
            .I(N__50487));
    LocalMux I__9110 (
            .O(N__50487),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__9109 (
            .O(N__50484),
            .I(N__50481));
    LocalMux I__9108 (
            .O(N__50481),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    InMux I__9107 (
            .O(N__50478),
            .I(N__50475));
    LocalMux I__9106 (
            .O(N__50475),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__9105 (
            .O(N__50472),
            .I(N__50469));
    LocalMux I__9104 (
            .O(N__50469),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__9103 (
            .O(N__50466),
            .I(N__50463));
    LocalMux I__9102 (
            .O(N__50463),
            .I(N__50460));
    Span4Mux_h I__9101 (
            .O(N__50460),
            .I(N__50456));
    InMux I__9100 (
            .O(N__50459),
            .I(N__50453));
    Odrv4 I__9099 (
            .O(N__50456),
            .I(scaler_4_data_10));
    LocalMux I__9098 (
            .O(N__50453),
            .I(scaler_4_data_10));
    InMux I__9097 (
            .O(N__50448),
            .I(N__50445));
    LocalMux I__9096 (
            .O(N__50445),
            .I(N__50441));
    InMux I__9095 (
            .O(N__50444),
            .I(N__50438));
    Span4Mux_h I__9094 (
            .O(N__50441),
            .I(N__50433));
    LocalMux I__9093 (
            .O(N__50438),
            .I(N__50433));
    Odrv4 I__9092 (
            .O(N__50433),
            .I(scaler_4_data_13));
    InMux I__9091 (
            .O(N__50430),
            .I(N__50427));
    LocalMux I__9090 (
            .O(N__50427),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    CascadeMux I__9089 (
            .O(N__50424),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ));
    InMux I__9088 (
            .O(N__50421),
            .I(N__50418));
    LocalMux I__9087 (
            .O(N__50418),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ));
    CascadeMux I__9086 (
            .O(N__50415),
            .I(\ppm_encoder_1.N_232_cascade_ ));
    CascadeMux I__9085 (
            .O(N__50412),
            .I(N__50409));
    InMux I__9084 (
            .O(N__50409),
            .I(N__50406));
    LocalMux I__9083 (
            .O(N__50406),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    CascadeMux I__9082 (
            .O(N__50403),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ));
    InMux I__9081 (
            .O(N__50400),
            .I(N__50394));
    InMux I__9080 (
            .O(N__50399),
            .I(N__50394));
    LocalMux I__9079 (
            .O(N__50394),
            .I(\ppm_encoder_1.N_139_17 ));
    InMux I__9078 (
            .O(N__50391),
            .I(N__50388));
    LocalMux I__9077 (
            .O(N__50388),
            .I(N__50385));
    Odrv4 I__9076 (
            .O(N__50385),
            .I(\ppm_encoder_1.N_139 ));
    InMux I__9075 (
            .O(N__50382),
            .I(N__50376));
    InMux I__9074 (
            .O(N__50381),
            .I(N__50376));
    LocalMux I__9073 (
            .O(N__50376),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    CascadeMux I__9072 (
            .O(N__50373),
            .I(\pid_front.m6_2_03_cascade_ ));
    InMux I__9071 (
            .O(N__50370),
            .I(N__50366));
    InMux I__9070 (
            .O(N__50369),
            .I(N__50363));
    LocalMux I__9069 (
            .O(N__50366),
            .I(N__50360));
    LocalMux I__9068 (
            .O(N__50363),
            .I(N__50357));
    Span12Mux_v I__9067 (
            .O(N__50360),
            .I(N__50350));
    Span4Mux_v I__9066 (
            .O(N__50357),
            .I(N__50347));
    InMux I__9065 (
            .O(N__50356),
            .I(N__50344));
    InMux I__9064 (
            .O(N__50355),
            .I(N__50341));
    InMux I__9063 (
            .O(N__50354),
            .I(N__50338));
    InMux I__9062 (
            .O(N__50353),
            .I(N__50335));
    Span12Mux_h I__9061 (
            .O(N__50350),
            .I(N__50332));
    Sp12to4 I__9060 (
            .O(N__50347),
            .I(N__50329));
    LocalMux I__9059 (
            .O(N__50344),
            .I(N__50326));
    LocalMux I__9058 (
            .O(N__50341),
            .I(N__50319));
    LocalMux I__9057 (
            .O(N__50338),
            .I(N__50319));
    LocalMux I__9056 (
            .O(N__50335),
            .I(N__50319));
    Odrv12 I__9055 (
            .O(N__50332),
            .I(\pid_front.error_5 ));
    Odrv12 I__9054 (
            .O(N__50329),
            .I(\pid_front.error_5 ));
    Odrv4 I__9053 (
            .O(N__50326),
            .I(\pid_front.error_5 ));
    Odrv4 I__9052 (
            .O(N__50319),
            .I(\pid_front.error_5 ));
    InMux I__9051 (
            .O(N__50310),
            .I(N__50307));
    LocalMux I__9050 (
            .O(N__50307),
            .I(N__50303));
    InMux I__9049 (
            .O(N__50306),
            .I(N__50300));
    Span4Mux_s3_h I__9048 (
            .O(N__50303),
            .I(N__50297));
    LocalMux I__9047 (
            .O(N__50300),
            .I(N__50292));
    Sp12to4 I__9046 (
            .O(N__50297),
            .I(N__50289));
    InMux I__9045 (
            .O(N__50296),
            .I(N__50286));
    InMux I__9044 (
            .O(N__50295),
            .I(N__50283));
    Span12Mux_h I__9043 (
            .O(N__50292),
            .I(N__50278));
    Span12Mux_s7_v I__9042 (
            .O(N__50289),
            .I(N__50275));
    LocalMux I__9041 (
            .O(N__50286),
            .I(N__50270));
    LocalMux I__9040 (
            .O(N__50283),
            .I(N__50270));
    InMux I__9039 (
            .O(N__50282),
            .I(N__50265));
    InMux I__9038 (
            .O(N__50281),
            .I(N__50265));
    Odrv12 I__9037 (
            .O(N__50278),
            .I(\pid_front.error_6 ));
    Odrv12 I__9036 (
            .O(N__50275),
            .I(\pid_front.error_6 ));
    Odrv4 I__9035 (
            .O(N__50270),
            .I(\pid_front.error_6 ));
    LocalMux I__9034 (
            .O(N__50265),
            .I(\pid_front.error_6 ));
    CascadeMux I__9033 (
            .O(N__50256),
            .I(\pid_front.N_27_1_cascade_ ));
    CascadeMux I__9032 (
            .O(N__50253),
            .I(\pid_front.N_63_cascade_ ));
    InMux I__9031 (
            .O(N__50250),
            .I(N__50247));
    LocalMux I__9030 (
            .O(N__50247),
            .I(\pid_front.N_41_0 ));
    CascadeMux I__9029 (
            .O(N__50244),
            .I(\pid_front.N_41_0_cascade_ ));
    CascadeMux I__9028 (
            .O(N__50241),
            .I(N__50238));
    InMux I__9027 (
            .O(N__50238),
            .I(N__50235));
    LocalMux I__9026 (
            .O(N__50235),
            .I(N__50232));
    Span4Mux_h I__9025 (
            .O(N__50232),
            .I(N__50229));
    Span4Mux_v I__9024 (
            .O(N__50229),
            .I(N__50226));
    Odrv4 I__9023 (
            .O(N__50226),
            .I(\pid_front.error_i_regZ0Z_10 ));
    InMux I__9022 (
            .O(N__50223),
            .I(N__50219));
    InMux I__9021 (
            .O(N__50222),
            .I(N__50216));
    LocalMux I__9020 (
            .O(N__50219),
            .I(N__50213));
    LocalMux I__9019 (
            .O(N__50216),
            .I(N__50210));
    Span4Mux_v I__9018 (
            .O(N__50213),
            .I(N__50207));
    Span4Mux_v I__9017 (
            .O(N__50210),
            .I(N__50204));
    Span4Mux_v I__9016 (
            .O(N__50207),
            .I(N__50200));
    Span4Mux_h I__9015 (
            .O(N__50204),
            .I(N__50197));
    InMux I__9014 (
            .O(N__50203),
            .I(N__50190));
    Span4Mux_h I__9013 (
            .O(N__50200),
            .I(N__50187));
    Span4Mux_h I__9012 (
            .O(N__50197),
            .I(N__50184));
    InMux I__9011 (
            .O(N__50196),
            .I(N__50181));
    InMux I__9010 (
            .O(N__50195),
            .I(N__50178));
    InMux I__9009 (
            .O(N__50194),
            .I(N__50175));
    InMux I__9008 (
            .O(N__50193),
            .I(N__50172));
    LocalMux I__9007 (
            .O(N__50190),
            .I(N__50165));
    Span4Mux_h I__9006 (
            .O(N__50187),
            .I(N__50165));
    Span4Mux_h I__9005 (
            .O(N__50184),
            .I(N__50165));
    LocalMux I__9004 (
            .O(N__50181),
            .I(N__50158));
    LocalMux I__9003 (
            .O(N__50178),
            .I(N__50158));
    LocalMux I__9002 (
            .O(N__50175),
            .I(N__50158));
    LocalMux I__9001 (
            .O(N__50172),
            .I(\pid_front.error_3 ));
    Odrv4 I__9000 (
            .O(N__50165),
            .I(\pid_front.error_3 ));
    Odrv4 I__8999 (
            .O(N__50158),
            .I(\pid_front.error_3 ));
    InMux I__8998 (
            .O(N__50151),
            .I(N__50147));
    InMux I__8997 (
            .O(N__50150),
            .I(N__50144));
    LocalMux I__8996 (
            .O(N__50147),
            .I(N__50141));
    LocalMux I__8995 (
            .O(N__50144),
            .I(N__50138));
    Span4Mux_s1_h I__8994 (
            .O(N__50141),
            .I(N__50135));
    Span12Mux_v I__8993 (
            .O(N__50138),
            .I(N__50128));
    Sp12to4 I__8992 (
            .O(N__50135),
            .I(N__50125));
    InMux I__8991 (
            .O(N__50134),
            .I(N__50122));
    InMux I__8990 (
            .O(N__50133),
            .I(N__50119));
    InMux I__8989 (
            .O(N__50132),
            .I(N__50116));
    InMux I__8988 (
            .O(N__50131),
            .I(N__50113));
    Span12Mux_h I__8987 (
            .O(N__50128),
            .I(N__50108));
    Span12Mux_s7_v I__8986 (
            .O(N__50125),
            .I(N__50108));
    LocalMux I__8985 (
            .O(N__50122),
            .I(N__50105));
    LocalMux I__8984 (
            .O(N__50119),
            .I(N__50098));
    LocalMux I__8983 (
            .O(N__50116),
            .I(N__50098));
    LocalMux I__8982 (
            .O(N__50113),
            .I(N__50098));
    Odrv12 I__8981 (
            .O(N__50108),
            .I(\pid_front.error_4 ));
    Odrv4 I__8980 (
            .O(N__50105),
            .I(\pid_front.error_4 ));
    Odrv4 I__8979 (
            .O(N__50098),
            .I(\pid_front.error_4 ));
    InMux I__8978 (
            .O(N__50091),
            .I(N__50088));
    LocalMux I__8977 (
            .O(N__50088),
            .I(N__50084));
    InMux I__8976 (
            .O(N__50087),
            .I(N__50081));
    Span4Mux_h I__8975 (
            .O(N__50084),
            .I(N__50078));
    LocalMux I__8974 (
            .O(N__50081),
            .I(\pid_front.N_30_1 ));
    Odrv4 I__8973 (
            .O(N__50078),
            .I(\pid_front.N_30_1 ));
    InMux I__8972 (
            .O(N__50073),
            .I(N__50069));
    InMux I__8971 (
            .O(N__50072),
            .I(N__50065));
    LocalMux I__8970 (
            .O(N__50069),
            .I(N__50062));
    CascadeMux I__8969 (
            .O(N__50068),
            .I(N__50058));
    LocalMux I__8968 (
            .O(N__50065),
            .I(N__50054));
    Span4Mux_v I__8967 (
            .O(N__50062),
            .I(N__50051));
    InMux I__8966 (
            .O(N__50061),
            .I(N__50046));
    InMux I__8965 (
            .O(N__50058),
            .I(N__50046));
    CascadeMux I__8964 (
            .O(N__50057),
            .I(N__50043));
    Span12Mux_h I__8963 (
            .O(N__50054),
            .I(N__50039));
    Span4Mux_h I__8962 (
            .O(N__50051),
            .I(N__50036));
    LocalMux I__8961 (
            .O(N__50046),
            .I(N__50033));
    InMux I__8960 (
            .O(N__50043),
            .I(N__50030));
    InMux I__8959 (
            .O(N__50042),
            .I(N__50027));
    Span12Mux_v I__8958 (
            .O(N__50039),
            .I(N__50024));
    Span4Mux_h I__8957 (
            .O(N__50036),
            .I(N__50019));
    Span4Mux_h I__8956 (
            .O(N__50033),
            .I(N__50019));
    LocalMux I__8955 (
            .O(N__50030),
            .I(N__50016));
    LocalMux I__8954 (
            .O(N__50027),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv12 I__8953 (
            .O(N__50024),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__8952 (
            .O(N__50019),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv12 I__8951 (
            .O(N__50016),
            .I(\pid_alt.stateZ0Z_0 ));
    IoInMux I__8950 (
            .O(N__50007),
            .I(N__50004));
    LocalMux I__8949 (
            .O(N__50004),
            .I(\pid_alt.state_0_0 ));
    InMux I__8948 (
            .O(N__50001),
            .I(\pid_front.error_cry_10 ));
    InMux I__8947 (
            .O(N__49998),
            .I(N__49994));
    InMux I__8946 (
            .O(N__49997),
            .I(N__49991));
    LocalMux I__8945 (
            .O(N__49994),
            .I(N__49988));
    LocalMux I__8944 (
            .O(N__49991),
            .I(N__49985));
    Span4Mux_v I__8943 (
            .O(N__49988),
            .I(N__49981));
    Span4Mux_v I__8942 (
            .O(N__49985),
            .I(N__49978));
    CascadeMux I__8941 (
            .O(N__49984),
            .I(N__49975));
    Span4Mux_v I__8940 (
            .O(N__49981),
            .I(N__49970));
    Span4Mux_h I__8939 (
            .O(N__49978),
            .I(N__49967));
    InMux I__8938 (
            .O(N__49975),
            .I(N__49964));
    InMux I__8937 (
            .O(N__49974),
            .I(N__49961));
    InMux I__8936 (
            .O(N__49973),
            .I(N__49956));
    Span4Mux_h I__8935 (
            .O(N__49970),
            .I(N__49953));
    Span4Mux_h I__8934 (
            .O(N__49967),
            .I(N__49950));
    LocalMux I__8933 (
            .O(N__49964),
            .I(N__49945));
    LocalMux I__8932 (
            .O(N__49961),
            .I(N__49945));
    InMux I__8931 (
            .O(N__49960),
            .I(N__49942));
    InMux I__8930 (
            .O(N__49959),
            .I(N__49939));
    LocalMux I__8929 (
            .O(N__49956),
            .I(N__49932));
    Span4Mux_h I__8928 (
            .O(N__49953),
            .I(N__49932));
    Span4Mux_h I__8927 (
            .O(N__49950),
            .I(N__49932));
    Span4Mux_v I__8926 (
            .O(N__49945),
            .I(N__49927));
    LocalMux I__8925 (
            .O(N__49942),
            .I(N__49927));
    LocalMux I__8924 (
            .O(N__49939),
            .I(\pid_front.error_2 ));
    Odrv4 I__8923 (
            .O(N__49932),
            .I(\pid_front.error_2 ));
    Odrv4 I__8922 (
            .O(N__49927),
            .I(\pid_front.error_2 ));
    CascadeMux I__8921 (
            .O(N__49920),
            .I(\pid_front.g0_11_1_cascade_ ));
    CascadeMux I__8920 (
            .O(N__49917),
            .I(\pid_front.N_12_1_0_cascade_ ));
    CascadeMux I__8919 (
            .O(N__49914),
            .I(\pid_front.N_116_0_0_cascade_ ));
    InMux I__8918 (
            .O(N__49911),
            .I(N__49908));
    LocalMux I__8917 (
            .O(N__49908),
            .I(N__49905));
    Span4Mux_h I__8916 (
            .O(N__49905),
            .I(N__49902));
    Odrv4 I__8915 (
            .O(N__49902),
            .I(\pid_front.N_117_0 ));
    InMux I__8914 (
            .O(N__49899),
            .I(N__49896));
    LocalMux I__8913 (
            .O(N__49896),
            .I(N__49893));
    Span4Mux_h I__8912 (
            .O(N__49893),
            .I(N__49890));
    Odrv4 I__8911 (
            .O(N__49890),
            .I(\pid_front.un4_error_i_reg_31_ns_1_0 ));
    InMux I__8910 (
            .O(N__49887),
            .I(N__49884));
    LocalMux I__8909 (
            .O(N__49884),
            .I(\pid_front.g0_3_1 ));
    InMux I__8908 (
            .O(N__49881),
            .I(N__49878));
    LocalMux I__8907 (
            .O(N__49878),
            .I(\pid_front.N_89_0_0 ));
    CascadeMux I__8906 (
            .O(N__49875),
            .I(N__49872));
    InMux I__8905 (
            .O(N__49872),
            .I(N__49869));
    LocalMux I__8904 (
            .O(N__49869),
            .I(N__49866));
    Span4Mux_h I__8903 (
            .O(N__49866),
            .I(N__49863));
    Span4Mux_h I__8902 (
            .O(N__49863),
            .I(N__49860));
    Odrv4 I__8901 (
            .O(N__49860),
            .I(front_command_3));
    InMux I__8900 (
            .O(N__49857),
            .I(\pid_front.error_cry_2_0 ));
    InMux I__8899 (
            .O(N__49854),
            .I(N__49851));
    LocalMux I__8898 (
            .O(N__49851),
            .I(N__49848));
    Odrv4 I__8897 (
            .O(N__49848),
            .I(drone_H_disp_front_i_8));
    CascadeMux I__8896 (
            .O(N__49845),
            .I(N__49842));
    InMux I__8895 (
            .O(N__49842),
            .I(N__49839));
    LocalMux I__8894 (
            .O(N__49839),
            .I(N__49836));
    Span4Mux_h I__8893 (
            .O(N__49836),
            .I(N__49833));
    Odrv4 I__8892 (
            .O(N__49833),
            .I(front_command_4));
    InMux I__8891 (
            .O(N__49830),
            .I(bfn_12_24_0_));
    InMux I__8890 (
            .O(N__49827),
            .I(N__49824));
    LocalMux I__8889 (
            .O(N__49824),
            .I(N__49821));
    Span4Mux_v I__8888 (
            .O(N__49821),
            .I(N__49818));
    Span4Mux_h I__8887 (
            .O(N__49818),
            .I(N__49815));
    Span4Mux_v I__8886 (
            .O(N__49815),
            .I(N__49812));
    Odrv4 I__8885 (
            .O(N__49812),
            .I(drone_H_disp_front_i_9));
    CascadeMux I__8884 (
            .O(N__49809),
            .I(N__49806));
    InMux I__8883 (
            .O(N__49806),
            .I(N__49803));
    LocalMux I__8882 (
            .O(N__49803),
            .I(N__49800));
    Span4Mux_h I__8881 (
            .O(N__49800),
            .I(N__49797));
    Span4Mux_v I__8880 (
            .O(N__49797),
            .I(N__49794));
    Odrv4 I__8879 (
            .O(N__49794),
            .I(front_command_5));
    InMux I__8878 (
            .O(N__49791),
            .I(\pid_front.error_cry_4 ));
    CascadeMux I__8877 (
            .O(N__49788),
            .I(N__49785));
    InMux I__8876 (
            .O(N__49785),
            .I(N__49782));
    LocalMux I__8875 (
            .O(N__49782),
            .I(N__49779));
    Span4Mux_h I__8874 (
            .O(N__49779),
            .I(N__49776));
    Span4Mux_v I__8873 (
            .O(N__49776),
            .I(N__49773));
    Odrv4 I__8872 (
            .O(N__49773),
            .I(front_command_6));
    InMux I__8871 (
            .O(N__49770),
            .I(\pid_front.error_cry_5 ));
    InMux I__8870 (
            .O(N__49767),
            .I(N__49764));
    LocalMux I__8869 (
            .O(N__49764),
            .I(N__49761));
    Span12Mux_s10_v I__8868 (
            .O(N__49761),
            .I(N__49758));
    Odrv12 I__8867 (
            .O(N__49758),
            .I(\pid_front.error_axbZ0Z_7 ));
    InMux I__8866 (
            .O(N__49755),
            .I(\pid_front.error_cry_6 ));
    InMux I__8865 (
            .O(N__49752),
            .I(N__49749));
    LocalMux I__8864 (
            .O(N__49749),
            .I(N__49746));
    Sp12to4 I__8863 (
            .O(N__49746),
            .I(N__49743));
    Span12Mux_v I__8862 (
            .O(N__49743),
            .I(N__49740));
    Odrv12 I__8861 (
            .O(N__49740),
            .I(\pid_front.error_axb_8_l_ofx_0 ));
    CascadeMux I__8860 (
            .O(N__49737),
            .I(N__49734));
    InMux I__8859 (
            .O(N__49734),
            .I(N__49731));
    LocalMux I__8858 (
            .O(N__49731),
            .I(N__49728));
    Span4Mux_h I__8857 (
            .O(N__49728),
            .I(N__49724));
    InMux I__8856 (
            .O(N__49727),
            .I(N__49720));
    Span4Mux_h I__8855 (
            .O(N__49724),
            .I(N__49717));
    InMux I__8854 (
            .O(N__49723),
            .I(N__49714));
    LocalMux I__8853 (
            .O(N__49720),
            .I(N__49711));
    Sp12to4 I__8852 (
            .O(N__49717),
            .I(N__49706));
    LocalMux I__8851 (
            .O(N__49714),
            .I(N__49706));
    Odrv12 I__8850 (
            .O(N__49711),
            .I(drone_H_disp_front_12));
    Odrv12 I__8849 (
            .O(N__49706),
            .I(drone_H_disp_front_12));
    InMux I__8848 (
            .O(N__49701),
            .I(\pid_front.error_cry_7 ));
    InMux I__8847 (
            .O(N__49698),
            .I(N__49695));
    LocalMux I__8846 (
            .O(N__49695),
            .I(N__49692));
    Odrv12 I__8845 (
            .O(N__49692),
            .I(drone_H_disp_front_i_12));
    InMux I__8844 (
            .O(N__49689),
            .I(\pid_front.error_cry_8 ));
    InMux I__8843 (
            .O(N__49686),
            .I(\pid_front.error_cry_9 ));
    InMux I__8842 (
            .O(N__49683),
            .I(N__49677));
    InMux I__8841 (
            .O(N__49682),
            .I(N__49677));
    LocalMux I__8840 (
            .O(N__49677),
            .I(drone_H_disp_front_2));
    InMux I__8839 (
            .O(N__49674),
            .I(N__49670));
    InMux I__8838 (
            .O(N__49673),
            .I(N__49667));
    LocalMux I__8837 (
            .O(N__49670),
            .I(dron_frame_decoder_1_source_H_disp_front_fast_0));
    LocalMux I__8836 (
            .O(N__49667),
            .I(dron_frame_decoder_1_source_H_disp_front_fast_0));
    InMux I__8835 (
            .O(N__49662),
            .I(N__49659));
    LocalMux I__8834 (
            .O(N__49659),
            .I(\pid_front.error_axb_0 ));
    InMux I__8833 (
            .O(N__49656),
            .I(N__49653));
    LocalMux I__8832 (
            .O(N__49653),
            .I(N__49650));
    Odrv4 I__8831 (
            .O(N__49650),
            .I(\pid_front.error_axbZ0Z_1 ));
    InMux I__8830 (
            .O(N__49647),
            .I(N__49643));
    InMux I__8829 (
            .O(N__49646),
            .I(N__49640));
    LocalMux I__8828 (
            .O(N__49643),
            .I(N__49637));
    LocalMux I__8827 (
            .O(N__49640),
            .I(N__49634));
    Span4Mux_v I__8826 (
            .O(N__49637),
            .I(N__49631));
    Span4Mux_v I__8825 (
            .O(N__49634),
            .I(N__49627));
    Span4Mux_h I__8824 (
            .O(N__49631),
            .I(N__49624));
    InMux I__8823 (
            .O(N__49630),
            .I(N__49621));
    Span4Mux_h I__8822 (
            .O(N__49627),
            .I(N__49617));
    Span4Mux_h I__8821 (
            .O(N__49624),
            .I(N__49613));
    LocalMux I__8820 (
            .O(N__49621),
            .I(N__49610));
    InMux I__8819 (
            .O(N__49620),
            .I(N__49606));
    Sp12to4 I__8818 (
            .O(N__49617),
            .I(N__49603));
    InMux I__8817 (
            .O(N__49616),
            .I(N__49600));
    Span4Mux_h I__8816 (
            .O(N__49613),
            .I(N__49595));
    Span4Mux_h I__8815 (
            .O(N__49610),
            .I(N__49595));
    InMux I__8814 (
            .O(N__49609),
            .I(N__49592));
    LocalMux I__8813 (
            .O(N__49606),
            .I(N__49589));
    Odrv12 I__8812 (
            .O(N__49603),
            .I(\pid_front.error_1 ));
    LocalMux I__8811 (
            .O(N__49600),
            .I(\pid_front.error_1 ));
    Odrv4 I__8810 (
            .O(N__49595),
            .I(\pid_front.error_1 ));
    LocalMux I__8809 (
            .O(N__49592),
            .I(\pid_front.error_1 ));
    Odrv4 I__8808 (
            .O(N__49589),
            .I(\pid_front.error_1 ));
    InMux I__8807 (
            .O(N__49578),
            .I(\pid_front.error_cry_0 ));
    InMux I__8806 (
            .O(N__49575),
            .I(N__49572));
    LocalMux I__8805 (
            .O(N__49572),
            .I(\pid_front.error_axbZ0Z_2 ));
    InMux I__8804 (
            .O(N__49569),
            .I(\pid_front.error_cry_1 ));
    InMux I__8803 (
            .O(N__49566),
            .I(N__49563));
    LocalMux I__8802 (
            .O(N__49563),
            .I(N__49560));
    Odrv12 I__8801 (
            .O(N__49560),
            .I(\pid_front.error_axbZ0Z_3 ));
    InMux I__8800 (
            .O(N__49557),
            .I(\pid_front.error_cry_2 ));
    InMux I__8799 (
            .O(N__49554),
            .I(N__49551));
    LocalMux I__8798 (
            .O(N__49551),
            .I(N__49548));
    Odrv4 I__8797 (
            .O(N__49548),
            .I(drone_H_disp_front_i_4));
    CascadeMux I__8796 (
            .O(N__49545),
            .I(N__49542));
    InMux I__8795 (
            .O(N__49542),
            .I(N__49539));
    LocalMux I__8794 (
            .O(N__49539),
            .I(N__49536));
    Span4Mux_v I__8793 (
            .O(N__49536),
            .I(N__49533));
    Span4Mux_h I__8792 (
            .O(N__49533),
            .I(N__49530));
    Odrv4 I__8791 (
            .O(N__49530),
            .I(front_command_0));
    InMux I__8790 (
            .O(N__49527),
            .I(\pid_front.error_cry_3 ));
    CascadeMux I__8789 (
            .O(N__49524),
            .I(N__49521));
    InMux I__8788 (
            .O(N__49521),
            .I(N__49518));
    LocalMux I__8787 (
            .O(N__49518),
            .I(N__49515));
    Span4Mux_v I__8786 (
            .O(N__49515),
            .I(N__49512));
    Span4Mux_h I__8785 (
            .O(N__49512),
            .I(N__49509));
    Odrv4 I__8784 (
            .O(N__49509),
            .I(front_command_1));
    InMux I__8783 (
            .O(N__49506),
            .I(\pid_front.error_cry_0_0 ));
    CascadeMux I__8782 (
            .O(N__49503),
            .I(N__49500));
    InMux I__8781 (
            .O(N__49500),
            .I(N__49497));
    LocalMux I__8780 (
            .O(N__49497),
            .I(N__49494));
    Span4Mux_h I__8779 (
            .O(N__49494),
            .I(N__49491));
    Span4Mux_h I__8778 (
            .O(N__49491),
            .I(N__49488));
    Odrv4 I__8777 (
            .O(N__49488),
            .I(front_command_2));
    InMux I__8776 (
            .O(N__49485),
            .I(\pid_front.error_cry_1_0 ));
    InMux I__8775 (
            .O(N__49482),
            .I(N__49479));
    LocalMux I__8774 (
            .O(N__49479),
            .I(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ));
    CascadeMux I__8773 (
            .O(N__49476),
            .I(\pid_front.g2_cascade_ ));
    InMux I__8772 (
            .O(N__49473),
            .I(N__49467));
    InMux I__8771 (
            .O(N__49472),
            .I(N__49467));
    LocalMux I__8770 (
            .O(N__49467),
            .I(\dron_frame_decoder_1.drone_H_disp_front_8 ));
    CascadeMux I__8769 (
            .O(N__49464),
            .I(\pid_front.un1_pid_prereg_0_7_cascade_ ));
    InMux I__8768 (
            .O(N__49461),
            .I(N__49457));
    InMux I__8767 (
            .O(N__49460),
            .I(N__49454));
    LocalMux I__8766 (
            .O(N__49457),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    LocalMux I__8765 (
            .O(N__49454),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    CascadeMux I__8764 (
            .O(N__49449),
            .I(N__49446));
    InMux I__8763 (
            .O(N__49446),
            .I(N__49443));
    LocalMux I__8762 (
            .O(N__49443),
            .I(N__49440));
    Span4Mux_v I__8761 (
            .O(N__49440),
            .I(N__49437));
    Odrv4 I__8760 (
            .O(N__49437),
            .I(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ));
    InMux I__8759 (
            .O(N__49434),
            .I(N__49428));
    InMux I__8758 (
            .O(N__49433),
            .I(N__49428));
    LocalMux I__8757 (
            .O(N__49428),
            .I(N__49425));
    Span4Mux_h I__8756 (
            .O(N__49425),
            .I(N__49422));
    Span4Mux_h I__8755 (
            .O(N__49422),
            .I(N__49419));
    Span4Mux_v I__8754 (
            .O(N__49419),
            .I(N__49416));
    Odrv4 I__8753 (
            .O(N__49416),
            .I(\pid_front.error_p_regZ0Z_17 ));
    InMux I__8752 (
            .O(N__49413),
            .I(N__49407));
    InMux I__8751 (
            .O(N__49412),
            .I(N__49407));
    LocalMux I__8750 (
            .O(N__49407),
            .I(N__49404));
    Span4Mux_v I__8749 (
            .O(N__49404),
            .I(N__49401));
    Span4Mux_h I__8748 (
            .O(N__49401),
            .I(N__49398));
    Odrv4 I__8747 (
            .O(N__49398),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ));
    CascadeMux I__8746 (
            .O(N__49395),
            .I(N__49392));
    InMux I__8745 (
            .O(N__49392),
            .I(N__49386));
    InMux I__8744 (
            .O(N__49391),
            .I(N__49386));
    LocalMux I__8743 (
            .O(N__49386),
            .I(\pid_front.error_d_reg_prevZ0Z_17 ));
    InMux I__8742 (
            .O(N__49383),
            .I(N__49380));
    LocalMux I__8741 (
            .O(N__49380),
            .I(N__49376));
    InMux I__8740 (
            .O(N__49379),
            .I(N__49373));
    Span4Mux_h I__8739 (
            .O(N__49376),
            .I(N__49370));
    LocalMux I__8738 (
            .O(N__49373),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    Odrv4 I__8737 (
            .O(N__49370),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    CascadeMux I__8736 (
            .O(N__49365),
            .I(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ));
    InMux I__8735 (
            .O(N__49362),
            .I(N__49359));
    LocalMux I__8734 (
            .O(N__49359),
            .I(N__49354));
    InMux I__8733 (
            .O(N__49358),
            .I(N__49351));
    CascadeMux I__8732 (
            .O(N__49357),
            .I(N__49348));
    Span4Mux_h I__8731 (
            .O(N__49354),
            .I(N__49345));
    LocalMux I__8730 (
            .O(N__49351),
            .I(N__49342));
    InMux I__8729 (
            .O(N__49348),
            .I(N__49339));
    Span4Mux_v I__8728 (
            .O(N__49345),
            .I(N__49336));
    Span4Mux_h I__8727 (
            .O(N__49342),
            .I(N__49333));
    LocalMux I__8726 (
            .O(N__49339),
            .I(N__49330));
    Odrv4 I__8725 (
            .O(N__49336),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    Odrv4 I__8724 (
            .O(N__49333),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    Odrv4 I__8723 (
            .O(N__49330),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    CascadeMux I__8722 (
            .O(N__49323),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ));
    InMux I__8721 (
            .O(N__49320),
            .I(N__49317));
    LocalMux I__8720 (
            .O(N__49317),
            .I(N__49314));
    Span4Mux_v I__8719 (
            .O(N__49314),
            .I(N__49311));
    Odrv4 I__8718 (
            .O(N__49311),
            .I(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ));
    InMux I__8717 (
            .O(N__49308),
            .I(N__49302));
    InMux I__8716 (
            .O(N__49307),
            .I(N__49302));
    LocalMux I__8715 (
            .O(N__49302),
            .I(N__49299));
    Span4Mux_v I__8714 (
            .O(N__49299),
            .I(N__49296));
    Odrv4 I__8713 (
            .O(N__49296),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    InMux I__8712 (
            .O(N__49293),
            .I(N__49290));
    LocalMux I__8711 (
            .O(N__49290),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ));
    CascadeMux I__8710 (
            .O(N__49287),
            .I(N__49284));
    InMux I__8709 (
            .O(N__49284),
            .I(N__49281));
    LocalMux I__8708 (
            .O(N__49281),
            .I(N__49277));
    InMux I__8707 (
            .O(N__49280),
            .I(N__49274));
    Span4Mux_h I__8706 (
            .O(N__49277),
            .I(N__49269));
    LocalMux I__8705 (
            .O(N__49274),
            .I(N__49269));
    Span4Mux_v I__8704 (
            .O(N__49269),
            .I(N__49266));
    Odrv4 I__8703 (
            .O(N__49266),
            .I(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ));
    InMux I__8702 (
            .O(N__49263),
            .I(N__49260));
    LocalMux I__8701 (
            .O(N__49260),
            .I(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ));
    CascadeMux I__8700 (
            .O(N__49257),
            .I(\pid_front.un1_pid_prereg_0_22_cascade_ ));
    InMux I__8699 (
            .O(N__49254),
            .I(N__49251));
    LocalMux I__8698 (
            .O(N__49251),
            .I(\pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ));
    InMux I__8697 (
            .O(N__49248),
            .I(N__49243));
    InMux I__8696 (
            .O(N__49247),
            .I(N__49238));
    InMux I__8695 (
            .O(N__49246),
            .I(N__49238));
    LocalMux I__8694 (
            .O(N__49243),
            .I(\pid_front.un1_pid_prereg_0_21 ));
    LocalMux I__8693 (
            .O(N__49238),
            .I(\pid_front.un1_pid_prereg_0_21 ));
    InMux I__8692 (
            .O(N__49233),
            .I(N__49227));
    InMux I__8691 (
            .O(N__49232),
            .I(N__49227));
    LocalMux I__8690 (
            .O(N__49227),
            .I(\pid_front.un1_pid_prereg_0_20 ));
    CascadeMux I__8689 (
            .O(N__49224),
            .I(N__49221));
    InMux I__8688 (
            .O(N__49221),
            .I(N__49218));
    LocalMux I__8687 (
            .O(N__49218),
            .I(\pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ));
    InMux I__8686 (
            .O(N__49215),
            .I(N__49212));
    LocalMux I__8685 (
            .O(N__49212),
            .I(N__49209));
    Span4Mux_h I__8684 (
            .O(N__49209),
            .I(N__49205));
    InMux I__8683 (
            .O(N__49208),
            .I(N__49202));
    Odrv4 I__8682 (
            .O(N__49205),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    LocalMux I__8681 (
            .O(N__49202),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    InMux I__8680 (
            .O(N__49197),
            .I(N__49194));
    LocalMux I__8679 (
            .O(N__49194),
            .I(N__49189));
    InMux I__8678 (
            .O(N__49193),
            .I(N__49184));
    InMux I__8677 (
            .O(N__49192),
            .I(N__49184));
    Odrv4 I__8676 (
            .O(N__49189),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    LocalMux I__8675 (
            .O(N__49184),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    CascadeMux I__8674 (
            .O(N__49179),
            .I(N__49176));
    InMux I__8673 (
            .O(N__49176),
            .I(N__49173));
    LocalMux I__8672 (
            .O(N__49173),
            .I(\pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ));
    CascadeMux I__8671 (
            .O(N__49170),
            .I(N__49163));
    CascadeMux I__8670 (
            .O(N__49169),
            .I(N__49159));
    CascadeMux I__8669 (
            .O(N__49168),
            .I(N__49156));
    CascadeMux I__8668 (
            .O(N__49167),
            .I(N__49153));
    CascadeMux I__8667 (
            .O(N__49166),
            .I(N__49149));
    InMux I__8666 (
            .O(N__49163),
            .I(N__49137));
    InMux I__8665 (
            .O(N__49162),
            .I(N__49137));
    InMux I__8664 (
            .O(N__49159),
            .I(N__49137));
    InMux I__8663 (
            .O(N__49156),
            .I(N__49126));
    InMux I__8662 (
            .O(N__49153),
            .I(N__49126));
    InMux I__8661 (
            .O(N__49152),
            .I(N__49126));
    InMux I__8660 (
            .O(N__49149),
            .I(N__49126));
    InMux I__8659 (
            .O(N__49148),
            .I(N__49126));
    CascadeMux I__8658 (
            .O(N__49147),
            .I(N__49123));
    CascadeMux I__8657 (
            .O(N__49146),
            .I(N__49119));
    CascadeMux I__8656 (
            .O(N__49145),
            .I(N__49116));
    CascadeMux I__8655 (
            .O(N__49144),
            .I(N__49113));
    LocalMux I__8654 (
            .O(N__49137),
            .I(N__49110));
    LocalMux I__8653 (
            .O(N__49126),
            .I(N__49107));
    InMux I__8652 (
            .O(N__49123),
            .I(N__49104));
    InMux I__8651 (
            .O(N__49122),
            .I(N__49099));
    InMux I__8650 (
            .O(N__49119),
            .I(N__49099));
    InMux I__8649 (
            .O(N__49116),
            .I(N__49096));
    InMux I__8648 (
            .O(N__49113),
            .I(N__49093));
    Span4Mux_v I__8647 (
            .O(N__49110),
            .I(N__49090));
    Span4Mux_h I__8646 (
            .O(N__49107),
            .I(N__49087));
    LocalMux I__8645 (
            .O(N__49104),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    LocalMux I__8644 (
            .O(N__49099),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    LocalMux I__8643 (
            .O(N__49096),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    LocalMux I__8642 (
            .O(N__49093),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__8641 (
            .O(N__49090),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__8640 (
            .O(N__49087),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    InMux I__8639 (
            .O(N__49074),
            .I(N__49071));
    LocalMux I__8638 (
            .O(N__49071),
            .I(N__49068));
    Span4Mux_h I__8637 (
            .O(N__49068),
            .I(N__49065));
    Odrv4 I__8636 (
            .O(N__49065),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ));
    CascadeMux I__8635 (
            .O(N__49062),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ));
    InMux I__8634 (
            .O(N__49059),
            .I(N__49056));
    LocalMux I__8633 (
            .O(N__49056),
            .I(N__49051));
    InMux I__8632 (
            .O(N__49055),
            .I(N__49048));
    InMux I__8631 (
            .O(N__49054),
            .I(N__49045));
    Span4Mux_v I__8630 (
            .O(N__49051),
            .I(N__49040));
    LocalMux I__8629 (
            .O(N__49048),
            .I(N__49040));
    LocalMux I__8628 (
            .O(N__49045),
            .I(N__49037));
    Odrv4 I__8627 (
            .O(N__49040),
            .I(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ));
    Odrv4 I__8626 (
            .O(N__49037),
            .I(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ));
    InMux I__8625 (
            .O(N__49032),
            .I(N__49029));
    LocalMux I__8624 (
            .O(N__49029),
            .I(N__49026));
    Span4Mux_v I__8623 (
            .O(N__49026),
            .I(N__49022));
    InMux I__8622 (
            .O(N__49025),
            .I(N__49019));
    Odrv4 I__8621 (
            .O(N__49022),
            .I(\pid_front.un1_pid_prereg_0_5 ));
    LocalMux I__8620 (
            .O(N__49019),
            .I(\pid_front.un1_pid_prereg_0_5 ));
    InMux I__8619 (
            .O(N__49014),
            .I(N__49011));
    LocalMux I__8618 (
            .O(N__49011),
            .I(N__49008));
    Span4Mux_v I__8617 (
            .O(N__49008),
            .I(N__49004));
    InMux I__8616 (
            .O(N__49007),
            .I(N__49001));
    Odrv4 I__8615 (
            .O(N__49004),
            .I(\pid_front.un1_pid_prereg_0_4 ));
    LocalMux I__8614 (
            .O(N__49001),
            .I(\pid_front.un1_pid_prereg_0_4 ));
    CascadeMux I__8613 (
            .O(N__48996),
            .I(\pid_front.un1_pid_prereg_0_6_cascade_ ));
    CascadeMux I__8612 (
            .O(N__48993),
            .I(N__48990));
    InMux I__8611 (
            .O(N__48990),
            .I(N__48987));
    LocalMux I__8610 (
            .O(N__48987),
            .I(N__48984));
    Odrv4 I__8609 (
            .O(N__48984),
            .I(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ));
    InMux I__8608 (
            .O(N__48981),
            .I(N__48977));
    InMux I__8607 (
            .O(N__48980),
            .I(N__48974));
    LocalMux I__8606 (
            .O(N__48977),
            .I(N__48971));
    LocalMux I__8605 (
            .O(N__48974),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    Odrv4 I__8604 (
            .O(N__48971),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    InMux I__8603 (
            .O(N__48966),
            .I(N__48963));
    LocalMux I__8602 (
            .O(N__48963),
            .I(N__48960));
    Span4Mux_h I__8601 (
            .O(N__48960),
            .I(N__48956));
    InMux I__8600 (
            .O(N__48959),
            .I(N__48952));
    Sp12to4 I__8599 (
            .O(N__48956),
            .I(N__48949));
    InMux I__8598 (
            .O(N__48955),
            .I(N__48946));
    LocalMux I__8597 (
            .O(N__48952),
            .I(N__48943));
    Odrv12 I__8596 (
            .O(N__48949),
            .I(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ));
    LocalMux I__8595 (
            .O(N__48946),
            .I(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ));
    Odrv4 I__8594 (
            .O(N__48943),
            .I(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ));
    InMux I__8593 (
            .O(N__48936),
            .I(N__48932));
    InMux I__8592 (
            .O(N__48935),
            .I(N__48929));
    LocalMux I__8591 (
            .O(N__48932),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    LocalMux I__8590 (
            .O(N__48929),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    InMux I__8589 (
            .O(N__48924),
            .I(N__48921));
    LocalMux I__8588 (
            .O(N__48921),
            .I(N__48918));
    Span4Mux_h I__8587 (
            .O(N__48918),
            .I(N__48913));
    InMux I__8586 (
            .O(N__48917),
            .I(N__48908));
    InMux I__8585 (
            .O(N__48916),
            .I(N__48908));
    Odrv4 I__8584 (
            .O(N__48913),
            .I(\pid_front.error_p_regZ0Z_11 ));
    LocalMux I__8583 (
            .O(N__48908),
            .I(\pid_front.error_p_regZ0Z_11 ));
    InMux I__8582 (
            .O(N__48903),
            .I(N__48900));
    LocalMux I__8581 (
            .O(N__48900),
            .I(N__48897));
    Span4Mux_h I__8580 (
            .O(N__48897),
            .I(N__48892));
    InMux I__8579 (
            .O(N__48896),
            .I(N__48887));
    InMux I__8578 (
            .O(N__48895),
            .I(N__48887));
    Odrv4 I__8577 (
            .O(N__48892),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    LocalMux I__8576 (
            .O(N__48887),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    InMux I__8575 (
            .O(N__48882),
            .I(N__48879));
    LocalMux I__8574 (
            .O(N__48879),
            .I(N__48875));
    CascadeMux I__8573 (
            .O(N__48878),
            .I(N__48872));
    Span4Mux_h I__8572 (
            .O(N__48875),
            .I(N__48868));
    InMux I__8571 (
            .O(N__48872),
            .I(N__48865));
    InMux I__8570 (
            .O(N__48871),
            .I(N__48862));
    Sp12to4 I__8569 (
            .O(N__48868),
            .I(N__48859));
    LocalMux I__8568 (
            .O(N__48865),
            .I(N__48854));
    LocalMux I__8567 (
            .O(N__48862),
            .I(N__48854));
    Span12Mux_v I__8566 (
            .O(N__48859),
            .I(N__48849));
    Sp12to4 I__8565 (
            .O(N__48854),
            .I(N__48849));
    Odrv12 I__8564 (
            .O(N__48849),
            .I(\pid_front.error_p_regZ0Z_13 ));
    CascadeMux I__8563 (
            .O(N__48846),
            .I(N__48843));
    InMux I__8562 (
            .O(N__48843),
            .I(N__48840));
    LocalMux I__8561 (
            .O(N__48840),
            .I(\pid_front.error_p_reg_esr_RNIETB61Z0Z_13 ));
    InMux I__8560 (
            .O(N__48837),
            .I(N__48831));
    InMux I__8559 (
            .O(N__48836),
            .I(N__48831));
    LocalMux I__8558 (
            .O(N__48831),
            .I(N__48827));
    InMux I__8557 (
            .O(N__48830),
            .I(N__48824));
    Span4Mux_h I__8556 (
            .O(N__48827),
            .I(N__48821));
    LocalMux I__8555 (
            .O(N__48824),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__8554 (
            .O(N__48821),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    InMux I__8553 (
            .O(N__48816),
            .I(N__48811));
    InMux I__8552 (
            .O(N__48815),
            .I(N__48808));
    InMux I__8551 (
            .O(N__48814),
            .I(N__48805));
    LocalMux I__8550 (
            .O(N__48811),
            .I(N__48802));
    LocalMux I__8549 (
            .O(N__48808),
            .I(N__48799));
    LocalMux I__8548 (
            .O(N__48805),
            .I(N__48796));
    Span4Mux_h I__8547 (
            .O(N__48802),
            .I(N__48793));
    Odrv4 I__8546 (
            .O(N__48799),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    Odrv4 I__8545 (
            .O(N__48796),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    Odrv4 I__8544 (
            .O(N__48793),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    CascadeMux I__8543 (
            .O(N__48786),
            .I(N__48783));
    InMux I__8542 (
            .O(N__48783),
            .I(N__48780));
    LocalMux I__8541 (
            .O(N__48780),
            .I(N__48777));
    Span4Mux_v I__8540 (
            .O(N__48777),
            .I(N__48773));
    InMux I__8539 (
            .O(N__48776),
            .I(N__48770));
    Odrv4 I__8538 (
            .O(N__48773),
            .I(\pid_front.un1_pid_prereg_0_1 ));
    LocalMux I__8537 (
            .O(N__48770),
            .I(\pid_front.un1_pid_prereg_0_1 ));
    CascadeMux I__8536 (
            .O(N__48765),
            .I(\pid_front.un1_pid_prereg_0_1_cascade_ ));
    InMux I__8535 (
            .O(N__48762),
            .I(N__48759));
    LocalMux I__8534 (
            .O(N__48759),
            .I(N__48756));
    Span4Mux_h I__8533 (
            .O(N__48756),
            .I(N__48752));
    InMux I__8532 (
            .O(N__48755),
            .I(N__48749));
    Odrv4 I__8531 (
            .O(N__48752),
            .I(\pid_front.un1_pid_prereg_0_0 ));
    LocalMux I__8530 (
            .O(N__48749),
            .I(\pid_front.un1_pid_prereg_0_0 ));
    CascadeMux I__8529 (
            .O(N__48744),
            .I(N__48741));
    InMux I__8528 (
            .O(N__48741),
            .I(N__48738));
    LocalMux I__8527 (
            .O(N__48738),
            .I(N__48735));
    Odrv4 I__8526 (
            .O(N__48735),
            .I(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ));
    InMux I__8525 (
            .O(N__48732),
            .I(N__48729));
    LocalMux I__8524 (
            .O(N__48729),
            .I(N__48724));
    CascadeMux I__8523 (
            .O(N__48728),
            .I(N__48721));
    InMux I__8522 (
            .O(N__48727),
            .I(N__48718));
    Span4Mux_h I__8521 (
            .O(N__48724),
            .I(N__48715));
    InMux I__8520 (
            .O(N__48721),
            .I(N__48712));
    LocalMux I__8519 (
            .O(N__48718),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    Odrv4 I__8518 (
            .O(N__48715),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    LocalMux I__8517 (
            .O(N__48712),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    InMux I__8516 (
            .O(N__48705),
            .I(N__48702));
    LocalMux I__8515 (
            .O(N__48702),
            .I(N__48699));
    Span4Mux_v I__8514 (
            .O(N__48699),
            .I(N__48694));
    InMux I__8513 (
            .O(N__48698),
            .I(N__48689));
    InMux I__8512 (
            .O(N__48697),
            .I(N__48689));
    Odrv4 I__8511 (
            .O(N__48694),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    LocalMux I__8510 (
            .O(N__48689),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    CascadeMux I__8509 (
            .O(N__48684),
            .I(\pid_front.un1_pid_prereg_0_20_cascade_ ));
    InMux I__8508 (
            .O(N__48681),
            .I(N__48678));
    LocalMux I__8507 (
            .O(N__48678),
            .I(N__48675));
    Span4Mux_h I__8506 (
            .O(N__48675),
            .I(N__48671));
    InMux I__8505 (
            .O(N__48674),
            .I(N__48668));
    Odrv4 I__8504 (
            .O(N__48671),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    LocalMux I__8503 (
            .O(N__48668),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    InMux I__8502 (
            .O(N__48663),
            .I(N__48660));
    LocalMux I__8501 (
            .O(N__48660),
            .I(\pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ));
    InMux I__8500 (
            .O(N__48657),
            .I(N__48652));
    InMux I__8499 (
            .O(N__48656),
            .I(N__48647));
    InMux I__8498 (
            .O(N__48655),
            .I(N__48647));
    LocalMux I__8497 (
            .O(N__48652),
            .I(N__48644));
    LocalMux I__8496 (
            .O(N__48647),
            .I(N__48641));
    Span4Mux_h I__8495 (
            .O(N__48644),
            .I(N__48636));
    Span4Mux_v I__8494 (
            .O(N__48641),
            .I(N__48636));
    Odrv4 I__8493 (
            .O(N__48636),
            .I(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ));
    InMux I__8492 (
            .O(N__48633),
            .I(N__48623));
    InMux I__8491 (
            .O(N__48632),
            .I(N__48623));
    InMux I__8490 (
            .O(N__48631),
            .I(N__48619));
    InMux I__8489 (
            .O(N__48630),
            .I(N__48612));
    InMux I__8488 (
            .O(N__48629),
            .I(N__48612));
    InMux I__8487 (
            .O(N__48628),
            .I(N__48612));
    LocalMux I__8486 (
            .O(N__48623),
            .I(N__48605));
    CascadeMux I__8485 (
            .O(N__48622),
            .I(N__48600));
    LocalMux I__8484 (
            .O(N__48619),
            .I(N__48595));
    LocalMux I__8483 (
            .O(N__48612),
            .I(N__48592));
    InMux I__8482 (
            .O(N__48611),
            .I(N__48589));
    InMux I__8481 (
            .O(N__48610),
            .I(N__48582));
    InMux I__8480 (
            .O(N__48609),
            .I(N__48582));
    InMux I__8479 (
            .O(N__48608),
            .I(N__48582));
    Span4Mux_h I__8478 (
            .O(N__48605),
            .I(N__48579));
    InMux I__8477 (
            .O(N__48604),
            .I(N__48568));
    InMux I__8476 (
            .O(N__48603),
            .I(N__48568));
    InMux I__8475 (
            .O(N__48600),
            .I(N__48568));
    InMux I__8474 (
            .O(N__48599),
            .I(N__48568));
    InMux I__8473 (
            .O(N__48598),
            .I(N__48568));
    Span4Mux_v I__8472 (
            .O(N__48595),
            .I(N__48565));
    Span4Mux_h I__8471 (
            .O(N__48592),
            .I(N__48560));
    LocalMux I__8470 (
            .O(N__48589),
            .I(N__48560));
    LocalMux I__8469 (
            .O(N__48582),
            .I(N__48553));
    Span4Mux_h I__8468 (
            .O(N__48579),
            .I(N__48553));
    LocalMux I__8467 (
            .O(N__48568),
            .I(N__48553));
    Span4Mux_h I__8466 (
            .O(N__48565),
            .I(N__48548));
    Span4Mux_h I__8465 (
            .O(N__48560),
            .I(N__48548));
    Span4Mux_v I__8464 (
            .O(N__48553),
            .I(N__48545));
    Span4Mux_h I__8463 (
            .O(N__48548),
            .I(N__48542));
    Span4Mux_h I__8462 (
            .O(N__48545),
            .I(N__48539));
    Span4Mux_v I__8461 (
            .O(N__48542),
            .I(N__48536));
    Span4Mux_h I__8460 (
            .O(N__48539),
            .I(N__48533));
    Odrv4 I__8459 (
            .O(N__48536),
            .I(\pid_front.error_p_regZ0Z_21 ));
    Odrv4 I__8458 (
            .O(N__48533),
            .I(\pid_front.error_p_regZ0Z_21 ));
    CascadeMux I__8457 (
            .O(N__48528),
            .I(\pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13_cascade_ ));
    InMux I__8456 (
            .O(N__48525),
            .I(N__48522));
    LocalMux I__8455 (
            .O(N__48522),
            .I(N__48518));
    CascadeMux I__8454 (
            .O(N__48521),
            .I(N__48515));
    Span4Mux_v I__8453 (
            .O(N__48518),
            .I(N__48512));
    InMux I__8452 (
            .O(N__48515),
            .I(N__48509));
    Odrv4 I__8451 (
            .O(N__48512),
            .I(\pid_front.error_d_reg_prev_esr_RNIUBM0GZ0Z_12 ));
    LocalMux I__8450 (
            .O(N__48509),
            .I(\pid_front.error_d_reg_prev_esr_RNIUBM0GZ0Z_12 ));
    InMux I__8449 (
            .O(N__48504),
            .I(N__48501));
    LocalMux I__8448 (
            .O(N__48501),
            .I(\pid_front.error_p_reg_esr_RNI3TJH01Z0Z_13 ));
    InMux I__8447 (
            .O(N__48498),
            .I(N__48495));
    LocalMux I__8446 (
            .O(N__48495),
            .I(\pid_front.error_p_reg_esr_RNI5HTGGZ0Z_13 ));
    InMux I__8445 (
            .O(N__48492),
            .I(N__48486));
    InMux I__8444 (
            .O(N__48491),
            .I(N__48486));
    LocalMux I__8443 (
            .O(N__48486),
            .I(\pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13 ));
    CascadeMux I__8442 (
            .O(N__48483),
            .I(\pid_front.un1_pid_prereg_0_0_cascade_ ));
    CascadeMux I__8441 (
            .O(N__48480),
            .I(N__48477));
    InMux I__8440 (
            .O(N__48477),
            .I(N__48474));
    LocalMux I__8439 (
            .O(N__48474),
            .I(\pid_front.error_p_reg_esr_RNI31A7NZ0Z_13 ));
    InMux I__8438 (
            .O(N__48471),
            .I(N__48465));
    InMux I__8437 (
            .O(N__48470),
            .I(N__48465));
    LocalMux I__8436 (
            .O(N__48465),
            .I(N__48462));
    Span4Mux_h I__8435 (
            .O(N__48462),
            .I(N__48459));
    Odrv4 I__8434 (
            .O(N__48459),
            .I(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ));
    InMux I__8433 (
            .O(N__48456),
            .I(N__48451));
    InMux I__8432 (
            .O(N__48455),
            .I(N__48446));
    InMux I__8431 (
            .O(N__48454),
            .I(N__48446));
    LocalMux I__8430 (
            .O(N__48451),
            .I(N__48443));
    LocalMux I__8429 (
            .O(N__48446),
            .I(N__48440));
    Span4Mux_h I__8428 (
            .O(N__48443),
            .I(N__48437));
    Span4Mux_h I__8427 (
            .O(N__48440),
            .I(N__48434));
    Odrv4 I__8426 (
            .O(N__48437),
            .I(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ));
    Odrv4 I__8425 (
            .O(N__48434),
            .I(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ));
    InMux I__8424 (
            .O(N__48429),
            .I(N__48420));
    InMux I__8423 (
            .O(N__48428),
            .I(N__48420));
    InMux I__8422 (
            .O(N__48427),
            .I(N__48420));
    LocalMux I__8421 (
            .O(N__48420),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    InMux I__8420 (
            .O(N__48417),
            .I(N__48411));
    InMux I__8419 (
            .O(N__48416),
            .I(N__48411));
    LocalMux I__8418 (
            .O(N__48411),
            .I(N__48408));
    Span4Mux_h I__8417 (
            .O(N__48408),
            .I(N__48405));
    Span4Mux_h I__8416 (
            .O(N__48405),
            .I(N__48402));
    Span4Mux_h I__8415 (
            .O(N__48402),
            .I(N__48399));
    Odrv4 I__8414 (
            .O(N__48399),
            .I(\pid_front.error_p_regZ0Z_19 ));
    InMux I__8413 (
            .O(N__48396),
            .I(N__48390));
    InMux I__8412 (
            .O(N__48395),
            .I(N__48390));
    LocalMux I__8411 (
            .O(N__48390),
            .I(\pid_front.error_d_reg_prevZ0Z_19 ));
    InMux I__8410 (
            .O(N__48387),
            .I(N__48384));
    LocalMux I__8409 (
            .O(N__48384),
            .I(N__48381));
    Span4Mux_v I__8408 (
            .O(N__48381),
            .I(N__48377));
    InMux I__8407 (
            .O(N__48380),
            .I(N__48374));
    Odrv4 I__8406 (
            .O(N__48377),
            .I(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ));
    LocalMux I__8405 (
            .O(N__48374),
            .I(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ));
    InMux I__8404 (
            .O(N__48369),
            .I(N__48366));
    LocalMux I__8403 (
            .O(N__48366),
            .I(N__48362));
    InMux I__8402 (
            .O(N__48365),
            .I(N__48359));
    Span4Mux_v I__8401 (
            .O(N__48362),
            .I(N__48356));
    LocalMux I__8400 (
            .O(N__48359),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    Odrv4 I__8399 (
            .O(N__48356),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    InMux I__8398 (
            .O(N__48351),
            .I(N__48341));
    InMux I__8397 (
            .O(N__48350),
            .I(N__48341));
    InMux I__8396 (
            .O(N__48349),
            .I(N__48337));
    InMux I__8395 (
            .O(N__48348),
            .I(N__48334));
    CascadeMux I__8394 (
            .O(N__48347),
            .I(N__48328));
    CascadeMux I__8393 (
            .O(N__48346),
            .I(N__48325));
    LocalMux I__8392 (
            .O(N__48341),
            .I(N__48322));
    InMux I__8391 (
            .O(N__48340),
            .I(N__48317));
    LocalMux I__8390 (
            .O(N__48337),
            .I(N__48313));
    LocalMux I__8389 (
            .O(N__48334),
            .I(N__48310));
    InMux I__8388 (
            .O(N__48333),
            .I(N__48307));
    InMux I__8387 (
            .O(N__48332),
            .I(N__48304));
    InMux I__8386 (
            .O(N__48331),
            .I(N__48301));
    InMux I__8385 (
            .O(N__48328),
            .I(N__48298));
    InMux I__8384 (
            .O(N__48325),
            .I(N__48295));
    Span4Mux_v I__8383 (
            .O(N__48322),
            .I(N__48292));
    InMux I__8382 (
            .O(N__48321),
            .I(N__48287));
    InMux I__8381 (
            .O(N__48320),
            .I(N__48287));
    LocalMux I__8380 (
            .O(N__48317),
            .I(N__48284));
    CascadeMux I__8379 (
            .O(N__48316),
            .I(N__48280));
    Span4Mux_v I__8378 (
            .O(N__48313),
            .I(N__48273));
    Span4Mux_v I__8377 (
            .O(N__48310),
            .I(N__48270));
    LocalMux I__8376 (
            .O(N__48307),
            .I(N__48256));
    LocalMux I__8375 (
            .O(N__48304),
            .I(N__48256));
    LocalMux I__8374 (
            .O(N__48301),
            .I(N__48256));
    LocalMux I__8373 (
            .O(N__48298),
            .I(N__48256));
    LocalMux I__8372 (
            .O(N__48295),
            .I(N__48249));
    Span4Mux_v I__8371 (
            .O(N__48292),
            .I(N__48249));
    LocalMux I__8370 (
            .O(N__48287),
            .I(N__48249));
    Span4Mux_v I__8369 (
            .O(N__48284),
            .I(N__48244));
    InMux I__8368 (
            .O(N__48283),
            .I(N__48241));
    InMux I__8367 (
            .O(N__48280),
            .I(N__48238));
    InMux I__8366 (
            .O(N__48279),
            .I(N__48227));
    InMux I__8365 (
            .O(N__48278),
            .I(N__48227));
    InMux I__8364 (
            .O(N__48277),
            .I(N__48227));
    InMux I__8363 (
            .O(N__48276),
            .I(N__48227));
    Span4Mux_v I__8362 (
            .O(N__48273),
            .I(N__48222));
    Span4Mux_v I__8361 (
            .O(N__48270),
            .I(N__48222));
    InMux I__8360 (
            .O(N__48269),
            .I(N__48211));
    InMux I__8359 (
            .O(N__48268),
            .I(N__48211));
    InMux I__8358 (
            .O(N__48267),
            .I(N__48211));
    InMux I__8357 (
            .O(N__48266),
            .I(N__48211));
    InMux I__8356 (
            .O(N__48265),
            .I(N__48211));
    Span4Mux_v I__8355 (
            .O(N__48256),
            .I(N__48208));
    Span4Mux_h I__8354 (
            .O(N__48249),
            .I(N__48205));
    InMux I__8353 (
            .O(N__48248),
            .I(N__48200));
    InMux I__8352 (
            .O(N__48247),
            .I(N__48200));
    Span4Mux_h I__8351 (
            .O(N__48244),
            .I(N__48197));
    LocalMux I__8350 (
            .O(N__48241),
            .I(N__48192));
    LocalMux I__8349 (
            .O(N__48238),
            .I(N__48192));
    InMux I__8348 (
            .O(N__48237),
            .I(N__48187));
    InMux I__8347 (
            .O(N__48236),
            .I(N__48187));
    LocalMux I__8346 (
            .O(N__48227),
            .I(uart_pc_data_rdy));
    Odrv4 I__8345 (
            .O(N__48222),
            .I(uart_pc_data_rdy));
    LocalMux I__8344 (
            .O(N__48211),
            .I(uart_pc_data_rdy));
    Odrv4 I__8343 (
            .O(N__48208),
            .I(uart_pc_data_rdy));
    Odrv4 I__8342 (
            .O(N__48205),
            .I(uart_pc_data_rdy));
    LocalMux I__8341 (
            .O(N__48200),
            .I(uart_pc_data_rdy));
    Odrv4 I__8340 (
            .O(N__48197),
            .I(uart_pc_data_rdy));
    Odrv12 I__8339 (
            .O(N__48192),
            .I(uart_pc_data_rdy));
    LocalMux I__8338 (
            .O(N__48187),
            .I(uart_pc_data_rdy));
    InMux I__8337 (
            .O(N__48168),
            .I(N__48165));
    LocalMux I__8336 (
            .O(N__48165),
            .I(N__48162));
    Span12Mux_h I__8335 (
            .O(N__48162),
            .I(N__48159));
    Odrv12 I__8334 (
            .O(N__48159),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ));
    CascadeMux I__8333 (
            .O(N__48156),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ));
    InMux I__8332 (
            .O(N__48153),
            .I(N__48149));
    InMux I__8331 (
            .O(N__48152),
            .I(N__48146));
    LocalMux I__8330 (
            .O(N__48149),
            .I(N__48143));
    LocalMux I__8329 (
            .O(N__48146),
            .I(N__48140));
    Span4Mux_h I__8328 (
            .O(N__48143),
            .I(N__48137));
    Span4Mux_h I__8327 (
            .O(N__48140),
            .I(N__48134));
    Span4Mux_v I__8326 (
            .O(N__48137),
            .I(N__48129));
    Span4Mux_v I__8325 (
            .O(N__48134),
            .I(N__48129));
    Odrv4 I__8324 (
            .O(N__48129),
            .I(front_command_7));
    InMux I__8323 (
            .O(N__48126),
            .I(N__48123));
    LocalMux I__8322 (
            .O(N__48123),
            .I(N__48119));
    InMux I__8321 (
            .O(N__48122),
            .I(N__48116));
    Span4Mux_h I__8320 (
            .O(N__48119),
            .I(N__48113));
    LocalMux I__8319 (
            .O(N__48116),
            .I(drone_H_disp_front_11));
    Odrv4 I__8318 (
            .O(N__48113),
            .I(drone_H_disp_front_11));
    InMux I__8317 (
            .O(N__48108),
            .I(N__48104));
    InMux I__8316 (
            .O(N__48107),
            .I(N__48101));
    LocalMux I__8315 (
            .O(N__48104),
            .I(\pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ));
    LocalMux I__8314 (
            .O(N__48101),
            .I(\pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ));
    CascadeMux I__8313 (
            .O(N__48096),
            .I(N__48093));
    InMux I__8312 (
            .O(N__48093),
            .I(N__48090));
    LocalMux I__8311 (
            .O(N__48090),
            .I(\pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ));
    InMux I__8310 (
            .O(N__48087),
            .I(N__48084));
    LocalMux I__8309 (
            .O(N__48084),
            .I(\pid_front.N_1686_i ));
    InMux I__8308 (
            .O(N__48081),
            .I(N__48078));
    LocalMux I__8307 (
            .O(N__48078),
            .I(N__48074));
    InMux I__8306 (
            .O(N__48077),
            .I(N__48070));
    Span4Mux_h I__8305 (
            .O(N__48074),
            .I(N__48067));
    InMux I__8304 (
            .O(N__48073),
            .I(N__48064));
    LocalMux I__8303 (
            .O(N__48070),
            .I(\pid_front.error_p_reg_esr_RNI6J6A4Z0Z_12 ));
    Odrv4 I__8302 (
            .O(N__48067),
            .I(\pid_front.error_p_reg_esr_RNI6J6A4Z0Z_12 ));
    LocalMux I__8301 (
            .O(N__48064),
            .I(\pid_front.error_p_reg_esr_RNI6J6A4Z0Z_12 ));
    InMux I__8300 (
            .O(N__48057),
            .I(N__48049));
    InMux I__8299 (
            .O(N__48056),
            .I(N__48049));
    InMux I__8298 (
            .O(N__48055),
            .I(N__48046));
    InMux I__8297 (
            .O(N__48054),
            .I(N__48043));
    LocalMux I__8296 (
            .O(N__48049),
            .I(N__48040));
    LocalMux I__8295 (
            .O(N__48046),
            .I(N__48037));
    LocalMux I__8294 (
            .O(N__48043),
            .I(N__48034));
    Span4Mux_v I__8293 (
            .O(N__48040),
            .I(N__48029));
    Span4Mux_h I__8292 (
            .O(N__48037),
            .I(N__48029));
    Odrv4 I__8291 (
            .O(N__48034),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    Odrv4 I__8290 (
            .O(N__48029),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    CascadeMux I__8289 (
            .O(N__48024),
            .I(\pid_front.error_d_reg_prev_esr_RNI4CD85Z0Z_12_cascade_ ));
    InMux I__8288 (
            .O(N__48021),
            .I(N__48016));
    CascadeMux I__8287 (
            .O(N__48020),
            .I(N__48012));
    CascadeMux I__8286 (
            .O(N__48019),
            .I(N__48009));
    LocalMux I__8285 (
            .O(N__48016),
            .I(N__48006));
    InMux I__8284 (
            .O(N__48015),
            .I(N__48002));
    InMux I__8283 (
            .O(N__48012),
            .I(N__47997));
    InMux I__8282 (
            .O(N__48009),
            .I(N__47997));
    Span4Mux_h I__8281 (
            .O(N__48006),
            .I(N__47994));
    InMux I__8280 (
            .O(N__48005),
            .I(N__47991));
    LocalMux I__8279 (
            .O(N__48002),
            .I(N__47986));
    LocalMux I__8278 (
            .O(N__47997),
            .I(N__47986));
    Odrv4 I__8277 (
            .O(N__47994),
            .I(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ));
    LocalMux I__8276 (
            .O(N__47991),
            .I(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ));
    Odrv4 I__8275 (
            .O(N__47986),
            .I(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ));
    InMux I__8274 (
            .O(N__47979),
            .I(N__47976));
    LocalMux I__8273 (
            .O(N__47976),
            .I(N__47973));
    Span4Mux_v I__8272 (
            .O(N__47973),
            .I(N__47970));
    Odrv4 I__8271 (
            .O(N__47970),
            .I(\pid_front.un1_pid_prereg_167_0 ));
    InMux I__8270 (
            .O(N__47967),
            .I(N__47964));
    LocalMux I__8269 (
            .O(N__47964),
            .I(N__47961));
    Span4Mux_v I__8268 (
            .O(N__47961),
            .I(N__47957));
    InMux I__8267 (
            .O(N__47960),
            .I(N__47954));
    Odrv4 I__8266 (
            .O(N__47957),
            .I(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ));
    LocalMux I__8265 (
            .O(N__47954),
            .I(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ));
    InMux I__8264 (
            .O(N__47949),
            .I(N__47946));
    LocalMux I__8263 (
            .O(N__47946),
            .I(N__47943));
    Odrv4 I__8262 (
            .O(N__47943),
            .I(\pid_front.un1_pid_prereg_97 ));
    CascadeMux I__8261 (
            .O(N__47940),
            .I(N__47937));
    InMux I__8260 (
            .O(N__47937),
            .I(N__47934));
    LocalMux I__8259 (
            .O(N__47934),
            .I(\pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ));
    CascadeMux I__8258 (
            .O(N__47931),
            .I(N__47928));
    InMux I__8257 (
            .O(N__47928),
            .I(N__47925));
    LocalMux I__8256 (
            .O(N__47925),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ));
    CascadeMux I__8255 (
            .O(N__47922),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ));
    InMux I__8254 (
            .O(N__47919),
            .I(N__47914));
    InMux I__8253 (
            .O(N__47918),
            .I(N__47909));
    InMux I__8252 (
            .O(N__47917),
            .I(N__47909));
    LocalMux I__8251 (
            .O(N__47914),
            .I(N__47906));
    LocalMux I__8250 (
            .O(N__47909),
            .I(N__47903));
    Span12Mux_s10_h I__8249 (
            .O(N__47906),
            .I(N__47900));
    Span4Mux_h I__8248 (
            .O(N__47903),
            .I(N__47897));
    Odrv12 I__8247 (
            .O(N__47900),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ));
    Odrv4 I__8246 (
            .O(N__47897),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ));
    InMux I__8245 (
            .O(N__47892),
            .I(N__47889));
    LocalMux I__8244 (
            .O(N__47889),
            .I(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ));
    CascadeMux I__8243 (
            .O(N__47886),
            .I(N__47882));
    InMux I__8242 (
            .O(N__47885),
            .I(N__47879));
    InMux I__8241 (
            .O(N__47882),
            .I(N__47876));
    LocalMux I__8240 (
            .O(N__47879),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    LocalMux I__8239 (
            .O(N__47876),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    CascadeMux I__8238 (
            .O(N__47871),
            .I(\pid_front.N_1680_i_cascade_ ));
    InMux I__8237 (
            .O(N__47868),
            .I(N__47862));
    InMux I__8236 (
            .O(N__47867),
            .I(N__47862));
    LocalMux I__8235 (
            .O(N__47862),
            .I(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ));
    InMux I__8234 (
            .O(N__47859),
            .I(N__47853));
    InMux I__8233 (
            .O(N__47858),
            .I(N__47853));
    LocalMux I__8232 (
            .O(N__47853),
            .I(N__47850));
    Span4Mux_h I__8231 (
            .O(N__47850),
            .I(N__47847));
    Span4Mux_h I__8230 (
            .O(N__47847),
            .I(N__47844));
    Odrv4 I__8229 (
            .O(N__47844),
            .I(\pid_front.error_p_regZ0Z_9 ));
    CascadeMux I__8228 (
            .O(N__47841),
            .I(N__47838));
    InMux I__8227 (
            .O(N__47838),
            .I(N__47832));
    InMux I__8226 (
            .O(N__47837),
            .I(N__47832));
    LocalMux I__8225 (
            .O(N__47832),
            .I(N__47829));
    Span4Mux_h I__8224 (
            .O(N__47829),
            .I(N__47825));
    InMux I__8223 (
            .O(N__47828),
            .I(N__47822));
    Odrv4 I__8222 (
            .O(N__47825),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    LocalMux I__8221 (
            .O(N__47822),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    InMux I__8220 (
            .O(N__47817),
            .I(N__47814));
    LocalMux I__8219 (
            .O(N__47814),
            .I(\pid_front.N_1680_i ));
    InMux I__8218 (
            .O(N__47811),
            .I(N__47808));
    LocalMux I__8217 (
            .O(N__47808),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ));
    InMux I__8216 (
            .O(N__47805),
            .I(N__47799));
    InMux I__8215 (
            .O(N__47804),
            .I(N__47799));
    LocalMux I__8214 (
            .O(N__47799),
            .I(N__47796));
    Span4Mux_v I__8213 (
            .O(N__47796),
            .I(N__47793));
    Odrv4 I__8212 (
            .O(N__47793),
            .I(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ));
    InMux I__8211 (
            .O(N__47790),
            .I(N__47786));
    CascadeMux I__8210 (
            .O(N__47789),
            .I(N__47783));
    LocalMux I__8209 (
            .O(N__47786),
            .I(N__47780));
    InMux I__8208 (
            .O(N__47783),
            .I(N__47777));
    Span4Mux_v I__8207 (
            .O(N__47780),
            .I(N__47772));
    LocalMux I__8206 (
            .O(N__47777),
            .I(N__47772));
    Odrv4 I__8205 (
            .O(N__47772),
            .I(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ));
    CascadeMux I__8204 (
            .O(N__47769),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ));
    InMux I__8203 (
            .O(N__47766),
            .I(N__47761));
    InMux I__8202 (
            .O(N__47765),
            .I(N__47756));
    InMux I__8201 (
            .O(N__47764),
            .I(N__47756));
    LocalMux I__8200 (
            .O(N__47761),
            .I(N__47753));
    LocalMux I__8199 (
            .O(N__47756),
            .I(N__47750));
    Span4Mux_h I__8198 (
            .O(N__47753),
            .I(N__47747));
    Span4Mux_h I__8197 (
            .O(N__47750),
            .I(N__47744));
    Odrv4 I__8196 (
            .O(N__47747),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ));
    Odrv4 I__8195 (
            .O(N__47744),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ));
    InMux I__8194 (
            .O(N__47739),
            .I(N__47736));
    LocalMux I__8193 (
            .O(N__47736),
            .I(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ));
    CascadeMux I__8192 (
            .O(N__47733),
            .I(N__47727));
    InMux I__8191 (
            .O(N__47732),
            .I(N__47717));
    InMux I__8190 (
            .O(N__47731),
            .I(N__47702));
    InMux I__8189 (
            .O(N__47730),
            .I(N__47702));
    InMux I__8188 (
            .O(N__47727),
            .I(N__47702));
    InMux I__8187 (
            .O(N__47726),
            .I(N__47702));
    InMux I__8186 (
            .O(N__47725),
            .I(N__47702));
    InMux I__8185 (
            .O(N__47724),
            .I(N__47702));
    InMux I__8184 (
            .O(N__47723),
            .I(N__47702));
    InMux I__8183 (
            .O(N__47722),
            .I(N__47689));
    InMux I__8182 (
            .O(N__47721),
            .I(N__47689));
    InMux I__8181 (
            .O(N__47720),
            .I(N__47689));
    LocalMux I__8180 (
            .O(N__47717),
            .I(N__47680));
    LocalMux I__8179 (
            .O(N__47702),
            .I(N__47677));
    InMux I__8178 (
            .O(N__47701),
            .I(N__47664));
    InMux I__8177 (
            .O(N__47700),
            .I(N__47664));
    InMux I__8176 (
            .O(N__47699),
            .I(N__47664));
    InMux I__8175 (
            .O(N__47698),
            .I(N__47664));
    InMux I__8174 (
            .O(N__47697),
            .I(N__47664));
    InMux I__8173 (
            .O(N__47696),
            .I(N__47664));
    LocalMux I__8172 (
            .O(N__47689),
            .I(N__47661));
    InMux I__8171 (
            .O(N__47688),
            .I(N__47656));
    InMux I__8170 (
            .O(N__47687),
            .I(N__47656));
    InMux I__8169 (
            .O(N__47686),
            .I(N__47653));
    InMux I__8168 (
            .O(N__47685),
            .I(N__47650));
    InMux I__8167 (
            .O(N__47684),
            .I(N__47647));
    InMux I__8166 (
            .O(N__47683),
            .I(N__47644));
    Span4Mux_v I__8165 (
            .O(N__47680),
            .I(N__47641));
    Span4Mux_v I__8164 (
            .O(N__47677),
            .I(N__47638));
    LocalMux I__8163 (
            .O(N__47664),
            .I(N__47635));
    Span4Mux_v I__8162 (
            .O(N__47661),
            .I(N__47630));
    LocalMux I__8161 (
            .O(N__47656),
            .I(N__47630));
    LocalMux I__8160 (
            .O(N__47653),
            .I(N__47627));
    LocalMux I__8159 (
            .O(N__47650),
            .I(N__47624));
    LocalMux I__8158 (
            .O(N__47647),
            .I(N__47621));
    LocalMux I__8157 (
            .O(N__47644),
            .I(N__47612));
    Span4Mux_v I__8156 (
            .O(N__47641),
            .I(N__47612));
    Span4Mux_h I__8155 (
            .O(N__47638),
            .I(N__47612));
    Span4Mux_v I__8154 (
            .O(N__47635),
            .I(N__47612));
    Span4Mux_h I__8153 (
            .O(N__47630),
            .I(N__47609));
    Span4Mux_h I__8152 (
            .O(N__47627),
            .I(N__47606));
    Span12Mux_v I__8151 (
            .O(N__47624),
            .I(N__47603));
    Span12Mux_v I__8150 (
            .O(N__47621),
            .I(N__47600));
    Span4Mux_h I__8149 (
            .O(N__47612),
            .I(N__47597));
    Span4Mux_h I__8148 (
            .O(N__47609),
            .I(N__47594));
    Span4Mux_h I__8147 (
            .O(N__47606),
            .I(N__47591));
    Odrv12 I__8146 (
            .O(N__47603),
            .I(\pid_alt.N_76_i ));
    Odrv12 I__8145 (
            .O(N__47600),
            .I(\pid_alt.N_76_i ));
    Odrv4 I__8144 (
            .O(N__47597),
            .I(\pid_alt.N_76_i ));
    Odrv4 I__8143 (
            .O(N__47594),
            .I(\pid_alt.N_76_i ));
    Odrv4 I__8142 (
            .O(N__47591),
            .I(\pid_alt.N_76_i ));
    CascadeMux I__8141 (
            .O(N__47580),
            .I(N__47577));
    InMux I__8140 (
            .O(N__47577),
            .I(N__47574));
    LocalMux I__8139 (
            .O(N__47574),
            .I(N__47571));
    Odrv4 I__8138 (
            .O(N__47571),
            .I(\pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ));
    InMux I__8137 (
            .O(N__47568),
            .I(N__47565));
    LocalMux I__8136 (
            .O(N__47565),
            .I(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ));
    CascadeMux I__8135 (
            .O(N__47562),
            .I(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ));
    InMux I__8134 (
            .O(N__47559),
            .I(N__47554));
    InMux I__8133 (
            .O(N__47558),
            .I(N__47549));
    InMux I__8132 (
            .O(N__47557),
            .I(N__47549));
    LocalMux I__8131 (
            .O(N__47554),
            .I(N__47546));
    LocalMux I__8130 (
            .O(N__47549),
            .I(N__47543));
    Span4Mux_v I__8129 (
            .O(N__47546),
            .I(N__47540));
    Span4Mux_h I__8128 (
            .O(N__47543),
            .I(N__47537));
    Odrv4 I__8127 (
            .O(N__47540),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ));
    Odrv4 I__8126 (
            .O(N__47537),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ));
    InMux I__8125 (
            .O(N__47532),
            .I(N__47529));
    LocalMux I__8124 (
            .O(N__47529),
            .I(N__47526));
    Span4Mux_h I__8123 (
            .O(N__47526),
            .I(N__47522));
    CascadeMux I__8122 (
            .O(N__47525),
            .I(N__47519));
    Span4Mux_v I__8121 (
            .O(N__47522),
            .I(N__47516));
    InMux I__8120 (
            .O(N__47519),
            .I(N__47513));
    Odrv4 I__8119 (
            .O(N__47516),
            .I(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ));
    LocalMux I__8118 (
            .O(N__47513),
            .I(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ));
    InMux I__8117 (
            .O(N__47508),
            .I(N__47502));
    InMux I__8116 (
            .O(N__47507),
            .I(N__47502));
    LocalMux I__8115 (
            .O(N__47502),
            .I(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ));
    InMux I__8114 (
            .O(N__47499),
            .I(N__47493));
    InMux I__8113 (
            .O(N__47498),
            .I(N__47493));
    LocalMux I__8112 (
            .O(N__47493),
            .I(N__47490));
    Span12Mux_v I__8111 (
            .O(N__47490),
            .I(N__47487));
    Odrv12 I__8110 (
            .O(N__47487),
            .I(\pid_front.error_p_regZ0Z_2 ));
    InMux I__8109 (
            .O(N__47484),
            .I(N__47478));
    InMux I__8108 (
            .O(N__47483),
            .I(N__47478));
    LocalMux I__8107 (
            .O(N__47478),
            .I(\pid_front.error_d_reg_prevZ0Z_2 ));
    InMux I__8106 (
            .O(N__47475),
            .I(N__47469));
    InMux I__8105 (
            .O(N__47474),
            .I(N__47469));
    LocalMux I__8104 (
            .O(N__47469),
            .I(N__47466));
    Odrv12 I__8103 (
            .O(N__47466),
            .I(\pid_front.error_p_regZ0Z_3 ));
    InMux I__8102 (
            .O(N__47463),
            .I(N__47457));
    InMux I__8101 (
            .O(N__47462),
            .I(N__47457));
    LocalMux I__8100 (
            .O(N__47457),
            .I(\pid_front.error_d_reg_prevZ0Z_3 ));
    InMux I__8099 (
            .O(N__47454),
            .I(N__47448));
    InMux I__8098 (
            .O(N__47453),
            .I(N__47448));
    LocalMux I__8097 (
            .O(N__47448),
            .I(N__47445));
    Span4Mux_v I__8096 (
            .O(N__47445),
            .I(N__47442));
    Odrv4 I__8095 (
            .O(N__47442),
            .I(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ));
    CascadeMux I__8094 (
            .O(N__47439),
            .I(N__47436));
    InMux I__8093 (
            .O(N__47436),
            .I(N__47433));
    LocalMux I__8092 (
            .O(N__47433),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__8091 (
            .O(N__47430),
            .I(N__47427));
    InMux I__8090 (
            .O(N__47427),
            .I(N__47424));
    LocalMux I__8089 (
            .O(N__47424),
            .I(frame_decoder_OFF4data_6));
    InMux I__8088 (
            .O(N__47421),
            .I(N__47418));
    LocalMux I__8087 (
            .O(N__47418),
            .I(N__47414));
    InMux I__8086 (
            .O(N__47417),
            .I(N__47411));
    Span4Mux_v I__8085 (
            .O(N__47414),
            .I(N__47408));
    LocalMux I__8084 (
            .O(N__47411),
            .I(frame_decoder_OFF4data_7));
    Odrv4 I__8083 (
            .O(N__47408),
            .I(frame_decoder_OFF4data_7));
    CEMux I__8082 (
            .O(N__47403),
            .I(N__47400));
    LocalMux I__8081 (
            .O(N__47400),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__8080 (
            .O(N__47397),
            .I(N__47394));
    LocalMux I__8079 (
            .O(N__47394),
            .I(N__47391));
    Span4Mux_v I__8078 (
            .O(N__47391),
            .I(N__47387));
    InMux I__8077 (
            .O(N__47390),
            .I(N__47384));
    Odrv4 I__8076 (
            .O(N__47387),
            .I(scaler_4_data_4));
    LocalMux I__8075 (
            .O(N__47384),
            .I(scaler_4_data_4));
    InMux I__8074 (
            .O(N__47379),
            .I(N__47376));
    LocalMux I__8073 (
            .O(N__47376),
            .I(N__47373));
    Span4Mux_h I__8072 (
            .O(N__47373),
            .I(N__47370));
    Odrv4 I__8071 (
            .O(N__47370),
            .I(scaler_4_data_5));
    CascadeMux I__8070 (
            .O(N__47367),
            .I(\pid_front.state_ns_0_cascade_ ));
    SRMux I__8069 (
            .O(N__47364),
            .I(N__47359));
    SRMux I__8068 (
            .O(N__47363),
            .I(N__47355));
    InMux I__8067 (
            .O(N__47362),
            .I(N__47352));
    LocalMux I__8066 (
            .O(N__47359),
            .I(N__47349));
    SRMux I__8065 (
            .O(N__47358),
            .I(N__47346));
    LocalMux I__8064 (
            .O(N__47355),
            .I(N__47343));
    LocalMux I__8063 (
            .O(N__47352),
            .I(N__47340));
    Span4Mux_h I__8062 (
            .O(N__47349),
            .I(N__47335));
    LocalMux I__8061 (
            .O(N__47346),
            .I(N__47335));
    Span4Mux_h I__8060 (
            .O(N__47343),
            .I(N__47332));
    Span4Mux_h I__8059 (
            .O(N__47340),
            .I(N__47329));
    Odrv4 I__8058 (
            .O(N__47335),
            .I(\pid_front.un1_reset_0_i ));
    Odrv4 I__8057 (
            .O(N__47332),
            .I(\pid_front.un1_reset_0_i ));
    Odrv4 I__8056 (
            .O(N__47329),
            .I(\pid_front.un1_reset_0_i ));
    CEMux I__8055 (
            .O(N__47322),
            .I(N__47317));
    CEMux I__8054 (
            .O(N__47321),
            .I(N__47314));
    CEMux I__8053 (
            .O(N__47320),
            .I(N__47311));
    LocalMux I__8052 (
            .O(N__47317),
            .I(\pid_front.state_0_1 ));
    LocalMux I__8051 (
            .O(N__47314),
            .I(\pid_front.state_0_1 ));
    LocalMux I__8050 (
            .O(N__47311),
            .I(\pid_front.state_0_1 ));
    InMux I__8049 (
            .O(N__47304),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__8048 (
            .O(N__47301),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__8047 (
            .O(N__47298),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__8046 (
            .O(N__47295),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__8045 (
            .O(N__47292),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    CascadeMux I__8044 (
            .O(N__47289),
            .I(N__47286));
    InMux I__8043 (
            .O(N__47286),
            .I(N__47279));
    InMux I__8042 (
            .O(N__47285),
            .I(N__47279));
    InMux I__8041 (
            .O(N__47284),
            .I(N__47275));
    LocalMux I__8040 (
            .O(N__47279),
            .I(N__47272));
    CascadeMux I__8039 (
            .O(N__47278),
            .I(N__47269));
    LocalMux I__8038 (
            .O(N__47275),
            .I(N__47264));
    Span4Mux_h I__8037 (
            .O(N__47272),
            .I(N__47264));
    InMux I__8036 (
            .O(N__47269),
            .I(N__47261));
    Odrv4 I__8035 (
            .O(N__47264),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__8034 (
            .O(N__47261),
            .I(frame_decoder_OFF4data_0));
    CascadeMux I__8033 (
            .O(N__47256),
            .I(N__47253));
    InMux I__8032 (
            .O(N__47253),
            .I(N__47250));
    LocalMux I__8031 (
            .O(N__47250),
            .I(frame_decoder_OFF4data_1));
    CascadeMux I__8030 (
            .O(N__47247),
            .I(N__47244));
    InMux I__8029 (
            .O(N__47244),
            .I(N__47241));
    LocalMux I__8028 (
            .O(N__47241),
            .I(frame_decoder_OFF4data_2));
    CascadeMux I__8027 (
            .O(N__47238),
            .I(N__47235));
    InMux I__8026 (
            .O(N__47235),
            .I(N__47232));
    LocalMux I__8025 (
            .O(N__47232),
            .I(frame_decoder_OFF4data_3));
    CascadeMux I__8024 (
            .O(N__47229),
            .I(N__47226));
    InMux I__8023 (
            .O(N__47226),
            .I(N__47223));
    LocalMux I__8022 (
            .O(N__47223),
            .I(frame_decoder_OFF4data_4));
    InMux I__8021 (
            .O(N__47220),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__8020 (
            .O(N__47217),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__8019 (
            .O(N__47214),
            .I(N__47211));
    LocalMux I__8018 (
            .O(N__47211),
            .I(N__47207));
    InMux I__8017 (
            .O(N__47210),
            .I(N__47204));
    Span4Mux_v I__8016 (
            .O(N__47207),
            .I(N__47201));
    LocalMux I__8015 (
            .O(N__47204),
            .I(N__47198));
    Span4Mux_v I__8014 (
            .O(N__47201),
            .I(N__47195));
    Span4Mux_h I__8013 (
            .O(N__47198),
            .I(N__47192));
    Span4Mux_h I__8012 (
            .O(N__47195),
            .I(N__47189));
    Span4Mux_h I__8011 (
            .O(N__47192),
            .I(N__47186));
    Odrv4 I__8010 (
            .O(N__47189),
            .I(throttle_order_4));
    Odrv4 I__8009 (
            .O(N__47186),
            .I(throttle_order_4));
    InMux I__8008 (
            .O(N__47181),
            .I(N__47178));
    LocalMux I__8007 (
            .O(N__47178),
            .I(N__47175));
    Odrv4 I__8006 (
            .O(N__47175),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__8005 (
            .O(N__47172),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__8004 (
            .O(N__47169),
            .I(N__47166));
    LocalMux I__8003 (
            .O(N__47166),
            .I(N__47162));
    InMux I__8002 (
            .O(N__47165),
            .I(N__47159));
    Span4Mux_h I__8001 (
            .O(N__47162),
            .I(N__47156));
    LocalMux I__8000 (
            .O(N__47159),
            .I(N__47153));
    Span4Mux_v I__7999 (
            .O(N__47156),
            .I(N__47150));
    Span4Mux_h I__7998 (
            .O(N__47153),
            .I(N__47147));
    Span4Mux_h I__7997 (
            .O(N__47150),
            .I(N__47144));
    Span4Mux_h I__7996 (
            .O(N__47147),
            .I(N__47141));
    Odrv4 I__7995 (
            .O(N__47144),
            .I(throttle_order_5));
    Odrv4 I__7994 (
            .O(N__47141),
            .I(throttle_order_5));
    InMux I__7993 (
            .O(N__47136),
            .I(N__47133));
    LocalMux I__7992 (
            .O(N__47133),
            .I(N__47130));
    Odrv4 I__7991 (
            .O(N__47130),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__7990 (
            .O(N__47127),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__7989 (
            .O(N__47124),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__7988 (
            .O(N__47121),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__7987 (
            .O(N__47118),
            .I(bfn_12_10_0_));
    InMux I__7986 (
            .O(N__47115),
            .I(N__47112));
    LocalMux I__7985 (
            .O(N__47112),
            .I(N__47108));
    CascadeMux I__7984 (
            .O(N__47111),
            .I(N__47104));
    Span4Mux_v I__7983 (
            .O(N__47108),
            .I(N__47101));
    InMux I__7982 (
            .O(N__47107),
            .I(N__47098));
    InMux I__7981 (
            .O(N__47104),
            .I(N__47095));
    Sp12to4 I__7980 (
            .O(N__47101),
            .I(N__47090));
    LocalMux I__7979 (
            .O(N__47098),
            .I(N__47090));
    LocalMux I__7978 (
            .O(N__47095),
            .I(throttle_order_9));
    Odrv12 I__7977 (
            .O(N__47090),
            .I(throttle_order_9));
    InMux I__7976 (
            .O(N__47085),
            .I(N__47082));
    LocalMux I__7975 (
            .O(N__47082),
            .I(N__47079));
    Odrv4 I__7974 (
            .O(N__47079),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__7973 (
            .O(N__47076),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__7972 (
            .O(N__47073),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__7971 (
            .O(N__47070),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__7970 (
            .O(N__47067),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__7969 (
            .O(N__47064),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__7968 (
            .O(N__47061),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__7967 (
            .O(N__47058),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__7966 (
            .O(N__47055),
            .I(N__47052));
    LocalMux I__7965 (
            .O(N__47052),
            .I(scaler_4_data_14));
    InMux I__7964 (
            .O(N__47049),
            .I(bfn_12_8_0_));
    InMux I__7963 (
            .O(N__47046),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    CascadeMux I__7962 (
            .O(N__47043),
            .I(\pid_front.g0_7_1_cascade_ ));
    CascadeMux I__7961 (
            .O(N__47040),
            .I(\pid_front.N_89_0_1_cascade_ ));
    InMux I__7960 (
            .O(N__47037),
            .I(N__47034));
    LocalMux I__7959 (
            .O(N__47034),
            .I(\pid_front.N_12_1_1 ));
    CascadeMux I__7958 (
            .O(N__47031),
            .I(\pid_front.N_116_0_cascade_ ));
    InMux I__7957 (
            .O(N__47028),
            .I(N__47022));
    InMux I__7956 (
            .O(N__47027),
            .I(N__47022));
    LocalMux I__7955 (
            .O(N__47022),
            .I(\pid_front.un4_error_i_reg_23_ns_1 ));
    CascadeMux I__7954 (
            .O(N__47019),
            .I(\pid_front.error_i_reg_9_1_13_cascade_ ));
    InMux I__7953 (
            .O(N__47016),
            .I(N__47013));
    LocalMux I__7952 (
            .O(N__47013),
            .I(\pid_front.N_127 ));
    CascadeMux I__7951 (
            .O(N__47010),
            .I(N__47007));
    InMux I__7950 (
            .O(N__47007),
            .I(N__47004));
    LocalMux I__7949 (
            .O(N__47004),
            .I(N__47001));
    Span4Mux_h I__7948 (
            .O(N__47001),
            .I(N__46998));
    Span4Mux_v I__7947 (
            .O(N__46998),
            .I(N__46995));
    Odrv4 I__7946 (
            .O(N__46995),
            .I(\pid_front.error_i_regZ0Z_13 ));
    IoInMux I__7945 (
            .O(N__46992),
            .I(N__46989));
    LocalMux I__7944 (
            .O(N__46989),
            .I(N__46986));
    Span4Mux_s3_v I__7943 (
            .O(N__46986),
            .I(N__46982));
    InMux I__7942 (
            .O(N__46985),
            .I(N__46979));
    Odrv4 I__7941 (
            .O(N__46982),
            .I(ppm_output_c));
    LocalMux I__7940 (
            .O(N__46979),
            .I(ppm_output_c));
    InMux I__7939 (
            .O(N__46974),
            .I(N__46971));
    LocalMux I__7938 (
            .O(N__46971),
            .I(\ppm_encoder_1.N_134_0 ));
    InMux I__7937 (
            .O(N__46968),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__7936 (
            .O(N__46965),
            .I(N__46962));
    LocalMux I__7935 (
            .O(N__46962),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_17 ));
    InMux I__7934 (
            .O(N__46959),
            .I(N__46956));
    LocalMux I__7933 (
            .O(N__46956),
            .I(\pid_front.N_51_1 ));
    CascadeMux I__7932 (
            .O(N__46953),
            .I(\pid_front.N_51_1_cascade_ ));
    CascadeMux I__7931 (
            .O(N__46950),
            .I(\pid_front.N_47_1_cascade_ ));
    InMux I__7930 (
            .O(N__46947),
            .I(N__46943));
    InMux I__7929 (
            .O(N__46946),
            .I(N__46940));
    LocalMux I__7928 (
            .O(N__46943),
            .I(N__46935));
    LocalMux I__7927 (
            .O(N__46940),
            .I(N__46935));
    Odrv4 I__7926 (
            .O(N__46935),
            .I(\pid_front.N_45_1 ));
    InMux I__7925 (
            .O(N__46932),
            .I(N__46929));
    LocalMux I__7924 (
            .O(N__46929),
            .I(\pid_front.N_126 ));
    CascadeMux I__7923 (
            .O(N__46926),
            .I(\pid_front.N_88_0_cascade_ ));
    InMux I__7922 (
            .O(N__46923),
            .I(N__46917));
    InMux I__7921 (
            .O(N__46922),
            .I(N__46917));
    LocalMux I__7920 (
            .O(N__46917),
            .I(\pid_front.N_89_0 ));
    InMux I__7919 (
            .O(N__46914),
            .I(N__46908));
    InMux I__7918 (
            .O(N__46913),
            .I(N__46908));
    LocalMux I__7917 (
            .O(N__46908),
            .I(\pid_front.N_88_0 ));
    InMux I__7916 (
            .O(N__46905),
            .I(N__46899));
    InMux I__7915 (
            .O(N__46904),
            .I(N__46899));
    LocalMux I__7914 (
            .O(N__46899),
            .I(\pid_front.N_90_0 ));
    InMux I__7913 (
            .O(N__46896),
            .I(N__46893));
    LocalMux I__7912 (
            .O(N__46893),
            .I(\pid_front.g0_6_1 ));
    InMux I__7911 (
            .O(N__46890),
            .I(N__46887));
    LocalMux I__7910 (
            .O(N__46887),
            .I(\pid_front.m5_2_03 ));
    CascadeMux I__7909 (
            .O(N__46884),
            .I(\pid_front.error_i_reg_9_rn_0_17_cascade_ ));
    InMux I__7908 (
            .O(N__46881),
            .I(N__46878));
    LocalMux I__7907 (
            .O(N__46878),
            .I(N__46875));
    Span4Mux_h I__7906 (
            .O(N__46875),
            .I(N__46872));
    Odrv4 I__7905 (
            .O(N__46872),
            .I(\pid_front.error_i_regZ0Z_17 ));
    CascadeMux I__7904 (
            .O(N__46869),
            .I(\pid_front.N_44_1_cascade_ ));
    CascadeMux I__7903 (
            .O(N__46866),
            .I(\pid_front.N_46_1_cascade_ ));
    InMux I__7902 (
            .O(N__46863),
            .I(N__46860));
    LocalMux I__7901 (
            .O(N__46860),
            .I(\pid_front.m27_2_03_0 ));
    InMux I__7900 (
            .O(N__46857),
            .I(N__46854));
    LocalMux I__7899 (
            .O(N__46854),
            .I(\pid_front.N_44_1 ));
    InMux I__7898 (
            .O(N__46851),
            .I(N__46848));
    LocalMux I__7897 (
            .O(N__46848),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_17 ));
    CascadeMux I__7896 (
            .O(N__46845),
            .I(\pid_front.N_50_1_cascade_ ));
    InMux I__7895 (
            .O(N__46842),
            .I(N__46839));
    LocalMux I__7894 (
            .O(N__46839),
            .I(\pid_front.error_i_reg_9_rn_0_19 ));
    InMux I__7893 (
            .O(N__46836),
            .I(N__46833));
    LocalMux I__7892 (
            .O(N__46833),
            .I(N__46830));
    Span4Mux_h I__7891 (
            .O(N__46830),
            .I(N__46827));
    Odrv4 I__7890 (
            .O(N__46827),
            .I(\pid_front.error_i_regZ0Z_19 ));
    InMux I__7889 (
            .O(N__46824),
            .I(N__46818));
    InMux I__7888 (
            .O(N__46823),
            .I(N__46818));
    LocalMux I__7887 (
            .O(N__46818),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ));
    InMux I__7886 (
            .O(N__46815),
            .I(N__46809));
    InMux I__7885 (
            .O(N__46814),
            .I(N__46809));
    LocalMux I__7884 (
            .O(N__46809),
            .I(N__46806));
    Span4Mux_v I__7883 (
            .O(N__46806),
            .I(N__46803));
    Span4Mux_h I__7882 (
            .O(N__46803),
            .I(N__46800));
    Span4Mux_h I__7881 (
            .O(N__46800),
            .I(N__46797));
    Span4Mux_v I__7880 (
            .O(N__46797),
            .I(N__46794));
    Odrv4 I__7879 (
            .O(N__46794),
            .I(\pid_front.error_p_regZ0Z_20 ));
    InMux I__7878 (
            .O(N__46791),
            .I(N__46787));
    InMux I__7877 (
            .O(N__46790),
            .I(N__46784));
    LocalMux I__7876 (
            .O(N__46787),
            .I(N__46781));
    LocalMux I__7875 (
            .O(N__46784),
            .I(\pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ));
    Odrv12 I__7874 (
            .O(N__46781),
            .I(\pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ));
    CascadeMux I__7873 (
            .O(N__46776),
            .I(\pid_front.m14_0_ns_1_cascade_ ));
    CascadeMux I__7872 (
            .O(N__46773),
            .I(\pid_front.N_15_1_cascade_ ));
    CascadeMux I__7871 (
            .O(N__46770),
            .I(\pid_front.m104_1_cascade_ ));
    InMux I__7870 (
            .O(N__46767),
            .I(N__46764));
    LocalMux I__7869 (
            .O(N__46764),
            .I(\pid_front.m11_2_03_3_i_0 ));
    CascadeMux I__7868 (
            .O(N__46761),
            .I(\pid_front.m11_2_03_3_i_0_cascade_ ));
    InMux I__7867 (
            .O(N__46758),
            .I(N__46755));
    LocalMux I__7866 (
            .O(N__46755),
            .I(N__46751));
    InMux I__7865 (
            .O(N__46754),
            .I(N__46748));
    Span4Mux_h I__7864 (
            .O(N__46751),
            .I(N__46745));
    LocalMux I__7863 (
            .O(N__46748),
            .I(\pid_front.error_i_regZ0Z_7 ));
    Odrv4 I__7862 (
            .O(N__46745),
            .I(\pid_front.error_i_regZ0Z_7 ));
    CascadeMux I__7861 (
            .O(N__46740),
            .I(\pid_front.m53_0_ns_1_cascade_ ));
    InMux I__7860 (
            .O(N__46737),
            .I(N__46731));
    InMux I__7859 (
            .O(N__46736),
            .I(N__46731));
    LocalMux I__7858 (
            .O(N__46731),
            .I(\pid_front.un1_pid_prereg_0_11 ));
    CascadeMux I__7857 (
            .O(N__46728),
            .I(\pid_front.un1_pid_prereg_0_11_cascade_ ));
    InMux I__7856 (
            .O(N__46725),
            .I(N__46722));
    LocalMux I__7855 (
            .O(N__46722),
            .I(N__46718));
    InMux I__7854 (
            .O(N__46721),
            .I(N__46715));
    Odrv4 I__7853 (
            .O(N__46718),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    LocalMux I__7852 (
            .O(N__46715),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    CascadeMux I__7851 (
            .O(N__46710),
            .I(N__46707));
    InMux I__7850 (
            .O(N__46707),
            .I(N__46704));
    LocalMux I__7849 (
            .O(N__46704),
            .I(N__46701));
    Span4Mux_h I__7848 (
            .O(N__46701),
            .I(N__46698));
    Odrv4 I__7847 (
            .O(N__46698),
            .I(\pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ));
    InMux I__7846 (
            .O(N__46695),
            .I(N__46689));
    InMux I__7845 (
            .O(N__46694),
            .I(N__46689));
    LocalMux I__7844 (
            .O(N__46689),
            .I(N__46686));
    Span4Mux_h I__7843 (
            .O(N__46686),
            .I(N__46683));
    Span4Mux_h I__7842 (
            .O(N__46683),
            .I(N__46680));
    Odrv4 I__7841 (
            .O(N__46680),
            .I(\pid_front.un1_pid_prereg_370_1 ));
    InMux I__7840 (
            .O(N__46677),
            .I(N__46674));
    LocalMux I__7839 (
            .O(N__46674),
            .I(N__46669));
    InMux I__7838 (
            .O(N__46673),
            .I(N__46664));
    InMux I__7837 (
            .O(N__46672),
            .I(N__46664));
    Odrv4 I__7836 (
            .O(N__46669),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    LocalMux I__7835 (
            .O(N__46664),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    InMux I__7834 (
            .O(N__46659),
            .I(N__46656));
    LocalMux I__7833 (
            .O(N__46656),
            .I(N__46651));
    InMux I__7832 (
            .O(N__46655),
            .I(N__46646));
    InMux I__7831 (
            .O(N__46654),
            .I(N__46646));
    Odrv4 I__7830 (
            .O(N__46651),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    LocalMux I__7829 (
            .O(N__46646),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    InMux I__7828 (
            .O(N__46641),
            .I(N__46637));
    InMux I__7827 (
            .O(N__46640),
            .I(N__46634));
    LocalMux I__7826 (
            .O(N__46637),
            .I(N__46631));
    LocalMux I__7825 (
            .O(N__46634),
            .I(N__46628));
    Span12Mux_h I__7824 (
            .O(N__46631),
            .I(N__46621));
    Span4Mux_h I__7823 (
            .O(N__46628),
            .I(N__46618));
    InMux I__7822 (
            .O(N__46627),
            .I(N__46609));
    InMux I__7821 (
            .O(N__46626),
            .I(N__46609));
    InMux I__7820 (
            .O(N__46625),
            .I(N__46609));
    InMux I__7819 (
            .O(N__46624),
            .I(N__46609));
    Odrv12 I__7818 (
            .O(N__46621),
            .I(\pid_alt.N_62_mux ));
    Odrv4 I__7817 (
            .O(N__46618),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__7816 (
            .O(N__46609),
            .I(\pid_alt.N_62_mux ));
    CascadeMux I__7815 (
            .O(N__46602),
            .I(N__46599));
    InMux I__7814 (
            .O(N__46599),
            .I(N__46596));
    LocalMux I__7813 (
            .O(N__46596),
            .I(N__46592));
    CascadeMux I__7812 (
            .O(N__46595),
            .I(N__46589));
    Span4Mux_h I__7811 (
            .O(N__46592),
            .I(N__46586));
    InMux I__7810 (
            .O(N__46589),
            .I(N__46583));
    Span4Mux_v I__7809 (
            .O(N__46586),
            .I(N__46580));
    LocalMux I__7808 (
            .O(N__46583),
            .I(N__46577));
    Span4Mux_v I__7807 (
            .O(N__46580),
            .I(N__46573));
    Span4Mux_v I__7806 (
            .O(N__46577),
            .I(N__46569));
    InMux I__7805 (
            .O(N__46576),
            .I(N__46566));
    Span4Mux_v I__7804 (
            .O(N__46573),
            .I(N__46563));
    InMux I__7803 (
            .O(N__46572),
            .I(N__46560));
    Span4Mux_h I__7802 (
            .O(N__46569),
            .I(N__46555));
    LocalMux I__7801 (
            .O(N__46566),
            .I(N__46555));
    Span4Mux_h I__7800 (
            .O(N__46563),
            .I(N__46550));
    LocalMux I__7799 (
            .O(N__46560),
            .I(N__46550));
    Odrv4 I__7798 (
            .O(N__46555),
            .I(\pid_alt.error_i_acumm7lto5 ));
    Odrv4 I__7797 (
            .O(N__46550),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__7796 (
            .O(N__46545),
            .I(N__46542));
    LocalMux I__7795 (
            .O(N__46542),
            .I(N__46539));
    Span4Mux_v I__7794 (
            .O(N__46539),
            .I(N__46536));
    Span4Mux_v I__7793 (
            .O(N__46536),
            .I(N__46533));
    Span4Mux_h I__7792 (
            .O(N__46533),
            .I(N__46529));
    InMux I__7791 (
            .O(N__46532),
            .I(N__46526));
    Span4Mux_h I__7790 (
            .O(N__46529),
            .I(N__46523));
    LocalMux I__7789 (
            .O(N__46526),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    Odrv4 I__7788 (
            .O(N__46523),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    SRMux I__7787 (
            .O(N__46518),
            .I(N__46515));
    LocalMux I__7786 (
            .O(N__46515),
            .I(N__46511));
    SRMux I__7785 (
            .O(N__46514),
            .I(N__46508));
    Span4Mux_v I__7784 (
            .O(N__46511),
            .I(N__46504));
    LocalMux I__7783 (
            .O(N__46508),
            .I(N__46500));
    SRMux I__7782 (
            .O(N__46507),
            .I(N__46497));
    Span4Mux_h I__7781 (
            .O(N__46504),
            .I(N__46494));
    SRMux I__7780 (
            .O(N__46503),
            .I(N__46491));
    Span4Mux_v I__7779 (
            .O(N__46500),
            .I(N__46485));
    LocalMux I__7778 (
            .O(N__46497),
            .I(N__46485));
    Span4Mux_v I__7777 (
            .O(N__46494),
            .I(N__46482));
    LocalMux I__7776 (
            .O(N__46491),
            .I(N__46479));
    SRMux I__7775 (
            .O(N__46490),
            .I(N__46476));
    Span4Mux_h I__7774 (
            .O(N__46485),
            .I(N__46473));
    Span4Mux_v I__7773 (
            .O(N__46482),
            .I(N__46466));
    Span4Mux_s3_h I__7772 (
            .O(N__46479),
            .I(N__46466));
    LocalMux I__7771 (
            .O(N__46476),
            .I(N__46466));
    Odrv4 I__7770 (
            .O(N__46473),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__7769 (
            .O(N__46466),
            .I(\pid_alt.un1_reset_1_0_i ));
    InMux I__7768 (
            .O(N__46461),
            .I(N__46458));
    LocalMux I__7767 (
            .O(N__46458),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ));
    CascadeMux I__7766 (
            .O(N__46455),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ));
    InMux I__7765 (
            .O(N__46452),
            .I(N__46449));
    LocalMux I__7764 (
            .O(N__46449),
            .I(N__46444));
    InMux I__7763 (
            .O(N__46448),
            .I(N__46441));
    InMux I__7762 (
            .O(N__46447),
            .I(N__46438));
    Odrv4 I__7761 (
            .O(N__46444),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    LocalMux I__7760 (
            .O(N__46441),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    LocalMux I__7759 (
            .O(N__46438),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    InMux I__7758 (
            .O(N__46431),
            .I(N__46427));
    InMux I__7757 (
            .O(N__46430),
            .I(N__46424));
    LocalMux I__7756 (
            .O(N__46427),
            .I(N__46418));
    LocalMux I__7755 (
            .O(N__46424),
            .I(N__46418));
    InMux I__7754 (
            .O(N__46423),
            .I(N__46415));
    Odrv4 I__7753 (
            .O(N__46418),
            .I(\pid_front.un1_pid_prereg_0_12 ));
    LocalMux I__7752 (
            .O(N__46415),
            .I(\pid_front.un1_pid_prereg_0_12 ));
    InMux I__7751 (
            .O(N__46410),
            .I(N__46406));
    InMux I__7750 (
            .O(N__46409),
            .I(N__46403));
    LocalMux I__7749 (
            .O(N__46406),
            .I(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ));
    LocalMux I__7748 (
            .O(N__46403),
            .I(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ));
    CascadeMux I__7747 (
            .O(N__46398),
            .I(\pid_front.un1_pid_prereg_0_8_cascade_ ));
    InMux I__7746 (
            .O(N__46395),
            .I(N__46392));
    LocalMux I__7745 (
            .O(N__46392),
            .I(N__46389));
    Odrv4 I__7744 (
            .O(N__46389),
            .I(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ));
    CascadeMux I__7743 (
            .O(N__46386),
            .I(N__46383));
    InMux I__7742 (
            .O(N__46383),
            .I(N__46380));
    LocalMux I__7741 (
            .O(N__46380),
            .I(\pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ));
    InMux I__7740 (
            .O(N__46377),
            .I(N__46372));
    InMux I__7739 (
            .O(N__46376),
            .I(N__46369));
    InMux I__7738 (
            .O(N__46375),
            .I(N__46366));
    LocalMux I__7737 (
            .O(N__46372),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    LocalMux I__7736 (
            .O(N__46369),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    LocalMux I__7735 (
            .O(N__46366),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    InMux I__7734 (
            .O(N__46359),
            .I(N__46353));
    InMux I__7733 (
            .O(N__46358),
            .I(N__46353));
    LocalMux I__7732 (
            .O(N__46353),
            .I(\pid_front.un1_pid_prereg_0_13 ));
    CascadeMux I__7731 (
            .O(N__46350),
            .I(\pid_front.un1_pid_prereg_0_13_cascade_ ));
    InMux I__7730 (
            .O(N__46347),
            .I(N__46344));
    LocalMux I__7729 (
            .O(N__46344),
            .I(N__46341));
    Odrv12 I__7728 (
            .O(N__46341),
            .I(\pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ));
    InMux I__7727 (
            .O(N__46338),
            .I(N__46335));
    LocalMux I__7726 (
            .O(N__46335),
            .I(N__46332));
    Span4Mux_h I__7725 (
            .O(N__46332),
            .I(N__46327));
    InMux I__7724 (
            .O(N__46331),
            .I(N__46324));
    InMux I__7723 (
            .O(N__46330),
            .I(N__46321));
    Odrv4 I__7722 (
            .O(N__46327),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    LocalMux I__7721 (
            .O(N__46324),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    LocalMux I__7720 (
            .O(N__46321),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    InMux I__7719 (
            .O(N__46314),
            .I(N__46311));
    LocalMux I__7718 (
            .O(N__46311),
            .I(N__46306));
    InMux I__7717 (
            .O(N__46310),
            .I(N__46301));
    InMux I__7716 (
            .O(N__46309),
            .I(N__46301));
    Odrv4 I__7715 (
            .O(N__46306),
            .I(\pid_front.un1_pid_prereg_0_9 ));
    LocalMux I__7714 (
            .O(N__46301),
            .I(\pid_front.un1_pid_prereg_0_9 ));
    InMux I__7713 (
            .O(N__46296),
            .I(N__46293));
    LocalMux I__7712 (
            .O(N__46293),
            .I(N__46289));
    InMux I__7711 (
            .O(N__46292),
            .I(N__46286));
    Odrv12 I__7710 (
            .O(N__46289),
            .I(\pid_front.un1_pid_prereg_0_8 ));
    LocalMux I__7709 (
            .O(N__46286),
            .I(\pid_front.un1_pid_prereg_0_8 ));
    CascadeMux I__7708 (
            .O(N__46281),
            .I(\pid_front.un1_pid_prereg_0_10_cascade_ ));
    InMux I__7707 (
            .O(N__46278),
            .I(N__46275));
    LocalMux I__7706 (
            .O(N__46275),
            .I(N__46272));
    Odrv4 I__7705 (
            .O(N__46272),
            .I(\pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ));
    CascadeMux I__7704 (
            .O(N__46269),
            .I(N__46266));
    InMux I__7703 (
            .O(N__46266),
            .I(N__46263));
    LocalMux I__7702 (
            .O(N__46263),
            .I(N__46260));
    Span4Mux_h I__7701 (
            .O(N__46260),
            .I(N__46257));
    Odrv4 I__7700 (
            .O(N__46257),
            .I(\pid_front.pid_preregZ0Z_27 ));
    InMux I__7699 (
            .O(N__46254),
            .I(\pid_front.un1_pid_prereg_0_cry_26 ));
    InMux I__7698 (
            .O(N__46251),
            .I(N__46248));
    LocalMux I__7697 (
            .O(N__46248),
            .I(N__46245));
    Span4Mux_v I__7696 (
            .O(N__46245),
            .I(N__46242));
    Odrv4 I__7695 (
            .O(N__46242),
            .I(\pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ));
    InMux I__7694 (
            .O(N__46239),
            .I(N__46236));
    LocalMux I__7693 (
            .O(N__46236),
            .I(N__46233));
    Span4Mux_h I__7692 (
            .O(N__46233),
            .I(N__46230));
    Odrv4 I__7691 (
            .O(N__46230),
            .I(\pid_front.pid_preregZ0Z_28 ));
    InMux I__7690 (
            .O(N__46227),
            .I(\pid_front.un1_pid_prereg_0_cry_27 ));
    InMux I__7689 (
            .O(N__46224),
            .I(N__46221));
    LocalMux I__7688 (
            .O(N__46221),
            .I(N__46218));
    Span4Mux_h I__7687 (
            .O(N__46218),
            .I(N__46215));
    Odrv4 I__7686 (
            .O(N__46215),
            .I(\pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ));
    CascadeMux I__7685 (
            .O(N__46212),
            .I(N__46209));
    InMux I__7684 (
            .O(N__46209),
            .I(N__46206));
    LocalMux I__7683 (
            .O(N__46206),
            .I(N__46203));
    Span4Mux_v I__7682 (
            .O(N__46203),
            .I(N__46200));
    Odrv4 I__7681 (
            .O(N__46200),
            .I(\pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ));
    InMux I__7680 (
            .O(N__46197),
            .I(N__46194));
    LocalMux I__7679 (
            .O(N__46194),
            .I(N__46191));
    Span4Mux_v I__7678 (
            .O(N__46191),
            .I(N__46188));
    Odrv4 I__7677 (
            .O(N__46188),
            .I(\pid_front.pid_preregZ0Z_29 ));
    InMux I__7676 (
            .O(N__46185),
            .I(\pid_front.un1_pid_prereg_0_cry_28 ));
    InMux I__7675 (
            .O(N__46182),
            .I(N__46179));
    LocalMux I__7674 (
            .O(N__46179),
            .I(N__46176));
    Span4Mux_v I__7673 (
            .O(N__46176),
            .I(N__46173));
    Odrv4 I__7672 (
            .O(N__46173),
            .I(\pid_front.un1_pid_prereg_0_axb_30 ));
    InMux I__7671 (
            .O(N__46170),
            .I(\pid_front.un1_pid_prereg_0_cry_29 ));
    CascadeMux I__7670 (
            .O(N__46167),
            .I(N__46161));
    CascadeMux I__7669 (
            .O(N__46166),
            .I(N__46158));
    CascadeMux I__7668 (
            .O(N__46165),
            .I(N__46146));
    CascadeMux I__7667 (
            .O(N__46164),
            .I(N__46143));
    InMux I__7666 (
            .O(N__46161),
            .I(N__46126));
    InMux I__7665 (
            .O(N__46158),
            .I(N__46126));
    InMux I__7664 (
            .O(N__46157),
            .I(N__46126));
    InMux I__7663 (
            .O(N__46156),
            .I(N__46126));
    InMux I__7662 (
            .O(N__46155),
            .I(N__46126));
    InMux I__7661 (
            .O(N__46154),
            .I(N__46126));
    InMux I__7660 (
            .O(N__46153),
            .I(N__46126));
    InMux I__7659 (
            .O(N__46152),
            .I(N__46126));
    CascadeMux I__7658 (
            .O(N__46151),
            .I(N__46119));
    InMux I__7657 (
            .O(N__46150),
            .I(N__46109));
    InMux I__7656 (
            .O(N__46149),
            .I(N__46109));
    InMux I__7655 (
            .O(N__46146),
            .I(N__46109));
    InMux I__7654 (
            .O(N__46143),
            .I(N__46109));
    LocalMux I__7653 (
            .O(N__46126),
            .I(N__46106));
    InMux I__7652 (
            .O(N__46125),
            .I(N__46097));
    InMux I__7651 (
            .O(N__46124),
            .I(N__46097));
    InMux I__7650 (
            .O(N__46123),
            .I(N__46097));
    InMux I__7649 (
            .O(N__46122),
            .I(N__46097));
    InMux I__7648 (
            .O(N__46119),
            .I(N__46092));
    InMux I__7647 (
            .O(N__46118),
            .I(N__46092));
    LocalMux I__7646 (
            .O(N__46109),
            .I(N__46083));
    Span4Mux_h I__7645 (
            .O(N__46106),
            .I(N__46083));
    LocalMux I__7644 (
            .O(N__46097),
            .I(N__46083));
    LocalMux I__7643 (
            .O(N__46092),
            .I(N__46083));
    Span4Mux_v I__7642 (
            .O(N__46083),
            .I(N__46080));
    Odrv4 I__7641 (
            .O(N__46080),
            .I(\pid_front.pid_preregZ0Z_30 ));
    InMux I__7640 (
            .O(N__46077),
            .I(N__46073));
    InMux I__7639 (
            .O(N__46076),
            .I(N__46070));
    LocalMux I__7638 (
            .O(N__46073),
            .I(N__46056));
    LocalMux I__7637 (
            .O(N__46070),
            .I(N__46053));
    CEMux I__7636 (
            .O(N__46069),
            .I(N__46026));
    CEMux I__7635 (
            .O(N__46068),
            .I(N__46026));
    CEMux I__7634 (
            .O(N__46067),
            .I(N__46026));
    CEMux I__7633 (
            .O(N__46066),
            .I(N__46026));
    CEMux I__7632 (
            .O(N__46065),
            .I(N__46026));
    CEMux I__7631 (
            .O(N__46064),
            .I(N__46026));
    CEMux I__7630 (
            .O(N__46063),
            .I(N__46026));
    CEMux I__7629 (
            .O(N__46062),
            .I(N__46026));
    CEMux I__7628 (
            .O(N__46061),
            .I(N__46026));
    CEMux I__7627 (
            .O(N__46060),
            .I(N__46026));
    CEMux I__7626 (
            .O(N__46059),
            .I(N__46026));
    Glb2LocalMux I__7625 (
            .O(N__46056),
            .I(N__46026));
    Glb2LocalMux I__7624 (
            .O(N__46053),
            .I(N__46026));
    GlobalMux I__7623 (
            .O(N__46026),
            .I(N__46023));
    gio2CtrlBuf I__7622 (
            .O(N__46023),
            .I(\pid_front.N_404_g ));
    CascadeMux I__7621 (
            .O(N__46020),
            .I(N__46017));
    InMux I__7620 (
            .O(N__46017),
            .I(N__46014));
    LocalMux I__7619 (
            .O(N__46014),
            .I(\pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ));
    InMux I__7618 (
            .O(N__46011),
            .I(N__46008));
    LocalMux I__7617 (
            .O(N__46008),
            .I(N__46003));
    InMux I__7616 (
            .O(N__46007),
            .I(N__46000));
    InMux I__7615 (
            .O(N__46006),
            .I(N__45997));
    Odrv4 I__7614 (
            .O(N__46003),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    LocalMux I__7613 (
            .O(N__46000),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    LocalMux I__7612 (
            .O(N__45997),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    InMux I__7611 (
            .O(N__45990),
            .I(N__45987));
    LocalMux I__7610 (
            .O(N__45987),
            .I(N__45984));
    Span4Mux_h I__7609 (
            .O(N__45984),
            .I(N__45980));
    InMux I__7608 (
            .O(N__45983),
            .I(N__45977));
    Odrv4 I__7607 (
            .O(N__45980),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    LocalMux I__7606 (
            .O(N__45977),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    CascadeMux I__7605 (
            .O(N__45972),
            .I(\pid_front.un1_pid_prereg_0_15_cascade_ ));
    InMux I__7604 (
            .O(N__45969),
            .I(N__45966));
    LocalMux I__7603 (
            .O(N__45966),
            .I(\pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ));
    CascadeMux I__7602 (
            .O(N__45963),
            .I(N__45960));
    InMux I__7601 (
            .O(N__45960),
            .I(N__45957));
    LocalMux I__7600 (
            .O(N__45957),
            .I(N__45954));
    Odrv4 I__7599 (
            .O(N__45954),
            .I(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ));
    InMux I__7598 (
            .O(N__45951),
            .I(N__45948));
    LocalMux I__7597 (
            .O(N__45948),
            .I(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ));
    CascadeMux I__7596 (
            .O(N__45945),
            .I(N__45941));
    InMux I__7595 (
            .O(N__45944),
            .I(N__45936));
    InMux I__7594 (
            .O(N__45941),
            .I(N__45936));
    LocalMux I__7593 (
            .O(N__45936),
            .I(N__45933));
    Span4Mux_h I__7592 (
            .O(N__45933),
            .I(N__45930));
    Odrv4 I__7591 (
            .O(N__45930),
            .I(\pid_front.pid_preregZ0Z_19 ));
    InMux I__7590 (
            .O(N__45927),
            .I(\pid_front.un1_pid_prereg_0_cry_18 ));
    CascadeMux I__7589 (
            .O(N__45924),
            .I(N__45921));
    InMux I__7588 (
            .O(N__45921),
            .I(N__45918));
    LocalMux I__7587 (
            .O(N__45918),
            .I(N__45915));
    Odrv4 I__7586 (
            .O(N__45915),
            .I(\pid_front.pid_preregZ0Z_20 ));
    InMux I__7585 (
            .O(N__45912),
            .I(\pid_front.un1_pid_prereg_0_cry_19 ));
    InMux I__7584 (
            .O(N__45909),
            .I(N__45906));
    LocalMux I__7583 (
            .O(N__45906),
            .I(N__45903));
    Odrv4 I__7582 (
            .O(N__45903),
            .I(\pid_front.pid_preregZ0Z_21 ));
    InMux I__7581 (
            .O(N__45900),
            .I(\pid_front.un1_pid_prereg_0_cry_20 ));
    InMux I__7580 (
            .O(N__45897),
            .I(N__45894));
    LocalMux I__7579 (
            .O(N__45894),
            .I(N__45891));
    Odrv4 I__7578 (
            .O(N__45891),
            .I(\pid_front.pid_preregZ0Z_22 ));
    InMux I__7577 (
            .O(N__45888),
            .I(\pid_front.un1_pid_prereg_0_cry_21 ));
    InMux I__7576 (
            .O(N__45885),
            .I(N__45882));
    LocalMux I__7575 (
            .O(N__45882),
            .I(N__45879));
    Odrv4 I__7574 (
            .O(N__45879),
            .I(\pid_front.pid_preregZ0Z_23 ));
    InMux I__7573 (
            .O(N__45876),
            .I(bfn_11_18_0_));
    InMux I__7572 (
            .O(N__45873),
            .I(N__45870));
    LocalMux I__7571 (
            .O(N__45870),
            .I(N__45867));
    Span4Mux_h I__7570 (
            .O(N__45867),
            .I(N__45864));
    Odrv4 I__7569 (
            .O(N__45864),
            .I(\pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ));
    InMux I__7568 (
            .O(N__45861),
            .I(N__45858));
    LocalMux I__7567 (
            .O(N__45858),
            .I(N__45855));
    Span4Mux_h I__7566 (
            .O(N__45855),
            .I(N__45852));
    Odrv4 I__7565 (
            .O(N__45852),
            .I(\pid_front.pid_preregZ0Z_24 ));
    InMux I__7564 (
            .O(N__45849),
            .I(\pid_front.un1_pid_prereg_0_cry_23 ));
    InMux I__7563 (
            .O(N__45846),
            .I(N__45843));
    LocalMux I__7562 (
            .O(N__45843),
            .I(N__45840));
    Span4Mux_v I__7561 (
            .O(N__45840),
            .I(N__45837));
    Odrv4 I__7560 (
            .O(N__45837),
            .I(\pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ));
    CascadeMux I__7559 (
            .O(N__45834),
            .I(N__45831));
    InMux I__7558 (
            .O(N__45831),
            .I(N__45828));
    LocalMux I__7557 (
            .O(N__45828),
            .I(N__45825));
    Span4Mux_h I__7556 (
            .O(N__45825),
            .I(N__45822));
    Odrv4 I__7555 (
            .O(N__45822),
            .I(\pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ));
    InMux I__7554 (
            .O(N__45819),
            .I(N__45816));
    LocalMux I__7553 (
            .O(N__45816),
            .I(N__45813));
    Span4Mux_h I__7552 (
            .O(N__45813),
            .I(N__45810));
    Odrv4 I__7551 (
            .O(N__45810),
            .I(\pid_front.pid_preregZ0Z_25 ));
    InMux I__7550 (
            .O(N__45807),
            .I(\pid_front.un1_pid_prereg_0_cry_24 ));
    CascadeMux I__7549 (
            .O(N__45804),
            .I(N__45801));
    InMux I__7548 (
            .O(N__45801),
            .I(N__45798));
    LocalMux I__7547 (
            .O(N__45798),
            .I(N__45795));
    Span4Mux_h I__7546 (
            .O(N__45795),
            .I(N__45792));
    Odrv4 I__7545 (
            .O(N__45792),
            .I(\pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ));
    InMux I__7544 (
            .O(N__45789),
            .I(N__45786));
    LocalMux I__7543 (
            .O(N__45786),
            .I(N__45783));
    Span4Mux_h I__7542 (
            .O(N__45783),
            .I(N__45780));
    Odrv4 I__7541 (
            .O(N__45780),
            .I(\pid_front.pid_preregZ0Z_26 ));
    InMux I__7540 (
            .O(N__45777),
            .I(\pid_front.un1_pid_prereg_0_cry_25 ));
    CascadeMux I__7539 (
            .O(N__45774),
            .I(N__45769));
    CascadeMux I__7538 (
            .O(N__45773),
            .I(N__45766));
    InMux I__7537 (
            .O(N__45772),
            .I(N__45763));
    InMux I__7536 (
            .O(N__45769),
            .I(N__45758));
    InMux I__7535 (
            .O(N__45766),
            .I(N__45758));
    LocalMux I__7534 (
            .O(N__45763),
            .I(N__45755));
    LocalMux I__7533 (
            .O(N__45758),
            .I(N__45752));
    Odrv12 I__7532 (
            .O(N__45755),
            .I(\pid_front.pid_preregZ0Z_11 ));
    Odrv4 I__7531 (
            .O(N__45752),
            .I(\pid_front.pid_preregZ0Z_11 ));
    InMux I__7530 (
            .O(N__45747),
            .I(\pid_front.un1_pid_prereg_0_cry_10 ));
    InMux I__7529 (
            .O(N__45744),
            .I(N__45737));
    InMux I__7528 (
            .O(N__45743),
            .I(N__45734));
    InMux I__7527 (
            .O(N__45742),
            .I(N__45731));
    InMux I__7526 (
            .O(N__45741),
            .I(N__45728));
    InMux I__7525 (
            .O(N__45740),
            .I(N__45725));
    LocalMux I__7524 (
            .O(N__45737),
            .I(N__45720));
    LocalMux I__7523 (
            .O(N__45734),
            .I(N__45720));
    LocalMux I__7522 (
            .O(N__45731),
            .I(N__45717));
    LocalMux I__7521 (
            .O(N__45728),
            .I(N__45712));
    LocalMux I__7520 (
            .O(N__45725),
            .I(N__45712));
    Span4Mux_h I__7519 (
            .O(N__45720),
            .I(N__45709));
    Odrv12 I__7518 (
            .O(N__45717),
            .I(\pid_front.pid_preregZ0Z_12 ));
    Odrv4 I__7517 (
            .O(N__45712),
            .I(\pid_front.pid_preregZ0Z_12 ));
    Odrv4 I__7516 (
            .O(N__45709),
            .I(\pid_front.pid_preregZ0Z_12 ));
    InMux I__7515 (
            .O(N__45702),
            .I(\pid_front.un1_pid_prereg_0_cry_11 ));
    CascadeMux I__7514 (
            .O(N__45699),
            .I(N__45696));
    InMux I__7513 (
            .O(N__45696),
            .I(N__45686));
    InMux I__7512 (
            .O(N__45695),
            .I(N__45686));
    InMux I__7511 (
            .O(N__45694),
            .I(N__45683));
    InMux I__7510 (
            .O(N__45693),
            .I(N__45678));
    InMux I__7509 (
            .O(N__45692),
            .I(N__45678));
    InMux I__7508 (
            .O(N__45691),
            .I(N__45675));
    LocalMux I__7507 (
            .O(N__45686),
            .I(N__45670));
    LocalMux I__7506 (
            .O(N__45683),
            .I(N__45670));
    LocalMux I__7505 (
            .O(N__45678),
            .I(N__45667));
    LocalMux I__7504 (
            .O(N__45675),
            .I(N__45664));
    Span4Mux_v I__7503 (
            .O(N__45670),
            .I(N__45659));
    Span4Mux_h I__7502 (
            .O(N__45667),
            .I(N__45659));
    Odrv4 I__7501 (
            .O(N__45664),
            .I(\pid_front.pid_preregZ0Z_13 ));
    Odrv4 I__7500 (
            .O(N__45659),
            .I(\pid_front.pid_preregZ0Z_13 ));
    InMux I__7499 (
            .O(N__45654),
            .I(\pid_front.un1_pid_prereg_0_cry_12 ));
    InMux I__7498 (
            .O(N__45651),
            .I(N__45647));
    InMux I__7497 (
            .O(N__45650),
            .I(N__45644));
    LocalMux I__7496 (
            .O(N__45647),
            .I(\pid_front.un1_pid_prereg_0_axb_14 ));
    LocalMux I__7495 (
            .O(N__45644),
            .I(\pid_front.un1_pid_prereg_0_axb_14 ));
    InMux I__7494 (
            .O(N__45639),
            .I(N__45636));
    LocalMux I__7493 (
            .O(N__45636),
            .I(N__45633));
    Span4Mux_h I__7492 (
            .O(N__45633),
            .I(N__45630));
    Odrv4 I__7491 (
            .O(N__45630),
            .I(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__7490 (
            .O(N__45627),
            .I(\pid_front.un1_pid_prereg_0_cry_13 ));
    CascadeMux I__7489 (
            .O(N__45624),
            .I(N__45620));
    InMux I__7488 (
            .O(N__45623),
            .I(N__45615));
    InMux I__7487 (
            .O(N__45620),
            .I(N__45615));
    LocalMux I__7486 (
            .O(N__45615),
            .I(N__45612));
    Span4Mux_h I__7485 (
            .O(N__45612),
            .I(N__45609));
    Odrv4 I__7484 (
            .O(N__45609),
            .I(\pid_front.pid_preregZ0Z_15 ));
    InMux I__7483 (
            .O(N__45606),
            .I(bfn_11_17_0_));
    InMux I__7482 (
            .O(N__45603),
            .I(N__45597));
    InMux I__7481 (
            .O(N__45602),
            .I(N__45597));
    LocalMux I__7480 (
            .O(N__45597),
            .I(N__45594));
    Span4Mux_h I__7479 (
            .O(N__45594),
            .I(N__45591));
    Odrv4 I__7478 (
            .O(N__45591),
            .I(\pid_front.pid_preregZ0Z_16 ));
    InMux I__7477 (
            .O(N__45588),
            .I(\pid_front.un1_pid_prereg_0_cry_15 ));
    InMux I__7476 (
            .O(N__45585),
            .I(N__45582));
    LocalMux I__7475 (
            .O(N__45582),
            .I(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ));
    InMux I__7474 (
            .O(N__45579),
            .I(N__45573));
    InMux I__7473 (
            .O(N__45578),
            .I(N__45573));
    LocalMux I__7472 (
            .O(N__45573),
            .I(N__45570));
    Span4Mux_v I__7471 (
            .O(N__45570),
            .I(N__45567));
    Odrv4 I__7470 (
            .O(N__45567),
            .I(\pid_front.pid_preregZ0Z_17 ));
    InMux I__7469 (
            .O(N__45564),
            .I(\pid_front.un1_pid_prereg_0_cry_16 ));
    InMux I__7468 (
            .O(N__45561),
            .I(N__45558));
    LocalMux I__7467 (
            .O(N__45558),
            .I(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ));
    CascadeMux I__7466 (
            .O(N__45555),
            .I(N__45552));
    InMux I__7465 (
            .O(N__45552),
            .I(N__45549));
    LocalMux I__7464 (
            .O(N__45549),
            .I(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ));
    InMux I__7463 (
            .O(N__45546),
            .I(N__45540));
    InMux I__7462 (
            .O(N__45545),
            .I(N__45540));
    LocalMux I__7461 (
            .O(N__45540),
            .I(N__45537));
    Span4Mux_v I__7460 (
            .O(N__45537),
            .I(N__45534));
    Span4Mux_h I__7459 (
            .O(N__45534),
            .I(N__45531));
    Odrv4 I__7458 (
            .O(N__45531),
            .I(\pid_front.pid_preregZ0Z_18 ));
    InMux I__7457 (
            .O(N__45528),
            .I(\pid_front.un1_pid_prereg_0_cry_17 ));
    CascadeMux I__7456 (
            .O(N__45525),
            .I(N__45521));
    CascadeMux I__7455 (
            .O(N__45524),
            .I(N__45517));
    InMux I__7454 (
            .O(N__45521),
            .I(N__45514));
    InMux I__7453 (
            .O(N__45520),
            .I(N__45509));
    InMux I__7452 (
            .O(N__45517),
            .I(N__45509));
    LocalMux I__7451 (
            .O(N__45514),
            .I(N__45504));
    LocalMux I__7450 (
            .O(N__45509),
            .I(N__45504));
    Odrv4 I__7449 (
            .O(N__45504),
            .I(\pid_front.pid_preregZ0Z_3 ));
    InMux I__7448 (
            .O(N__45501),
            .I(\pid_front.un1_pid_prereg_0_cry_2 ));
    InMux I__7447 (
            .O(N__45498),
            .I(N__45495));
    LocalMux I__7446 (
            .O(N__45495),
            .I(N__45492));
    Span4Mux_h I__7445 (
            .O(N__45492),
            .I(N__45489));
    Odrv4 I__7444 (
            .O(N__45489),
            .I(\pid_front.error_p_reg_esr_RNI4U472Z0Z_3 ));
    InMux I__7443 (
            .O(N__45486),
            .I(N__45481));
    InMux I__7442 (
            .O(N__45485),
            .I(N__45475));
    InMux I__7441 (
            .O(N__45484),
            .I(N__45475));
    LocalMux I__7440 (
            .O(N__45481),
            .I(N__45472));
    InMux I__7439 (
            .O(N__45480),
            .I(N__45469));
    LocalMux I__7438 (
            .O(N__45475),
            .I(\pid_front.pid_preregZ0Z_4 ));
    Odrv4 I__7437 (
            .O(N__45472),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__7436 (
            .O(N__45469),
            .I(\pid_front.pid_preregZ0Z_4 ));
    InMux I__7435 (
            .O(N__45462),
            .I(\pid_front.un1_pid_prereg_0_cry_3 ));
    InMux I__7434 (
            .O(N__45459),
            .I(N__45455));
    CascadeMux I__7433 (
            .O(N__45458),
            .I(N__45452));
    LocalMux I__7432 (
            .O(N__45455),
            .I(N__45449));
    InMux I__7431 (
            .O(N__45452),
            .I(N__45446));
    Span4Mux_h I__7430 (
            .O(N__45449),
            .I(N__45443));
    LocalMux I__7429 (
            .O(N__45446),
            .I(\pid_front.error_p_reg_esr_RNIKJHV_0Z0Z_5 ));
    Odrv4 I__7428 (
            .O(N__45443),
            .I(\pid_front.error_p_reg_esr_RNIKJHV_0Z0Z_5 ));
    CascadeMux I__7427 (
            .O(N__45438),
            .I(N__45435));
    InMux I__7426 (
            .O(N__45435),
            .I(N__45432));
    LocalMux I__7425 (
            .O(N__45432),
            .I(N__45429));
    Span4Mux_h I__7424 (
            .O(N__45429),
            .I(N__45426));
    Odrv4 I__7423 (
            .O(N__45426),
            .I(\pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ));
    InMux I__7422 (
            .O(N__45423),
            .I(N__45417));
    CascadeMux I__7421 (
            .O(N__45422),
            .I(N__45414));
    InMux I__7420 (
            .O(N__45421),
            .I(N__45409));
    InMux I__7419 (
            .O(N__45420),
            .I(N__45409));
    LocalMux I__7418 (
            .O(N__45417),
            .I(N__45406));
    InMux I__7417 (
            .O(N__45414),
            .I(N__45403));
    LocalMux I__7416 (
            .O(N__45409),
            .I(\pid_front.pid_preregZ0Z_5 ));
    Odrv12 I__7415 (
            .O(N__45406),
            .I(\pid_front.pid_preregZ0Z_5 ));
    LocalMux I__7414 (
            .O(N__45403),
            .I(\pid_front.pid_preregZ0Z_5 ));
    InMux I__7413 (
            .O(N__45396),
            .I(\pid_front.un1_pid_prereg_0_cry_4 ));
    InMux I__7412 (
            .O(N__45393),
            .I(N__45390));
    LocalMux I__7411 (
            .O(N__45390),
            .I(N__45387));
    Span4Mux_v I__7410 (
            .O(N__45387),
            .I(N__45384));
    Odrv4 I__7409 (
            .O(N__45384),
            .I(\pid_front.error_p_reg_esr_RNIHMAE2Z0Z_5 ));
    CascadeMux I__7408 (
            .O(N__45381),
            .I(N__45378));
    InMux I__7407 (
            .O(N__45378),
            .I(N__45375));
    LocalMux I__7406 (
            .O(N__45375),
            .I(N__45372));
    Span4Mux_h I__7405 (
            .O(N__45372),
            .I(N__45369));
    Odrv4 I__7404 (
            .O(N__45369),
            .I(\pid_front.error_p_reg_esr_RNIKJHVZ0Z_5 ));
    InMux I__7403 (
            .O(N__45366),
            .I(N__45363));
    LocalMux I__7402 (
            .O(N__45363),
            .I(N__45358));
    InMux I__7401 (
            .O(N__45362),
            .I(N__45355));
    InMux I__7400 (
            .O(N__45361),
            .I(N__45352));
    Odrv12 I__7399 (
            .O(N__45358),
            .I(\pid_front.pid_preregZ0Z_6 ));
    LocalMux I__7398 (
            .O(N__45355),
            .I(\pid_front.pid_preregZ0Z_6 ));
    LocalMux I__7397 (
            .O(N__45352),
            .I(\pid_front.pid_preregZ0Z_6 ));
    InMux I__7396 (
            .O(N__45345),
            .I(\pid_front.un1_pid_prereg_0_cry_5 ));
    InMux I__7395 (
            .O(N__45342),
            .I(N__45339));
    LocalMux I__7394 (
            .O(N__45339),
            .I(N__45336));
    Odrv4 I__7393 (
            .O(N__45336),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ));
    CascadeMux I__7392 (
            .O(N__45333),
            .I(N__45330));
    InMux I__7391 (
            .O(N__45330),
            .I(N__45327));
    LocalMux I__7390 (
            .O(N__45327),
            .I(N__45324));
    Span4Mux_v I__7389 (
            .O(N__45324),
            .I(N__45321));
    Span4Mux_h I__7388 (
            .O(N__45321),
            .I(N__45318));
    Odrv4 I__7387 (
            .O(N__45318),
            .I(\pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ));
    InMux I__7386 (
            .O(N__45315),
            .I(N__45310));
    InMux I__7385 (
            .O(N__45314),
            .I(N__45307));
    InMux I__7384 (
            .O(N__45313),
            .I(N__45304));
    LocalMux I__7383 (
            .O(N__45310),
            .I(N__45301));
    LocalMux I__7382 (
            .O(N__45307),
            .I(N__45296));
    LocalMux I__7381 (
            .O(N__45304),
            .I(N__45296));
    Odrv12 I__7380 (
            .O(N__45301),
            .I(\pid_front.pid_preregZ0Z_7 ));
    Odrv4 I__7379 (
            .O(N__45296),
            .I(\pid_front.pid_preregZ0Z_7 ));
    InMux I__7378 (
            .O(N__45291),
            .I(bfn_11_16_0_));
    InMux I__7377 (
            .O(N__45288),
            .I(N__45285));
    LocalMux I__7376 (
            .O(N__45285),
            .I(N__45282));
    Odrv4 I__7375 (
            .O(N__45282),
            .I(\pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ));
    CascadeMux I__7374 (
            .O(N__45279),
            .I(N__45276));
    InMux I__7373 (
            .O(N__45276),
            .I(N__45273));
    LocalMux I__7372 (
            .O(N__45273),
            .I(N__45269));
    InMux I__7371 (
            .O(N__45272),
            .I(N__45266));
    Span4Mux_h I__7370 (
            .O(N__45269),
            .I(N__45263));
    LocalMux I__7369 (
            .O(N__45266),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ));
    Odrv4 I__7368 (
            .O(N__45263),
            .I(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ));
    InMux I__7367 (
            .O(N__45258),
            .I(N__45253));
    InMux I__7366 (
            .O(N__45257),
            .I(N__45248));
    InMux I__7365 (
            .O(N__45256),
            .I(N__45248));
    LocalMux I__7364 (
            .O(N__45253),
            .I(N__45245));
    LocalMux I__7363 (
            .O(N__45248),
            .I(N__45242));
    Odrv12 I__7362 (
            .O(N__45245),
            .I(\pid_front.pid_preregZ0Z_8 ));
    Odrv4 I__7361 (
            .O(N__45242),
            .I(\pid_front.pid_preregZ0Z_8 ));
    InMux I__7360 (
            .O(N__45237),
            .I(\pid_front.un1_pid_prereg_0_cry_7 ));
    InMux I__7359 (
            .O(N__45234),
            .I(N__45229));
    InMux I__7358 (
            .O(N__45233),
            .I(N__45224));
    InMux I__7357 (
            .O(N__45232),
            .I(N__45224));
    LocalMux I__7356 (
            .O(N__45229),
            .I(N__45221));
    LocalMux I__7355 (
            .O(N__45224),
            .I(N__45218));
    Odrv12 I__7354 (
            .O(N__45221),
            .I(\pid_front.pid_preregZ0Z_9 ));
    Odrv4 I__7353 (
            .O(N__45218),
            .I(\pid_front.pid_preregZ0Z_9 ));
    InMux I__7352 (
            .O(N__45213),
            .I(\pid_front.un1_pid_prereg_0_cry_8 ));
    InMux I__7351 (
            .O(N__45210),
            .I(N__45205));
    InMux I__7350 (
            .O(N__45209),
            .I(N__45200));
    InMux I__7349 (
            .O(N__45208),
            .I(N__45200));
    LocalMux I__7348 (
            .O(N__45205),
            .I(N__45197));
    LocalMux I__7347 (
            .O(N__45200),
            .I(N__45194));
    Odrv12 I__7346 (
            .O(N__45197),
            .I(\pid_front.pid_preregZ0Z_10 ));
    Odrv4 I__7345 (
            .O(N__45194),
            .I(\pid_front.pid_preregZ0Z_10 ));
    InMux I__7344 (
            .O(N__45189),
            .I(\pid_front.un1_pid_prereg_0_cry_9 ));
    InMux I__7343 (
            .O(N__45186),
            .I(N__45180));
    InMux I__7342 (
            .O(N__45185),
            .I(N__45180));
    LocalMux I__7341 (
            .O(N__45180),
            .I(N__45176));
    InMux I__7340 (
            .O(N__45179),
            .I(N__45173));
    Odrv4 I__7339 (
            .O(N__45176),
            .I(\pid_front.N_98 ));
    LocalMux I__7338 (
            .O(N__45173),
            .I(\pid_front.N_98 ));
    InMux I__7337 (
            .O(N__45168),
            .I(N__45165));
    LocalMux I__7336 (
            .O(N__45165),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_o2_sx ));
    CascadeMux I__7335 (
            .O(N__45162),
            .I(\pid_front.N_75_cascade_ ));
    InMux I__7334 (
            .O(N__45159),
            .I(N__45156));
    LocalMux I__7333 (
            .O(N__45156),
            .I(\pid_front.N_102 ));
    InMux I__7332 (
            .O(N__45153),
            .I(N__45149));
    CascadeMux I__7331 (
            .O(N__45152),
            .I(N__45146));
    LocalMux I__7330 (
            .O(N__45149),
            .I(N__45143));
    InMux I__7329 (
            .O(N__45146),
            .I(N__45140));
    Span4Mux_h I__7328 (
            .O(N__45143),
            .I(N__45137));
    LocalMux I__7327 (
            .O(N__45140),
            .I(\pid_front.N_99 ));
    Odrv4 I__7326 (
            .O(N__45137),
            .I(\pid_front.N_99 ));
    InMux I__7325 (
            .O(N__45132),
            .I(N__45129));
    LocalMux I__7324 (
            .O(N__45129),
            .I(\pid_front.N_11_i ));
    CascadeMux I__7323 (
            .O(N__45126),
            .I(N__45120));
    CascadeMux I__7322 (
            .O(N__45125),
            .I(N__45117));
    InMux I__7321 (
            .O(N__45124),
            .I(N__45100));
    InMux I__7320 (
            .O(N__45123),
            .I(N__45100));
    InMux I__7319 (
            .O(N__45120),
            .I(N__45100));
    InMux I__7318 (
            .O(N__45117),
            .I(N__45100));
    InMux I__7317 (
            .O(N__45116),
            .I(N__45095));
    InMux I__7316 (
            .O(N__45115),
            .I(N__45095));
    InMux I__7315 (
            .O(N__45114),
            .I(N__45082));
    InMux I__7314 (
            .O(N__45113),
            .I(N__45082));
    InMux I__7313 (
            .O(N__45112),
            .I(N__45082));
    InMux I__7312 (
            .O(N__45111),
            .I(N__45082));
    InMux I__7311 (
            .O(N__45110),
            .I(N__45082));
    InMux I__7310 (
            .O(N__45109),
            .I(N__45082));
    LocalMux I__7309 (
            .O(N__45100),
            .I(N__45079));
    LocalMux I__7308 (
            .O(N__45095),
            .I(N__45074));
    LocalMux I__7307 (
            .O(N__45082),
            .I(N__45074));
    Span4Mux_h I__7306 (
            .O(N__45079),
            .I(N__45071));
    Span4Mux_v I__7305 (
            .O(N__45074),
            .I(N__45068));
    Odrv4 I__7304 (
            .O(N__45071),
            .I(\pid_front.N_76 ));
    Odrv4 I__7303 (
            .O(N__45068),
            .I(\pid_front.N_76 ));
    CascadeMux I__7302 (
            .O(N__45063),
            .I(N__45058));
    InMux I__7301 (
            .O(N__45062),
            .I(N__45051));
    InMux I__7300 (
            .O(N__45061),
            .I(N__45051));
    InMux I__7299 (
            .O(N__45058),
            .I(N__45048));
    InMux I__7298 (
            .O(N__45057),
            .I(N__45043));
    InMux I__7297 (
            .O(N__45056),
            .I(N__45043));
    LocalMux I__7296 (
            .O(N__45051),
            .I(N__45040));
    LocalMux I__7295 (
            .O(N__45048),
            .I(\pid_front.N_75 ));
    LocalMux I__7294 (
            .O(N__45043),
            .I(\pid_front.N_75 ));
    Odrv4 I__7293 (
            .O(N__45040),
            .I(\pid_front.N_75 ));
    CascadeMux I__7292 (
            .O(N__45033),
            .I(N__45030));
    InMux I__7291 (
            .O(N__45030),
            .I(N__45026));
    InMux I__7290 (
            .O(N__45029),
            .I(N__45023));
    LocalMux I__7289 (
            .O(N__45026),
            .I(N__45020));
    LocalMux I__7288 (
            .O(N__45023),
            .I(N__45017));
    Span4Mux_v I__7287 (
            .O(N__45020),
            .I(N__45014));
    Span4Mux_v I__7286 (
            .O(N__45017),
            .I(N__45011));
    Span4Mux_h I__7285 (
            .O(N__45014),
            .I(N__45006));
    Span4Mux_h I__7284 (
            .O(N__45011),
            .I(N__45006));
    Odrv4 I__7283 (
            .O(N__45006),
            .I(\pid_front.error_p_regZ0Z_0 ));
    InMux I__7282 (
            .O(N__45003),
            .I(N__44994));
    InMux I__7281 (
            .O(N__45002),
            .I(N__44994));
    InMux I__7280 (
            .O(N__45001),
            .I(N__44994));
    LocalMux I__7279 (
            .O(N__44994),
            .I(N__44991));
    Odrv4 I__7278 (
            .O(N__44991),
            .I(\pid_front.pid_preregZ0Z_0 ));
    InMux I__7277 (
            .O(N__44988),
            .I(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__7276 (
            .O(N__44985),
            .I(N__44976));
    InMux I__7275 (
            .O(N__44984),
            .I(N__44976));
    InMux I__7274 (
            .O(N__44983),
            .I(N__44976));
    LocalMux I__7273 (
            .O(N__44976),
            .I(N__44973));
    Odrv4 I__7272 (
            .O(N__44973),
            .I(\pid_front.pid_preregZ0Z_1 ));
    InMux I__7271 (
            .O(N__44970),
            .I(\pid_front.un1_pid_prereg_0_cry_0 ));
    InMux I__7270 (
            .O(N__44967),
            .I(N__44958));
    InMux I__7269 (
            .O(N__44966),
            .I(N__44958));
    InMux I__7268 (
            .O(N__44965),
            .I(N__44958));
    LocalMux I__7267 (
            .O(N__44958),
            .I(N__44955));
    Odrv4 I__7266 (
            .O(N__44955),
            .I(\pid_front.pid_preregZ0Z_2 ));
    InMux I__7265 (
            .O(N__44952),
            .I(\pid_front.un1_pid_prereg_0_cry_1 ));
    InMux I__7264 (
            .O(N__44949),
            .I(N__44946));
    LocalMux I__7263 (
            .O(N__44946),
            .I(N__44943));
    Span4Mux_h I__7262 (
            .O(N__44943),
            .I(N__44940));
    Odrv4 I__7261 (
            .O(N__44940),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a4_4 ));
    InMux I__7260 (
            .O(N__44937),
            .I(N__44934));
    LocalMux I__7259 (
            .O(N__44934),
            .I(\pid_front.source_pid10lt4_0 ));
    InMux I__7258 (
            .O(N__44931),
            .I(N__44928));
    LocalMux I__7257 (
            .O(N__44928),
            .I(N__44925));
    Span4Mux_v I__7256 (
            .O(N__44925),
            .I(N__44922));
    Odrv4 I__7255 (
            .O(N__44922),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a4_3 ));
    CascadeMux I__7254 (
            .O(N__44919),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ));
    CascadeMux I__7253 (
            .O(N__44916),
            .I(\pid_front.N_99_cascade_ ));
    InMux I__7252 (
            .O(N__44913),
            .I(N__44908));
    InMux I__7251 (
            .O(N__44912),
            .I(N__44899));
    InMux I__7250 (
            .O(N__44911),
            .I(N__44899));
    LocalMux I__7249 (
            .O(N__44908),
            .I(N__44896));
    InMux I__7248 (
            .O(N__44907),
            .I(N__44887));
    InMux I__7247 (
            .O(N__44906),
            .I(N__44887));
    InMux I__7246 (
            .O(N__44905),
            .I(N__44887));
    InMux I__7245 (
            .O(N__44904),
            .I(N__44887));
    LocalMux I__7244 (
            .O(N__44899),
            .I(N__44880));
    Span4Mux_h I__7243 (
            .O(N__44896),
            .I(N__44875));
    LocalMux I__7242 (
            .O(N__44887),
            .I(N__44875));
    InMux I__7241 (
            .O(N__44886),
            .I(N__44866));
    InMux I__7240 (
            .O(N__44885),
            .I(N__44866));
    InMux I__7239 (
            .O(N__44884),
            .I(N__44866));
    InMux I__7238 (
            .O(N__44883),
            .I(N__44866));
    Odrv4 I__7237 (
            .O(N__44880),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__7236 (
            .O(N__44875),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__7235 (
            .O(N__44866),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    CascadeMux I__7234 (
            .O(N__44859),
            .I(N__44852));
    CascadeMux I__7233 (
            .O(N__44858),
            .I(N__44848));
    CascadeMux I__7232 (
            .O(N__44857),
            .I(N__44845));
    CascadeMux I__7231 (
            .O(N__44856),
            .I(N__44842));
    CascadeMux I__7230 (
            .O(N__44855),
            .I(N__44838));
    InMux I__7229 (
            .O(N__44852),
            .I(N__44833));
    InMux I__7228 (
            .O(N__44851),
            .I(N__44833));
    InMux I__7227 (
            .O(N__44848),
            .I(N__44830));
    InMux I__7226 (
            .O(N__44845),
            .I(N__44821));
    InMux I__7225 (
            .O(N__44842),
            .I(N__44821));
    InMux I__7224 (
            .O(N__44841),
            .I(N__44821));
    InMux I__7223 (
            .O(N__44838),
            .I(N__44821));
    LocalMux I__7222 (
            .O(N__44833),
            .I(N__44816));
    LocalMux I__7221 (
            .O(N__44830),
            .I(N__44811));
    LocalMux I__7220 (
            .O(N__44821),
            .I(N__44811));
    InMux I__7219 (
            .O(N__44820),
            .I(N__44806));
    InMux I__7218 (
            .O(N__44819),
            .I(N__44806));
    Odrv4 I__7217 (
            .O(N__44816),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__7216 (
            .O(N__44811),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__7215 (
            .O(N__44806),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__7214 (
            .O(N__44799),
            .I(N__44788));
    InMux I__7213 (
            .O(N__44798),
            .I(N__44788));
    InMux I__7212 (
            .O(N__44797),
            .I(N__44785));
    InMux I__7211 (
            .O(N__44796),
            .I(N__44776));
    InMux I__7210 (
            .O(N__44795),
            .I(N__44776));
    InMux I__7209 (
            .O(N__44794),
            .I(N__44776));
    InMux I__7208 (
            .O(N__44793),
            .I(N__44776));
    LocalMux I__7207 (
            .O(N__44788),
            .I(N__44770));
    LocalMux I__7206 (
            .O(N__44785),
            .I(N__44765));
    LocalMux I__7205 (
            .O(N__44776),
            .I(N__44765));
    InMux I__7204 (
            .O(N__44775),
            .I(N__44758));
    InMux I__7203 (
            .O(N__44774),
            .I(N__44758));
    InMux I__7202 (
            .O(N__44773),
            .I(N__44758));
    Odrv4 I__7201 (
            .O(N__44770),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__7200 (
            .O(N__44765),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__7199 (
            .O(N__44758),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__7198 (
            .O(N__44751),
            .I(N__44748));
    LocalMux I__7197 (
            .O(N__44748),
            .I(\uart_drone.data_Auxce_0_5 ));
    CascadeMux I__7196 (
            .O(N__44745),
            .I(N__44742));
    InMux I__7195 (
            .O(N__44742),
            .I(N__44736));
    InMux I__7194 (
            .O(N__44741),
            .I(N__44736));
    LocalMux I__7193 (
            .O(N__44736),
            .I(N__44733));
    Odrv4 I__7192 (
            .O(N__44733),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__7191 (
            .O(N__44730),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__7190 (
            .O(N__44727),
            .I(N__44724));
    LocalMux I__7189 (
            .O(N__44724),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__7188 (
            .O(N__44721),
            .I(N__44718));
    InMux I__7187 (
            .O(N__44718),
            .I(N__44712));
    InMux I__7186 (
            .O(N__44717),
            .I(N__44712));
    LocalMux I__7185 (
            .O(N__44712),
            .I(N__44709));
    Odrv4 I__7184 (
            .O(N__44709),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__7183 (
            .O(N__44706),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__7182 (
            .O(N__44703),
            .I(N__44700));
    LocalMux I__7181 (
            .O(N__44700),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__7180 (
            .O(N__44697),
            .I(N__44694));
    InMux I__7179 (
            .O(N__44694),
            .I(N__44688));
    InMux I__7178 (
            .O(N__44693),
            .I(N__44688));
    LocalMux I__7177 (
            .O(N__44688),
            .I(N__44685));
    Odrv4 I__7176 (
            .O(N__44685),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__7175 (
            .O(N__44682),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__7174 (
            .O(N__44679),
            .I(N__44676));
    LocalMux I__7173 (
            .O(N__44676),
            .I(N__44673));
    Span4Mux_h I__7172 (
            .O(N__44673),
            .I(N__44670));
    Span4Mux_v I__7171 (
            .O(N__44670),
            .I(N__44667));
    Odrv4 I__7170 (
            .O(N__44667),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    CascadeMux I__7169 (
            .O(N__44664),
            .I(N__44661));
    InMux I__7168 (
            .O(N__44661),
            .I(N__44655));
    InMux I__7167 (
            .O(N__44660),
            .I(N__44655));
    LocalMux I__7166 (
            .O(N__44655),
            .I(N__44652));
    Odrv4 I__7165 (
            .O(N__44652),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__7164 (
            .O(N__44649),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__7163 (
            .O(N__44646),
            .I(N__44642));
    InMux I__7162 (
            .O(N__44645),
            .I(N__44639));
    LocalMux I__7161 (
            .O(N__44642),
            .I(N__44634));
    LocalMux I__7160 (
            .O(N__44639),
            .I(N__44634));
    Odrv4 I__7159 (
            .O(N__44634),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    InMux I__7158 (
            .O(N__44631),
            .I(bfn_11_11_0_));
    InMux I__7157 (
            .O(N__44628),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CascadeMux I__7156 (
            .O(N__44625),
            .I(N__44622));
    InMux I__7155 (
            .O(N__44622),
            .I(N__44619));
    LocalMux I__7154 (
            .O(N__44619),
            .I(N__44616));
    Odrv4 I__7153 (
            .O(N__44616),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__7152 (
            .O(N__44613),
            .I(N__44610));
    LocalMux I__7151 (
            .O(N__44610),
            .I(N__44606));
    InMux I__7150 (
            .O(N__44609),
            .I(N__44603));
    Span4Mux_v I__7149 (
            .O(N__44606),
            .I(N__44600));
    LocalMux I__7148 (
            .O(N__44603),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    Odrv4 I__7147 (
            .O(N__44600),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    InMux I__7146 (
            .O(N__44595),
            .I(N__44592));
    LocalMux I__7145 (
            .O(N__44592),
            .I(N__44589));
    Span4Mux_h I__7144 (
            .O(N__44589),
            .I(N__44585));
    InMux I__7143 (
            .O(N__44588),
            .I(N__44582));
    Odrv4 I__7142 (
            .O(N__44585),
            .I(frame_decoder_CH4data_7));
    LocalMux I__7141 (
            .O(N__44582),
            .I(frame_decoder_CH4data_7));
    InMux I__7140 (
            .O(N__44577),
            .I(N__44574));
    LocalMux I__7139 (
            .O(N__44574),
            .I(\scaler_4.N_2232_i_l_ofxZ0 ));
    InMux I__7138 (
            .O(N__44571),
            .I(N__44568));
    LocalMux I__7137 (
            .O(N__44568),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__7136 (
            .O(N__44565),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__7135 (
            .O(N__44562),
            .I(bfn_11_9_0_));
    InMux I__7134 (
            .O(N__44559),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    CEMux I__7133 (
            .O(N__44556),
            .I(N__44553));
    LocalMux I__7132 (
            .O(N__44553),
            .I(N__44550));
    Span4Mux_v I__7131 (
            .O(N__44550),
            .I(N__44546));
    CEMux I__7130 (
            .O(N__44549),
            .I(N__44543));
    Span4Mux_v I__7129 (
            .O(N__44546),
            .I(N__44538));
    LocalMux I__7128 (
            .O(N__44543),
            .I(N__44538));
    Odrv4 I__7127 (
            .O(N__44538),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    InMux I__7126 (
            .O(N__44535),
            .I(N__44531));
    InMux I__7125 (
            .O(N__44534),
            .I(N__44528));
    LocalMux I__7124 (
            .O(N__44531),
            .I(N__44522));
    LocalMux I__7123 (
            .O(N__44528),
            .I(N__44522));
    InMux I__7122 (
            .O(N__44527),
            .I(N__44518));
    Span4Mux_h I__7121 (
            .O(N__44522),
            .I(N__44515));
    InMux I__7120 (
            .O(N__44521),
            .I(N__44512));
    LocalMux I__7119 (
            .O(N__44518),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__7118 (
            .O(N__44515),
            .I(frame_decoder_CH4data_0));
    LocalMux I__7117 (
            .O(N__44512),
            .I(frame_decoder_CH4data_0));
    InMux I__7116 (
            .O(N__44505),
            .I(N__44502));
    LocalMux I__7115 (
            .O(N__44502),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__7114 (
            .O(N__44499),
            .I(N__44495));
    InMux I__7113 (
            .O(N__44498),
            .I(N__44490));
    InMux I__7112 (
            .O(N__44495),
            .I(N__44485));
    InMux I__7111 (
            .O(N__44494),
            .I(N__44485));
    InMux I__7110 (
            .O(N__44493),
            .I(N__44482));
    LocalMux I__7109 (
            .O(N__44490),
            .I(N__44477));
    LocalMux I__7108 (
            .O(N__44485),
            .I(N__44477));
    LocalMux I__7107 (
            .O(N__44482),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__7106 (
            .O(N__44477),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__7105 (
            .O(N__44472),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__7104 (
            .O(N__44469),
            .I(N__44466));
    LocalMux I__7103 (
            .O(N__44466),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__7102 (
            .O(N__44463),
            .I(N__44460));
    InMux I__7101 (
            .O(N__44460),
            .I(N__44454));
    InMux I__7100 (
            .O(N__44459),
            .I(N__44454));
    LocalMux I__7099 (
            .O(N__44454),
            .I(N__44451));
    Odrv4 I__7098 (
            .O(N__44451),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__7097 (
            .O(N__44448),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__7096 (
            .O(N__44445),
            .I(N__44442));
    LocalMux I__7095 (
            .O(N__44442),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__7094 (
            .O(N__44439),
            .I(N__44436));
    InMux I__7093 (
            .O(N__44436),
            .I(N__44430));
    InMux I__7092 (
            .O(N__44435),
            .I(N__44430));
    LocalMux I__7091 (
            .O(N__44430),
            .I(N__44427));
    Odrv4 I__7090 (
            .O(N__44427),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__7089 (
            .O(N__44424),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__7088 (
            .O(N__44421),
            .I(N__44418));
    LocalMux I__7087 (
            .O(N__44418),
            .I(frame_decoder_CH4data_4));
    IoInMux I__7086 (
            .O(N__44415),
            .I(N__44412));
    LocalMux I__7085 (
            .O(N__44412),
            .I(N__44409));
    IoSpan4Mux I__7084 (
            .O(N__44409),
            .I(N__44405));
    CascadeMux I__7083 (
            .O(N__44408),
            .I(N__44400));
    IoSpan4Mux I__7082 (
            .O(N__44405),
            .I(N__44397));
    InMux I__7081 (
            .O(N__44404),
            .I(N__44392));
    InMux I__7080 (
            .O(N__44403),
            .I(N__44392));
    InMux I__7079 (
            .O(N__44400),
            .I(N__44389));
    Span4Mux_s3_v I__7078 (
            .O(N__44397),
            .I(N__44384));
    LocalMux I__7077 (
            .O(N__44392),
            .I(N__44384));
    LocalMux I__7076 (
            .O(N__44389),
            .I(debug_CH3_20A_c));
    Odrv4 I__7075 (
            .O(N__44384),
            .I(debug_CH3_20A_c));
    CascadeMux I__7074 (
            .O(N__44379),
            .I(N__44376));
    InMux I__7073 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__7072 (
            .O(N__44373),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__7071 (
            .O(N__44370),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    InMux I__7070 (
            .O(N__44367),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    InMux I__7069 (
            .O(N__44364),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    InMux I__7068 (
            .O(N__44361),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    InMux I__7067 (
            .O(N__44358),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    InMux I__7066 (
            .O(N__44355),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__7065 (
            .O(N__44352),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ));
    CascadeMux I__7064 (
            .O(N__44349),
            .I(\pid_front.error_i_reg_9_rn_0_16_cascade_ ));
    CascadeMux I__7063 (
            .O(N__44346),
            .I(N__44343));
    InMux I__7062 (
            .O(N__44343),
            .I(N__44340));
    LocalMux I__7061 (
            .O(N__44340),
            .I(N__44337));
    Odrv12 I__7060 (
            .O(N__44337),
            .I(\pid_front.error_i_regZ0Z_16 ));
    InMux I__7059 (
            .O(N__44334),
            .I(N__44331));
    LocalMux I__7058 (
            .O(N__44331),
            .I(\pid_front.m4_2_03 ));
    InMux I__7057 (
            .O(N__44328),
            .I(N__44325));
    LocalMux I__7056 (
            .O(N__44325),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ));
    CascadeMux I__7055 (
            .O(N__44322),
            .I(N__44319));
    InMux I__7054 (
            .O(N__44319),
            .I(N__44316));
    LocalMux I__7053 (
            .O(N__44316),
            .I(N__44313));
    Odrv12 I__7052 (
            .O(N__44313),
            .I(\pid_front.error_i_regZ0Z_2 ));
    CascadeMux I__7051 (
            .O(N__44310),
            .I(\pid_front.N_126_cascade_ ));
    InMux I__7050 (
            .O(N__44307),
            .I(N__44303));
    InMux I__7049 (
            .O(N__44306),
            .I(N__44300));
    LocalMux I__7048 (
            .O(N__44303),
            .I(\pid_front.N_12_1 ));
    LocalMux I__7047 (
            .O(N__44300),
            .I(\pid_front.N_12_1 ));
    CascadeMux I__7046 (
            .O(N__44295),
            .I(\pid_front.m1_0_03_cascade_ ));
    CascadeMux I__7045 (
            .O(N__44292),
            .I(\pid_front.N_93_0_cascade_ ));
    InMux I__7044 (
            .O(N__44289),
            .I(N__44286));
    LocalMux I__7043 (
            .O(N__44286),
            .I(\pid_front.m29_2_03_0 ));
    CascadeMux I__7042 (
            .O(N__44283),
            .I(\pid_front.error_i_reg_9_rn_0_25_cascade_ ));
    InMux I__7041 (
            .O(N__44280),
            .I(N__44277));
    LocalMux I__7040 (
            .O(N__44277),
            .I(N__44274));
    Odrv12 I__7039 (
            .O(N__44274),
            .I(\pid_front.error_i_regZ0Z_25 ));
    InMux I__7038 (
            .O(N__44271),
            .I(N__44268));
    LocalMux I__7037 (
            .O(N__44268),
            .I(\pid_front.N_93_0 ));
    CascadeMux I__7036 (
            .O(N__44265),
            .I(N__44262));
    InMux I__7035 (
            .O(N__44262),
            .I(N__44259));
    LocalMux I__7034 (
            .O(N__44259),
            .I(N__44256));
    Span4Mux_v I__7033 (
            .O(N__44256),
            .I(N__44253));
    Odrv4 I__7032 (
            .O(N__44253),
            .I(\pid_front.error_i_regZ0Z_9 ));
    CascadeMux I__7031 (
            .O(N__44250),
            .I(N__44246));
    InMux I__7030 (
            .O(N__44249),
            .I(N__44243));
    InMux I__7029 (
            .O(N__44246),
            .I(N__44240));
    LocalMux I__7028 (
            .O(N__44243),
            .I(N__44237));
    LocalMux I__7027 (
            .O(N__44240),
            .I(N__44234));
    Odrv4 I__7026 (
            .O(N__44237),
            .I(\pid_front.error_i_regZ0Z_0 ));
    Odrv12 I__7025 (
            .O(N__44234),
            .I(\pid_front.error_i_regZ0Z_0 ));
    CascadeMux I__7024 (
            .O(N__44229),
            .I(\pid_front.N_11_0_cascade_ ));
    CascadeMux I__7023 (
            .O(N__44226),
            .I(\pid_front.N_12_1_cascade_ ));
    CascadeMux I__7022 (
            .O(N__44223),
            .I(N__44220));
    InMux I__7021 (
            .O(N__44220),
            .I(N__44217));
    LocalMux I__7020 (
            .O(N__44217),
            .I(N__44214));
    Odrv12 I__7019 (
            .O(N__44214),
            .I(\pid_front.error_i_regZ0Z_1 ));
    InMux I__7018 (
            .O(N__44211),
            .I(N__44208));
    LocalMux I__7017 (
            .O(N__44208),
            .I(\pid_front.N_9_1 ));
    CascadeMux I__7016 (
            .O(N__44205),
            .I(\pid_front.N_9_1_cascade_ ));
    CascadeMux I__7015 (
            .O(N__44202),
            .I(\pid_front.N_39_0_cascade_ ));
    CascadeMux I__7014 (
            .O(N__44199),
            .I(\pid_front.m7_2_03_cascade_ ));
    CascadeMux I__7013 (
            .O(N__44196),
            .I(N__44193));
    InMux I__7012 (
            .O(N__44193),
            .I(N__44187));
    InMux I__7011 (
            .O(N__44192),
            .I(N__44187));
    LocalMux I__7010 (
            .O(N__44187),
            .I(N__44184));
    Odrv4 I__7009 (
            .O(N__44184),
            .I(\pid_front.error_i_acumm_preregZ0Z_27 ));
    CascadeMux I__7008 (
            .O(N__44181),
            .I(\pid_front.g0_8_1_cascade_ ));
    CascadeMux I__7007 (
            .O(N__44178),
            .I(\pid_front.N_88_0_0_cascade_ ));
    CascadeMux I__7006 (
            .O(N__44175),
            .I(\pid_front.g1_cascade_ ));
    InMux I__7005 (
            .O(N__44172),
            .I(N__44169));
    LocalMux I__7004 (
            .O(N__44169),
            .I(N__44166));
    Odrv4 I__7003 (
            .O(N__44166),
            .I(\pid_front.error_i_regZ0Z_21 ));
    InMux I__7002 (
            .O(N__44163),
            .I(N__44160));
    LocalMux I__7001 (
            .O(N__44160),
            .I(\pid_front.N_126_0 ));
    InMux I__7000 (
            .O(N__44157),
            .I(N__44154));
    LocalMux I__6999 (
            .O(N__44154),
            .I(\pid_front.g3 ));
    InMux I__6998 (
            .O(N__44151),
            .I(N__44145));
    InMux I__6997 (
            .O(N__44150),
            .I(N__44145));
    LocalMux I__6996 (
            .O(N__44145),
            .I(\pid_front.error_i_regZ0Z_27 ));
    InMux I__6995 (
            .O(N__44142),
            .I(N__44139));
    LocalMux I__6994 (
            .O(N__44139),
            .I(N__44136));
    Span4Mux_h I__6993 (
            .O(N__44136),
            .I(N__44133));
    Odrv4 I__6992 (
            .O(N__44133),
            .I(\pid_front.error_i_regZ0Z_23 ));
    InMux I__6991 (
            .O(N__44130),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__6990 (
            .O(N__44127),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__6989 (
            .O(N__44124),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_22 ));
    InMux I__6988 (
            .O(N__44121),
            .I(N__44116));
    InMux I__6987 (
            .O(N__44120),
            .I(N__44111));
    InMux I__6986 (
            .O(N__44119),
            .I(N__44111));
    LocalMux I__6985 (
            .O(N__44116),
            .I(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ));
    LocalMux I__6984 (
            .O(N__44111),
            .I(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ));
    InMux I__6983 (
            .O(N__44106),
            .I(bfn_10_21_0_));
    InMux I__6982 (
            .O(N__44103),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_24 ));
    InMux I__6981 (
            .O(N__44100),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_25 ));
    InMux I__6980 (
            .O(N__44097),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26 ));
    CascadeMux I__6979 (
            .O(N__44094),
            .I(N__44089));
    CascadeMux I__6978 (
            .O(N__44093),
            .I(N__44085));
    InMux I__6977 (
            .O(N__44092),
            .I(N__44068));
    InMux I__6976 (
            .O(N__44089),
            .I(N__44068));
    InMux I__6975 (
            .O(N__44088),
            .I(N__44068));
    InMux I__6974 (
            .O(N__44085),
            .I(N__44068));
    InMux I__6973 (
            .O(N__44084),
            .I(N__44068));
    CascadeMux I__6972 (
            .O(N__44083),
            .I(N__44065));
    CascadeMux I__6971 (
            .O(N__44082),
            .I(N__44061));
    CascadeMux I__6970 (
            .O(N__44081),
            .I(N__44057));
    CascadeMux I__6969 (
            .O(N__44080),
            .I(N__44053));
    CascadeMux I__6968 (
            .O(N__44079),
            .I(N__44048));
    LocalMux I__6967 (
            .O(N__44068),
            .I(N__44044));
    InMux I__6966 (
            .O(N__44065),
            .I(N__44027));
    InMux I__6965 (
            .O(N__44064),
            .I(N__44027));
    InMux I__6964 (
            .O(N__44061),
            .I(N__44027));
    InMux I__6963 (
            .O(N__44060),
            .I(N__44027));
    InMux I__6962 (
            .O(N__44057),
            .I(N__44027));
    InMux I__6961 (
            .O(N__44056),
            .I(N__44027));
    InMux I__6960 (
            .O(N__44053),
            .I(N__44027));
    InMux I__6959 (
            .O(N__44052),
            .I(N__44027));
    InMux I__6958 (
            .O(N__44051),
            .I(N__44020));
    InMux I__6957 (
            .O(N__44048),
            .I(N__44020));
    InMux I__6956 (
            .O(N__44047),
            .I(N__44020));
    Odrv4 I__6955 (
            .O(N__44044),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    LocalMux I__6954 (
            .O(N__44027),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    LocalMux I__6953 (
            .O(N__44020),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    InMux I__6952 (
            .O(N__44013),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__6951 (
            .O(N__44010),
            .I(N__44005));
    InMux I__6950 (
            .O(N__44009),
            .I(N__44000));
    InMux I__6949 (
            .O(N__44008),
            .I(N__44000));
    LocalMux I__6948 (
            .O(N__44005),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    LocalMux I__6947 (
            .O(N__44000),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    CascadeMux I__6946 (
            .O(N__43995),
            .I(N__43990));
    InMux I__6945 (
            .O(N__43994),
            .I(N__43987));
    InMux I__6944 (
            .O(N__43993),
            .I(N__43982));
    InMux I__6943 (
            .O(N__43990),
            .I(N__43982));
    LocalMux I__6942 (
            .O(N__43987),
            .I(N__43977));
    LocalMux I__6941 (
            .O(N__43982),
            .I(N__43977));
    Odrv4 I__6940 (
            .O(N__43977),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    InMux I__6939 (
            .O(N__43974),
            .I(N__43971));
    LocalMux I__6938 (
            .O(N__43971),
            .I(\pid_front.error_i_acummZ0Z_12 ));
    InMux I__6937 (
            .O(N__43968),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__6936 (
            .O(N__43965),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__6935 (
            .O(N__43962),
            .I(N__43957));
    InMux I__6934 (
            .O(N__43961),
            .I(N__43952));
    InMux I__6933 (
            .O(N__43960),
            .I(N__43952));
    LocalMux I__6932 (
            .O(N__43957),
            .I(N__43949));
    LocalMux I__6931 (
            .O(N__43952),
            .I(N__43946));
    Span4Mux_v I__6930 (
            .O(N__43949),
            .I(N__43943));
    Span4Mux_h I__6929 (
            .O(N__43946),
            .I(N__43940));
    Odrv4 I__6928 (
            .O(N__43943),
            .I(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ));
    Odrv4 I__6927 (
            .O(N__43940),
            .I(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ));
    InMux I__6926 (
            .O(N__43935),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__6925 (
            .O(N__43932),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__6924 (
            .O(N__43929),
            .I(bfn_10_20_0_));
    InMux I__6923 (
            .O(N__43926),
            .I(N__43921));
    InMux I__6922 (
            .O(N__43925),
            .I(N__43916));
    InMux I__6921 (
            .O(N__43924),
            .I(N__43916));
    LocalMux I__6920 (
            .O(N__43921),
            .I(N__43913));
    LocalMux I__6919 (
            .O(N__43916),
            .I(N__43910));
    Odrv4 I__6918 (
            .O(N__43913),
            .I(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ));
    Odrv4 I__6917 (
            .O(N__43910),
            .I(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ));
    InMux I__6916 (
            .O(N__43905),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__6915 (
            .O(N__43902),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__6914 (
            .O(N__43899),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__6913 (
            .O(N__43896),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__6912 (
            .O(N__43893),
            .I(N__43890));
    LocalMux I__6911 (
            .O(N__43890),
            .I(\pid_front.error_i_acummZ0Z_4 ));
    InMux I__6910 (
            .O(N__43887),
            .I(N__43884));
    LocalMux I__6909 (
            .O(N__43884),
            .I(N__43879));
    InMux I__6908 (
            .O(N__43883),
            .I(N__43874));
    InMux I__6907 (
            .O(N__43882),
            .I(N__43874));
    Span4Mux_v I__6906 (
            .O(N__43879),
            .I(N__43869));
    LocalMux I__6905 (
            .O(N__43874),
            .I(N__43869));
    Odrv4 I__6904 (
            .O(N__43869),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ));
    InMux I__6903 (
            .O(N__43866),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__6902 (
            .O(N__43863),
            .I(N__43860));
    LocalMux I__6901 (
            .O(N__43860),
            .I(\pid_front.error_i_acummZ0Z_5 ));
    InMux I__6900 (
            .O(N__43857),
            .I(N__43852));
    InMux I__6899 (
            .O(N__43856),
            .I(N__43849));
    InMux I__6898 (
            .O(N__43855),
            .I(N__43845));
    LocalMux I__6897 (
            .O(N__43852),
            .I(N__43840));
    LocalMux I__6896 (
            .O(N__43849),
            .I(N__43840));
    InMux I__6895 (
            .O(N__43848),
            .I(N__43837));
    LocalMux I__6894 (
            .O(N__43845),
            .I(N__43834));
    Span4Mux_v I__6893 (
            .O(N__43840),
            .I(N__43829));
    LocalMux I__6892 (
            .O(N__43837),
            .I(N__43829));
    Odrv12 I__6891 (
            .O(N__43834),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNILQKE ));
    Odrv4 I__6890 (
            .O(N__43829),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNILQKE ));
    InMux I__6889 (
            .O(N__43824),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__6888 (
            .O(N__43821),
            .I(N__43818));
    LocalMux I__6887 (
            .O(N__43818),
            .I(\pid_front.error_i_acummZ0Z_6 ));
    InMux I__6886 (
            .O(N__43815),
            .I(N__43812));
    LocalMux I__6885 (
            .O(N__43812),
            .I(N__43807));
    InMux I__6884 (
            .O(N__43811),
            .I(N__43802));
    InMux I__6883 (
            .O(N__43810),
            .I(N__43802));
    Span4Mux_v I__6882 (
            .O(N__43807),
            .I(N__43797));
    LocalMux I__6881 (
            .O(N__43802),
            .I(N__43797));
    Odrv4 I__6880 (
            .O(N__43797),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ));
    InMux I__6879 (
            .O(N__43794),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5 ));
    CascadeMux I__6878 (
            .O(N__43791),
            .I(N__43788));
    InMux I__6877 (
            .O(N__43788),
            .I(N__43785));
    LocalMux I__6876 (
            .O(N__43785),
            .I(\pid_front.error_i_acummZ0Z_7 ));
    InMux I__6875 (
            .O(N__43782),
            .I(N__43777));
    InMux I__6874 (
            .O(N__43781),
            .I(N__43772));
    InMux I__6873 (
            .O(N__43780),
            .I(N__43772));
    LocalMux I__6872 (
            .O(N__43777),
            .I(N__43769));
    LocalMux I__6871 (
            .O(N__43772),
            .I(N__43766));
    Span4Mux_h I__6870 (
            .O(N__43769),
            .I(N__43763));
    Span4Mux_h I__6869 (
            .O(N__43766),
            .I(N__43760));
    Odrv4 I__6868 (
            .O(N__43763),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ));
    Odrv4 I__6867 (
            .O(N__43760),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ));
    InMux I__6866 (
            .O(N__43755),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__6865 (
            .O(N__43752),
            .I(N__43749));
    LocalMux I__6864 (
            .O(N__43749),
            .I(\pid_front.error_i_acummZ0Z_8 ));
    InMux I__6863 (
            .O(N__43746),
            .I(N__43741));
    InMux I__6862 (
            .O(N__43745),
            .I(N__43736));
    InMux I__6861 (
            .O(N__43744),
            .I(N__43736));
    LocalMux I__6860 (
            .O(N__43741),
            .I(N__43733));
    LocalMux I__6859 (
            .O(N__43736),
            .I(N__43730));
    Span4Mux_h I__6858 (
            .O(N__43733),
            .I(N__43727));
    Span4Mux_v I__6857 (
            .O(N__43730),
            .I(N__43724));
    Odrv4 I__6856 (
            .O(N__43727),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    Odrv4 I__6855 (
            .O(N__43724),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    InMux I__6854 (
            .O(N__43719),
            .I(bfn_10_19_0_));
    InMux I__6853 (
            .O(N__43716),
            .I(N__43713));
    LocalMux I__6852 (
            .O(N__43713),
            .I(\pid_front.error_i_acummZ0Z_9 ));
    InMux I__6851 (
            .O(N__43710),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__6850 (
            .O(N__43707),
            .I(N__43704));
    LocalMux I__6849 (
            .O(N__43704),
            .I(\pid_front.error_i_acummZ0Z_10 ));
    InMux I__6848 (
            .O(N__43701),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__6847 (
            .O(N__43698),
            .I(N__43695));
    LocalMux I__6846 (
            .O(N__43695),
            .I(\pid_front.error_i_acummZ0Z_11 ));
    InMux I__6845 (
            .O(N__43692),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__6844 (
            .O(N__43689),
            .I(N__43685));
    InMux I__6843 (
            .O(N__43688),
            .I(N__43682));
    LocalMux I__6842 (
            .O(N__43685),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    LocalMux I__6841 (
            .O(N__43682),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    CascadeMux I__6840 (
            .O(N__43677),
            .I(\pid_front.un1_pid_prereg_0_4_cascade_ ));
    CascadeMux I__6839 (
            .O(N__43674),
            .I(\pid_front.un1_pid_prereg_0_5_cascade_ ));
    InMux I__6838 (
            .O(N__43671),
            .I(N__43666));
    InMux I__6837 (
            .O(N__43670),
            .I(N__43661));
    InMux I__6836 (
            .O(N__43669),
            .I(N__43661));
    LocalMux I__6835 (
            .O(N__43666),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    LocalMux I__6834 (
            .O(N__43661),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    InMux I__6833 (
            .O(N__43656),
            .I(N__43653));
    LocalMux I__6832 (
            .O(N__43653),
            .I(N__43649));
    InMux I__6831 (
            .O(N__43652),
            .I(N__43646));
    Odrv12 I__6830 (
            .O(N__43649),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    LocalMux I__6829 (
            .O(N__43646),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    InMux I__6828 (
            .O(N__43641),
            .I(N__43638));
    LocalMux I__6827 (
            .O(N__43638),
            .I(\pid_front.error_i_acummZ0Z_1 ));
    InMux I__6826 (
            .O(N__43635),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__6825 (
            .O(N__43632),
            .I(N__43629));
    LocalMux I__6824 (
            .O(N__43629),
            .I(\pid_front.error_i_acummZ0Z_2 ));
    InMux I__6823 (
            .O(N__43626),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__6822 (
            .O(N__43623),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2 ));
    CascadeMux I__6821 (
            .O(N__43620),
            .I(N__43615));
    InMux I__6820 (
            .O(N__43619),
            .I(N__43612));
    InMux I__6819 (
            .O(N__43618),
            .I(N__43609));
    InMux I__6818 (
            .O(N__43615),
            .I(N__43606));
    LocalMux I__6817 (
            .O(N__43612),
            .I(N__43603));
    LocalMux I__6816 (
            .O(N__43609),
            .I(\pid_front.un1_pid_prereg_79 ));
    LocalMux I__6815 (
            .O(N__43606),
            .I(\pid_front.un1_pid_prereg_79 ));
    Odrv4 I__6814 (
            .O(N__43603),
            .I(\pid_front.un1_pid_prereg_79 ));
    InMux I__6813 (
            .O(N__43596),
            .I(N__43590));
    InMux I__6812 (
            .O(N__43595),
            .I(N__43587));
    InMux I__6811 (
            .O(N__43594),
            .I(N__43584));
    InMux I__6810 (
            .O(N__43593),
            .I(N__43581));
    LocalMux I__6809 (
            .O(N__43590),
            .I(N__43578));
    LocalMux I__6808 (
            .O(N__43587),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    LocalMux I__6807 (
            .O(N__43584),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    LocalMux I__6806 (
            .O(N__43581),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    Odrv4 I__6805 (
            .O(N__43578),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    CascadeMux I__6804 (
            .O(N__43569),
            .I(\pid_front.error_p_reg_esr_RNIJ1FT1Z0Z_12_cascade_ ));
    InMux I__6803 (
            .O(N__43566),
            .I(N__43563));
    LocalMux I__6802 (
            .O(N__43563),
            .I(\pid_front.un1_pid_prereg_167_0_1 ));
    InMux I__6801 (
            .O(N__43560),
            .I(N__43556));
    InMux I__6800 (
            .O(N__43559),
            .I(N__43550));
    LocalMux I__6799 (
            .O(N__43556),
            .I(N__43547));
    InMux I__6798 (
            .O(N__43555),
            .I(N__43544));
    InMux I__6797 (
            .O(N__43554),
            .I(N__43539));
    InMux I__6796 (
            .O(N__43553),
            .I(N__43539));
    LocalMux I__6795 (
            .O(N__43550),
            .I(\pid_front.error_p_regZ0Z_12 ));
    Odrv4 I__6794 (
            .O(N__43547),
            .I(\pid_front.error_p_regZ0Z_12 ));
    LocalMux I__6793 (
            .O(N__43544),
            .I(\pid_front.error_p_regZ0Z_12 ));
    LocalMux I__6792 (
            .O(N__43539),
            .I(\pid_front.error_p_regZ0Z_12 ));
    InMux I__6791 (
            .O(N__43530),
            .I(N__43527));
    LocalMux I__6790 (
            .O(N__43527),
            .I(\pid_front.error_p_reg_esr_RNIBQB61Z0Z_12 ));
    InMux I__6789 (
            .O(N__43524),
            .I(N__43518));
    InMux I__6788 (
            .O(N__43523),
            .I(N__43518));
    LocalMux I__6787 (
            .O(N__43518),
            .I(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12 ));
    CascadeMux I__6786 (
            .O(N__43515),
            .I(N__43512));
    InMux I__6785 (
            .O(N__43512),
            .I(N__43509));
    LocalMux I__6784 (
            .O(N__43509),
            .I(\pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12 ));
    CascadeMux I__6783 (
            .O(N__43506),
            .I(\pid_front.un1_pid_prereg_0_3_cascade_ ));
    CascadeMux I__6782 (
            .O(N__43503),
            .I(N__43499));
    InMux I__6781 (
            .O(N__43502),
            .I(N__43496));
    InMux I__6780 (
            .O(N__43499),
            .I(N__43493));
    LocalMux I__6779 (
            .O(N__43496),
            .I(\pid_front.N_1698_i ));
    LocalMux I__6778 (
            .O(N__43493),
            .I(\pid_front.N_1698_i ));
    InMux I__6777 (
            .O(N__43488),
            .I(N__43485));
    LocalMux I__6776 (
            .O(N__43485),
            .I(N__43482));
    Span4Mux_h I__6775 (
            .O(N__43482),
            .I(N__43479));
    Span4Mux_h I__6774 (
            .O(N__43479),
            .I(N__43476));
    Span4Mux_h I__6773 (
            .O(N__43476),
            .I(N__43473));
    Odrv4 I__6772 (
            .O(N__43473),
            .I(\pid_front.O_0_15 ));
    InMux I__6771 (
            .O(N__43470),
            .I(N__43467));
    LocalMux I__6770 (
            .O(N__43467),
            .I(\pid_front.pid_prereg_esr_RNIBQKJ3Z0Z_20 ));
    InMux I__6769 (
            .O(N__43464),
            .I(N__43460));
    InMux I__6768 (
            .O(N__43463),
            .I(N__43457));
    LocalMux I__6767 (
            .O(N__43460),
            .I(N__43454));
    LocalMux I__6766 (
            .O(N__43457),
            .I(\pid_front.un11lto30_i_a2_4_and ));
    Odrv4 I__6765 (
            .O(N__43454),
            .I(\pid_front.un11lto30_i_a2_4_and ));
    InMux I__6764 (
            .O(N__43449),
            .I(N__43442));
    InMux I__6763 (
            .O(N__43448),
            .I(N__43442));
    InMux I__6762 (
            .O(N__43447),
            .I(N__43439));
    LocalMux I__6761 (
            .O(N__43442),
            .I(\pid_front.un11lto30_i_a2_6_and ));
    LocalMux I__6760 (
            .O(N__43439),
            .I(\pid_front.un11lto30_i_a2_6_and ));
    InMux I__6759 (
            .O(N__43434),
            .I(N__43427));
    InMux I__6758 (
            .O(N__43433),
            .I(N__43427));
    InMux I__6757 (
            .O(N__43432),
            .I(N__43424));
    LocalMux I__6756 (
            .O(N__43427),
            .I(\pid_front.un11lto30_i_a2_5_and ));
    LocalMux I__6755 (
            .O(N__43424),
            .I(\pid_front.un11lto30_i_a2_5_and ));
    CascadeMux I__6754 (
            .O(N__43419),
            .I(\pid_front.un11lto30_i_a2_4_and_cascade_ ));
    InMux I__6753 (
            .O(N__43416),
            .I(N__43413));
    LocalMux I__6752 (
            .O(N__43413),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ));
    CascadeMux I__6751 (
            .O(N__43410),
            .I(\pid_front.N_98_cascade_ ));
    CascadeMux I__6750 (
            .O(N__43407),
            .I(\pid_front.N_389_cascade_ ));
    CascadeMux I__6749 (
            .O(N__43404),
            .I(\pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12_cascade_ ));
    InMux I__6748 (
            .O(N__43401),
            .I(N__43398));
    LocalMux I__6747 (
            .O(N__43398),
            .I(N__43395));
    Odrv4 I__6746 (
            .O(N__43395),
            .I(\pid_front.un11lto30_i_a2_2_and ));
    InMux I__6745 (
            .O(N__43392),
            .I(N__43389));
    LocalMux I__6744 (
            .O(N__43389),
            .I(N__43386));
    Odrv4 I__6743 (
            .O(N__43386),
            .I(\pid_front.un11lto30_i_a2_3_and ));
    InMux I__6742 (
            .O(N__43383),
            .I(bfn_10_14_0_));
    InMux I__6741 (
            .O(N__43380),
            .I(N__43377));
    LocalMux I__6740 (
            .O(N__43377),
            .I(\pid_front.un11lto30_i_a2_0_and ));
    CascadeMux I__6739 (
            .O(N__43374),
            .I(N__43370));
    InMux I__6738 (
            .O(N__43373),
            .I(N__43367));
    InMux I__6737 (
            .O(N__43370),
            .I(N__43364));
    LocalMux I__6736 (
            .O(N__43367),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__6735 (
            .O(N__43364),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    CascadeMux I__6734 (
            .O(N__43359),
            .I(N__43355));
    InMux I__6733 (
            .O(N__43358),
            .I(N__43352));
    InMux I__6732 (
            .O(N__43355),
            .I(N__43349));
    LocalMux I__6731 (
            .O(N__43352),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__6730 (
            .O(N__43349),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__6729 (
            .O(N__43344),
            .I(N__43340));
    InMux I__6728 (
            .O(N__43343),
            .I(N__43337));
    LocalMux I__6727 (
            .O(N__43340),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__6726 (
            .O(N__43337),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    CascadeMux I__6725 (
            .O(N__43332),
            .I(N__43328));
    InMux I__6724 (
            .O(N__43331),
            .I(N__43325));
    InMux I__6723 (
            .O(N__43328),
            .I(N__43322));
    LocalMux I__6722 (
            .O(N__43325),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__6721 (
            .O(N__43322),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__6720 (
            .O(N__43317),
            .I(N__43313));
    InMux I__6719 (
            .O(N__43316),
            .I(N__43310));
    InMux I__6718 (
            .O(N__43313),
            .I(N__43307));
    LocalMux I__6717 (
            .O(N__43310),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__6716 (
            .O(N__43307),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__6715 (
            .O(N__43302),
            .I(N__43298));
    InMux I__6714 (
            .O(N__43301),
            .I(N__43295));
    InMux I__6713 (
            .O(N__43298),
            .I(N__43292));
    LocalMux I__6712 (
            .O(N__43295),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__6711 (
            .O(N__43292),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CEMux I__6710 (
            .O(N__43287),
            .I(N__43284));
    LocalMux I__6709 (
            .O(N__43284),
            .I(N__43281));
    Span4Mux_v I__6708 (
            .O(N__43281),
            .I(N__43278));
    Odrv4 I__6707 (
            .O(N__43278),
            .I(\uart_drone.data_rdyc_1_0 ));
    SRMux I__6706 (
            .O(N__43275),
            .I(N__43272));
    LocalMux I__6705 (
            .O(N__43272),
            .I(N__43269));
    Span4Mux_v I__6704 (
            .O(N__43269),
            .I(N__43266));
    Span4Mux_h I__6703 (
            .O(N__43266),
            .I(N__43263));
    Odrv4 I__6702 (
            .O(N__43263),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    InMux I__6701 (
            .O(N__43260),
            .I(N__43257));
    LocalMux I__6700 (
            .O(N__43257),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__6699 (
            .O(N__43254),
            .I(N__43251));
    LocalMux I__6698 (
            .O(N__43251),
            .I(\uart_drone.data_Auxce_0_3 ));
    InMux I__6697 (
            .O(N__43248),
            .I(N__43245));
    LocalMux I__6696 (
            .O(N__43245),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__6695 (
            .O(N__43242),
            .I(N__43239));
    LocalMux I__6694 (
            .O(N__43239),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__6693 (
            .O(N__43236),
            .I(N__43212));
    InMux I__6692 (
            .O(N__43235),
            .I(N__43212));
    InMux I__6691 (
            .O(N__43234),
            .I(N__43212));
    InMux I__6690 (
            .O(N__43233),
            .I(N__43212));
    InMux I__6689 (
            .O(N__43232),
            .I(N__43212));
    InMux I__6688 (
            .O(N__43231),
            .I(N__43212));
    InMux I__6687 (
            .O(N__43230),
            .I(N__43212));
    InMux I__6686 (
            .O(N__43229),
            .I(N__43212));
    LocalMux I__6685 (
            .O(N__43212),
            .I(N__43209));
    Odrv12 I__6684 (
            .O(N__43209),
            .I(\uart_drone.un1_state_2_0 ));
    InMux I__6683 (
            .O(N__43206),
            .I(N__43203));
    LocalMux I__6682 (
            .O(N__43203),
            .I(N__43198));
    InMux I__6681 (
            .O(N__43202),
            .I(N__43193));
    InMux I__6680 (
            .O(N__43201),
            .I(N__43193));
    Odrv4 I__6679 (
            .O(N__43198),
            .I(\uart_drone.N_152 ));
    LocalMux I__6678 (
            .O(N__43193),
            .I(\uart_drone.N_152 ));
    IoInMux I__6677 (
            .O(N__43188),
            .I(N__43185));
    LocalMux I__6676 (
            .O(N__43185),
            .I(N__43180));
    CascadeMux I__6675 (
            .O(N__43184),
            .I(N__43170));
    CascadeMux I__6674 (
            .O(N__43183),
            .I(N__43167));
    Span4Mux_s1_v I__6673 (
            .O(N__43180),
            .I(N__43164));
    InMux I__6672 (
            .O(N__43179),
            .I(N__43161));
    InMux I__6671 (
            .O(N__43178),
            .I(N__43156));
    InMux I__6670 (
            .O(N__43177),
            .I(N__43156));
    InMux I__6669 (
            .O(N__43176),
            .I(N__43143));
    InMux I__6668 (
            .O(N__43175),
            .I(N__43143));
    InMux I__6667 (
            .O(N__43174),
            .I(N__43143));
    InMux I__6666 (
            .O(N__43173),
            .I(N__43143));
    InMux I__6665 (
            .O(N__43170),
            .I(N__43143));
    InMux I__6664 (
            .O(N__43167),
            .I(N__43143));
    Sp12to4 I__6663 (
            .O(N__43164),
            .I(N__43138));
    LocalMux I__6662 (
            .O(N__43161),
            .I(N__43135));
    LocalMux I__6661 (
            .O(N__43156),
            .I(N__43128));
    LocalMux I__6660 (
            .O(N__43143),
            .I(N__43128));
    InMux I__6659 (
            .O(N__43142),
            .I(N__43123));
    InMux I__6658 (
            .O(N__43141),
            .I(N__43123));
    Span12Mux_h I__6657 (
            .O(N__43138),
            .I(N__43118));
    Span12Mux_s10_h I__6656 (
            .O(N__43135),
            .I(N__43118));
    InMux I__6655 (
            .O(N__43134),
            .I(N__43113));
    InMux I__6654 (
            .O(N__43133),
            .I(N__43113));
    Odrv4 I__6653 (
            .O(N__43128),
            .I(debug_CH0_16A_c));
    LocalMux I__6652 (
            .O(N__43123),
            .I(debug_CH0_16A_c));
    Odrv12 I__6651 (
            .O(N__43118),
            .I(debug_CH0_16A_c));
    LocalMux I__6650 (
            .O(N__43113),
            .I(debug_CH0_16A_c));
    SRMux I__6649 (
            .O(N__43104),
            .I(N__43101));
    LocalMux I__6648 (
            .O(N__43101),
            .I(N__43098));
    Span4Mux_h I__6647 (
            .O(N__43098),
            .I(N__43095));
    Odrv4 I__6646 (
            .O(N__43095),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__6645 (
            .O(N__43092),
            .I(N__43088));
    InMux I__6644 (
            .O(N__43091),
            .I(N__43085));
    LocalMux I__6643 (
            .O(N__43088),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__6642 (
            .O(N__43085),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    CascadeMux I__6641 (
            .O(N__43080),
            .I(N__43076));
    InMux I__6640 (
            .O(N__43079),
            .I(N__43073));
    InMux I__6639 (
            .O(N__43076),
            .I(N__43070));
    LocalMux I__6638 (
            .O(N__43073),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__6637 (
            .O(N__43070),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__6636 (
            .O(N__43065),
            .I(N__43058));
    CascadeMux I__6635 (
            .O(N__43064),
            .I(N__43055));
    CascadeMux I__6634 (
            .O(N__43063),
            .I(N__43051));
    InMux I__6633 (
            .O(N__43062),
            .I(N__43042));
    InMux I__6632 (
            .O(N__43061),
            .I(N__43042));
    InMux I__6631 (
            .O(N__43058),
            .I(N__43042));
    InMux I__6630 (
            .O(N__43055),
            .I(N__43039));
    InMux I__6629 (
            .O(N__43054),
            .I(N__43036));
    InMux I__6628 (
            .O(N__43051),
            .I(N__43031));
    InMux I__6627 (
            .O(N__43050),
            .I(N__43031));
    InMux I__6626 (
            .O(N__43049),
            .I(N__43028));
    LocalMux I__6625 (
            .O(N__43042),
            .I(N__43025));
    LocalMux I__6624 (
            .O(N__43039),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__6623 (
            .O(N__43036),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__6622 (
            .O(N__43031),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__6621 (
            .O(N__43028),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__6620 (
            .O(N__43025),
            .I(\uart_drone.stateZ0Z_3 ));
    CascadeMux I__6619 (
            .O(N__43014),
            .I(N__43010));
    InMux I__6618 (
            .O(N__43013),
            .I(N__43002));
    InMux I__6617 (
            .O(N__43010),
            .I(N__43002));
    InMux I__6616 (
            .O(N__43009),
            .I(N__43002));
    LocalMux I__6615 (
            .O(N__43002),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__6614 (
            .O(N__42999),
            .I(N__42990));
    InMux I__6613 (
            .O(N__42998),
            .I(N__42990));
    InMux I__6612 (
            .O(N__42997),
            .I(N__42984));
    InMux I__6611 (
            .O(N__42996),
            .I(N__42981));
    InMux I__6610 (
            .O(N__42995),
            .I(N__42978));
    LocalMux I__6609 (
            .O(N__42990),
            .I(N__42975));
    InMux I__6608 (
            .O(N__42989),
            .I(N__42968));
    InMux I__6607 (
            .O(N__42988),
            .I(N__42968));
    InMux I__6606 (
            .O(N__42987),
            .I(N__42968));
    LocalMux I__6605 (
            .O(N__42984),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__6604 (
            .O(N__42981),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__6603 (
            .O(N__42978),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__6602 (
            .O(N__42975),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__6601 (
            .O(N__42968),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__6600 (
            .O(N__42957),
            .I(N__42952));
    InMux I__6599 (
            .O(N__42956),
            .I(N__42944));
    InMux I__6598 (
            .O(N__42955),
            .I(N__42944));
    LocalMux I__6597 (
            .O(N__42952),
            .I(N__42941));
    InMux I__6596 (
            .O(N__42951),
            .I(N__42938));
    InMux I__6595 (
            .O(N__42950),
            .I(N__42933));
    InMux I__6594 (
            .O(N__42949),
            .I(N__42933));
    LocalMux I__6593 (
            .O(N__42944),
            .I(N__42927));
    Span4Mux_v I__6592 (
            .O(N__42941),
            .I(N__42920));
    LocalMux I__6591 (
            .O(N__42938),
            .I(N__42920));
    LocalMux I__6590 (
            .O(N__42933),
            .I(N__42920));
    InMux I__6589 (
            .O(N__42932),
            .I(N__42913));
    InMux I__6588 (
            .O(N__42931),
            .I(N__42913));
    InMux I__6587 (
            .O(N__42930),
            .I(N__42913));
    Span4Mux_h I__6586 (
            .O(N__42927),
            .I(N__42910));
    Odrv4 I__6585 (
            .O(N__42920),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__6584 (
            .O(N__42913),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__6583 (
            .O(N__42910),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__6582 (
            .O(N__42903),
            .I(N__42897));
    InMux I__6581 (
            .O(N__42902),
            .I(N__42897));
    LocalMux I__6580 (
            .O(N__42897),
            .I(N__42894));
    Odrv4 I__6579 (
            .O(N__42894),
            .I(\uart_drone.N_144_1 ));
    CEMux I__6578 (
            .O(N__42891),
            .I(N__42888));
    LocalMux I__6577 (
            .O(N__42888),
            .I(N__42884));
    CEMux I__6576 (
            .O(N__42887),
            .I(N__42881));
    Span4Mux_v I__6575 (
            .O(N__42884),
            .I(N__42878));
    LocalMux I__6574 (
            .O(N__42881),
            .I(N__42875));
    Span4Mux_v I__6573 (
            .O(N__42878),
            .I(N__42870));
    Span4Mux_h I__6572 (
            .O(N__42875),
            .I(N__42870));
    Span4Mux_h I__6571 (
            .O(N__42870),
            .I(N__42867));
    Odrv4 I__6570 (
            .O(N__42867),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__6569 (
            .O(N__42864),
            .I(N__42861));
    LocalMux I__6568 (
            .O(N__42861),
            .I(N__42858));
    Odrv4 I__6567 (
            .O(N__42858),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__6566 (
            .O(N__42855),
            .I(N__42852));
    LocalMux I__6565 (
            .O(N__42852),
            .I(N__42849));
    Odrv12 I__6564 (
            .O(N__42849),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__6563 (
            .O(N__42846),
            .I(N__42843));
    LocalMux I__6562 (
            .O(N__42843),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    CascadeMux I__6561 (
            .O(N__42840),
            .I(\uart_drone.N_152_cascade_ ));
    CascadeMux I__6560 (
            .O(N__42837),
            .I(\uart_drone.un1_state_7_0_cascade_ ));
    InMux I__6559 (
            .O(N__42834),
            .I(N__42827));
    InMux I__6558 (
            .O(N__42833),
            .I(N__42823));
    InMux I__6557 (
            .O(N__42832),
            .I(N__42820));
    InMux I__6556 (
            .O(N__42831),
            .I(N__42817));
    InMux I__6555 (
            .O(N__42830),
            .I(N__42814));
    LocalMux I__6554 (
            .O(N__42827),
            .I(N__42811));
    InMux I__6553 (
            .O(N__42826),
            .I(N__42808));
    LocalMux I__6552 (
            .O(N__42823),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6551 (
            .O(N__42820),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6550 (
            .O(N__42817),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6549 (
            .O(N__42814),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__6548 (
            .O(N__42811),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6547 (
            .O(N__42808),
            .I(\uart_drone.stateZ0Z_4 ));
    CascadeMux I__6546 (
            .O(N__42795),
            .I(\uart_drone.un1_state_4_0_cascade_ ));
    InMux I__6545 (
            .O(N__42792),
            .I(N__42789));
    LocalMux I__6544 (
            .O(N__42789),
            .I(\uart_drone.un1_state_7_0 ));
    CascadeMux I__6543 (
            .O(N__42786),
            .I(\uart_drone.CO0_cascade_ ));
    CascadeMux I__6542 (
            .O(N__42783),
            .I(N__42780));
    InMux I__6541 (
            .O(N__42780),
            .I(N__42777));
    LocalMux I__6540 (
            .O(N__42777),
            .I(N__42774));
    Odrv4 I__6539 (
            .O(N__42774),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    CascadeMux I__6538 (
            .O(N__42771),
            .I(N__42766));
    InMux I__6537 (
            .O(N__42770),
            .I(N__42759));
    InMux I__6536 (
            .O(N__42769),
            .I(N__42759));
    InMux I__6535 (
            .O(N__42766),
            .I(N__42759));
    LocalMux I__6534 (
            .O(N__42759),
            .I(\uart_drone.stateZ0Z_1 ));
    CascadeMux I__6533 (
            .O(N__42756),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__6532 (
            .O(N__42753),
            .I(N__42750));
    LocalMux I__6531 (
            .O(N__42750),
            .I(\uart_drone.N_145 ));
    CascadeMux I__6530 (
            .O(N__42747),
            .I(N__42743));
    CascadeMux I__6529 (
            .O(N__42746),
            .I(N__42739));
    InMux I__6528 (
            .O(N__42743),
            .I(N__42732));
    InMux I__6527 (
            .O(N__42742),
            .I(N__42732));
    InMux I__6526 (
            .O(N__42739),
            .I(N__42732));
    LocalMux I__6525 (
            .O(N__42732),
            .I(N__42728));
    InMux I__6524 (
            .O(N__42731),
            .I(N__42725));
    Odrv4 I__6523 (
            .O(N__42728),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__6522 (
            .O(N__42725),
            .I(\uart_drone.stateZ0Z_2 ));
    InMux I__6521 (
            .O(N__42720),
            .I(N__42716));
    InMux I__6520 (
            .O(N__42719),
            .I(N__42713));
    LocalMux I__6519 (
            .O(N__42716),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__6518 (
            .O(N__42713),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__6517 (
            .O(N__42708),
            .I(N__42704));
    InMux I__6516 (
            .O(N__42707),
            .I(N__42701));
    LocalMux I__6515 (
            .O(N__42704),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__6514 (
            .O(N__42701),
            .I(\reset_module_System.countZ0Z_7 ));
    CascadeMux I__6513 (
            .O(N__42696),
            .I(N__42692));
    InMux I__6512 (
            .O(N__42695),
            .I(N__42689));
    InMux I__6511 (
            .O(N__42692),
            .I(N__42686));
    LocalMux I__6510 (
            .O(N__42689),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__6509 (
            .O(N__42686),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__6508 (
            .O(N__42681),
            .I(N__42677));
    InMux I__6507 (
            .O(N__42680),
            .I(N__42674));
    LocalMux I__6506 (
            .O(N__42677),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__6505 (
            .O(N__42674),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__6504 (
            .O(N__42669),
            .I(N__42666));
    LocalMux I__6503 (
            .O(N__42666),
            .I(N__42663));
    Odrv4 I__6502 (
            .O(N__42663),
            .I(\reset_module_System.reset6_13 ));
    InMux I__6501 (
            .O(N__42660),
            .I(N__42656));
    InMux I__6500 (
            .O(N__42659),
            .I(N__42653));
    LocalMux I__6499 (
            .O(N__42656),
            .I(\uart_drone.N_126_li ));
    LocalMux I__6498 (
            .O(N__42653),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__6497 (
            .O(N__42648),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__6496 (
            .O(N__42645),
            .I(N__42642));
    InMux I__6495 (
            .O(N__42642),
            .I(N__42638));
    InMux I__6494 (
            .O(N__42641),
            .I(N__42635));
    LocalMux I__6493 (
            .O(N__42638),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__6492 (
            .O(N__42635),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__6491 (
            .O(N__42630),
            .I(N__42627));
    LocalMux I__6490 (
            .O(N__42627),
            .I(N__42624));
    Span4Mux_v I__6489 (
            .O(N__42624),
            .I(N__42619));
    InMux I__6488 (
            .O(N__42623),
            .I(N__42614));
    InMux I__6487 (
            .O(N__42622),
            .I(N__42614));
    Odrv4 I__6486 (
            .O(N__42619),
            .I(\uart_drone.data_rdyc_1 ));
    LocalMux I__6485 (
            .O(N__42614),
            .I(\uart_drone.data_rdyc_1 ));
    CascadeMux I__6484 (
            .O(N__42609),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    InMux I__6483 (
            .O(N__42606),
            .I(N__42601));
    InMux I__6482 (
            .O(N__42605),
            .I(N__42598));
    InMux I__6481 (
            .O(N__42604),
            .I(N__42595));
    LocalMux I__6480 (
            .O(N__42601),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__6479 (
            .O(N__42598),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__6478 (
            .O(N__42595),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__6477 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__6476 (
            .O(N__42585),
            .I(\Commands_frame_decoder.WDT8lto9_3 ));
    CascadeMux I__6475 (
            .O(N__42582),
            .I(N__42577));
    CascadeMux I__6474 (
            .O(N__42581),
            .I(N__42574));
    InMux I__6473 (
            .O(N__42580),
            .I(N__42571));
    InMux I__6472 (
            .O(N__42577),
            .I(N__42568));
    InMux I__6471 (
            .O(N__42574),
            .I(N__42565));
    LocalMux I__6470 (
            .O(N__42571),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__6469 (
            .O(N__42568),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__6468 (
            .O(N__42565),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__6467 (
            .O(N__42558),
            .I(N__42553));
    InMux I__6466 (
            .O(N__42557),
            .I(N__42550));
    InMux I__6465 (
            .O(N__42556),
            .I(N__42547));
    LocalMux I__6464 (
            .O(N__42553),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__6463 (
            .O(N__42550),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__6462 (
            .O(N__42547),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__6461 (
            .O(N__42540),
            .I(N__42537));
    LocalMux I__6460 (
            .O(N__42537),
            .I(\Commands_frame_decoder.state_0_sqmuxacf1 ));
    CascadeMux I__6459 (
            .O(N__42534),
            .I(\Commands_frame_decoder.WDT8lt12_0_cascade_ ));
    InMux I__6458 (
            .O(N__42531),
            .I(N__42527));
    CascadeMux I__6457 (
            .O(N__42530),
            .I(N__42524));
    LocalMux I__6456 (
            .O(N__42527),
            .I(N__42521));
    InMux I__6455 (
            .O(N__42524),
            .I(N__42518));
    Odrv4 I__6454 (
            .O(N__42521),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__6453 (
            .O(N__42518),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__6452 (
            .O(N__42513),
            .I(N__42507));
    InMux I__6451 (
            .O(N__42512),
            .I(N__42504));
    InMux I__6450 (
            .O(N__42511),
            .I(N__42499));
    InMux I__6449 (
            .O(N__42510),
            .I(N__42499));
    LocalMux I__6448 (
            .O(N__42507),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__6447 (
            .O(N__42504),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__6446 (
            .O(N__42499),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__6445 (
            .O(N__42492),
            .I(N__42486));
    InMux I__6444 (
            .O(N__42491),
            .I(N__42481));
    InMux I__6443 (
            .O(N__42490),
            .I(N__42481));
    InMux I__6442 (
            .O(N__42489),
            .I(N__42478));
    LocalMux I__6441 (
            .O(N__42486),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__6440 (
            .O(N__42481),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__6439 (
            .O(N__42478),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__6438 (
            .O(N__42471),
            .I(N__42465));
    InMux I__6437 (
            .O(N__42470),
            .I(N__42460));
    InMux I__6436 (
            .O(N__42469),
            .I(N__42460));
    InMux I__6435 (
            .O(N__42468),
            .I(N__42457));
    LocalMux I__6434 (
            .O(N__42465),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__6433 (
            .O(N__42460),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__6432 (
            .O(N__42457),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__6431 (
            .O(N__42450),
            .I(N__42442));
    InMux I__6430 (
            .O(N__42449),
            .I(N__42442));
    InMux I__6429 (
            .O(N__42448),
            .I(N__42437));
    InMux I__6428 (
            .O(N__42447),
            .I(N__42437));
    LocalMux I__6427 (
            .O(N__42442),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__6426 (
            .O(N__42437),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__6425 (
            .O(N__42432),
            .I(N__42429));
    LocalMux I__6424 (
            .O(N__42429),
            .I(N__42424));
    InMux I__6423 (
            .O(N__42428),
            .I(N__42419));
    InMux I__6422 (
            .O(N__42427),
            .I(N__42416));
    Span4Mux_h I__6421 (
            .O(N__42424),
            .I(N__42413));
    InMux I__6420 (
            .O(N__42423),
            .I(N__42410));
    InMux I__6419 (
            .O(N__42422),
            .I(N__42407));
    LocalMux I__6418 (
            .O(N__42419),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__6417 (
            .O(N__42416),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__6416 (
            .O(N__42413),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__6415 (
            .O(N__42410),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__6414 (
            .O(N__42407),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    CascadeMux I__6413 (
            .O(N__42396),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ));
    InMux I__6412 (
            .O(N__42393),
            .I(N__42387));
    CascadeMux I__6411 (
            .O(N__42392),
            .I(N__42384));
    InMux I__6410 (
            .O(N__42391),
            .I(N__42380));
    InMux I__6409 (
            .O(N__42390),
            .I(N__42377));
    LocalMux I__6408 (
            .O(N__42387),
            .I(N__42374));
    InMux I__6407 (
            .O(N__42384),
            .I(N__42369));
    InMux I__6406 (
            .O(N__42383),
            .I(N__42369));
    LocalMux I__6405 (
            .O(N__42380),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__6404 (
            .O(N__42377),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__6403 (
            .O(N__42374),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__6402 (
            .O(N__42369),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__6401 (
            .O(N__42360),
            .I(N__42357));
    LocalMux I__6400 (
            .O(N__42357),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0 ));
    CascadeMux I__6399 (
            .O(N__42354),
            .I(N__42349));
    InMux I__6398 (
            .O(N__42353),
            .I(N__42343));
    InMux I__6397 (
            .O(N__42352),
            .I(N__42343));
    InMux I__6396 (
            .O(N__42349),
            .I(N__42337));
    InMux I__6395 (
            .O(N__42348),
            .I(N__42337));
    LocalMux I__6394 (
            .O(N__42343),
            .I(N__42334));
    InMux I__6393 (
            .O(N__42342),
            .I(N__42331));
    LocalMux I__6392 (
            .O(N__42337),
            .I(\uart_drone.N_143 ));
    Odrv4 I__6391 (
            .O(N__42334),
            .I(\uart_drone.N_143 ));
    LocalMux I__6390 (
            .O(N__42331),
            .I(\uart_drone.N_143 ));
    CascadeMux I__6389 (
            .O(N__42324),
            .I(N__42320));
    InMux I__6388 (
            .O(N__42323),
            .I(N__42313));
    InMux I__6387 (
            .O(N__42320),
            .I(N__42313));
    InMux I__6386 (
            .O(N__42319),
            .I(N__42308));
    InMux I__6385 (
            .O(N__42318),
            .I(N__42308));
    LocalMux I__6384 (
            .O(N__42313),
            .I(N__42302));
    LocalMux I__6383 (
            .O(N__42308),
            .I(N__42302));
    InMux I__6382 (
            .O(N__42307),
            .I(N__42299));
    Odrv12 I__6381 (
            .O(N__42302),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__6380 (
            .O(N__42299),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    InMux I__6379 (
            .O(N__42294),
            .I(N__42291));
    LocalMux I__6378 (
            .O(N__42291),
            .I(N__42288));
    Span4Mux_h I__6377 (
            .O(N__42288),
            .I(N__42285));
    Odrv4 I__6376 (
            .O(N__42285),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10 ));
    InMux I__6375 (
            .O(N__42282),
            .I(N__42279));
    LocalMux I__6374 (
            .O(N__42279),
            .I(N__42276));
    Odrv4 I__6373 (
            .O(N__42276),
            .I(\pid_front.un10lt11_0 ));
    CascadeMux I__6372 (
            .O(N__42273),
            .I(N__42268));
    InMux I__6371 (
            .O(N__42272),
            .I(N__42265));
    InMux I__6370 (
            .O(N__42271),
            .I(N__42262));
    InMux I__6369 (
            .O(N__42268),
            .I(N__42259));
    LocalMux I__6368 (
            .O(N__42265),
            .I(N__42256));
    LocalMux I__6367 (
            .O(N__42262),
            .I(N__42253));
    LocalMux I__6366 (
            .O(N__42259),
            .I(N__42250));
    Span4Mux_h I__6365 (
            .O(N__42256),
            .I(N__42247));
    Span4Mux_v I__6364 (
            .O(N__42253),
            .I(N__42242));
    Span4Mux_v I__6363 (
            .O(N__42250),
            .I(N__42242));
    Odrv4 I__6362 (
            .O(N__42247),
            .I(\pid_front.un10lto12 ));
    Odrv4 I__6361 (
            .O(N__42242),
            .I(\pid_front.un10lto12 ));
    InMux I__6360 (
            .O(N__42237),
            .I(N__42234));
    LocalMux I__6359 (
            .O(N__42234),
            .I(\pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ));
    InMux I__6358 (
            .O(N__42231),
            .I(N__42228));
    LocalMux I__6357 (
            .O(N__42228),
            .I(N__42225));
    Odrv12 I__6356 (
            .O(N__42225),
            .I(\pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ));
    InMux I__6355 (
            .O(N__42222),
            .I(N__42218));
    InMux I__6354 (
            .O(N__42221),
            .I(N__42215));
    LocalMux I__6353 (
            .O(N__42218),
            .I(drone_H_disp_front_1));
    LocalMux I__6352 (
            .O(N__42215),
            .I(drone_H_disp_front_1));
    InMux I__6351 (
            .O(N__42210),
            .I(N__42206));
    InMux I__6350 (
            .O(N__42209),
            .I(N__42203));
    LocalMux I__6349 (
            .O(N__42206),
            .I(drone_H_disp_front_3));
    LocalMux I__6348 (
            .O(N__42203),
            .I(drone_H_disp_front_3));
    IoInMux I__6347 (
            .O(N__42198),
            .I(N__42195));
    LocalMux I__6346 (
            .O(N__42195),
            .I(N__42192));
    Span4Mux_s0_v I__6345 (
            .O(N__42192),
            .I(N__42189));
    Span4Mux_h I__6344 (
            .O(N__42189),
            .I(N__42186));
    Odrv4 I__6343 (
            .O(N__42186),
            .I(\pid_front.state_RNIPKTDZ0Z_0 ));
    InMux I__6342 (
            .O(N__42183),
            .I(N__42180));
    LocalMux I__6341 (
            .O(N__42180),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__6340 (
            .O(N__42177),
            .I(N__42174));
    LocalMux I__6339 (
            .O(N__42174),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__6338 (
            .O(N__42171),
            .I(N__42166));
    InMux I__6337 (
            .O(N__42170),
            .I(N__42163));
    InMux I__6336 (
            .O(N__42169),
            .I(N__42160));
    LocalMux I__6335 (
            .O(N__42166),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__6334 (
            .O(N__42163),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__6333 (
            .O(N__42160),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__6332 (
            .O(N__42153),
            .I(N__42148));
    InMux I__6331 (
            .O(N__42152),
            .I(N__42145));
    InMux I__6330 (
            .O(N__42151),
            .I(N__42142));
    LocalMux I__6329 (
            .O(N__42148),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__6328 (
            .O(N__42145),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__6327 (
            .O(N__42142),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    CascadeMux I__6326 (
            .O(N__42135),
            .I(N__42130));
    CascadeMux I__6325 (
            .O(N__42134),
            .I(N__42127));
    InMux I__6324 (
            .O(N__42133),
            .I(N__42124));
    InMux I__6323 (
            .O(N__42130),
            .I(N__42121));
    InMux I__6322 (
            .O(N__42127),
            .I(N__42118));
    LocalMux I__6321 (
            .O(N__42124),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__6320 (
            .O(N__42121),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__6319 (
            .O(N__42118),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__6318 (
            .O(N__42111),
            .I(N__42106));
    InMux I__6317 (
            .O(N__42110),
            .I(N__42103));
    InMux I__6316 (
            .O(N__42109),
            .I(N__42100));
    LocalMux I__6315 (
            .O(N__42106),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__6314 (
            .O(N__42103),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__6313 (
            .O(N__42100),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__6312 (
            .O(N__42093),
            .I(N__42090));
    LocalMux I__6311 (
            .O(N__42090),
            .I(N__42087));
    Odrv12 I__6310 (
            .O(N__42087),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    InMux I__6309 (
            .O(N__42084),
            .I(N__42080));
    InMux I__6308 (
            .O(N__42083),
            .I(N__42077));
    LocalMux I__6307 (
            .O(N__42080),
            .I(N__42074));
    LocalMux I__6306 (
            .O(N__42077),
            .I(N__42071));
    Odrv12 I__6305 (
            .O(N__42074),
            .I(\pid_front.error_i_acumm_preregZ0Z_0 ));
    Odrv4 I__6304 (
            .O(N__42071),
            .I(\pid_front.error_i_acumm_preregZ0Z_0 ));
    CascadeMux I__6303 (
            .O(N__42066),
            .I(N__42062));
    CascadeMux I__6302 (
            .O(N__42065),
            .I(N__42059));
    InMux I__6301 (
            .O(N__42062),
            .I(N__42056));
    InMux I__6300 (
            .O(N__42059),
            .I(N__42053));
    LocalMux I__6299 (
            .O(N__42056),
            .I(\pid_front.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__6298 (
            .O(N__42053),
            .I(\pid_front.error_i_acumm_preregZ0Z_21 ));
    CascadeMux I__6297 (
            .O(N__42048),
            .I(N__42045));
    InMux I__6296 (
            .O(N__42045),
            .I(N__42041));
    InMux I__6295 (
            .O(N__42044),
            .I(N__42038));
    LocalMux I__6294 (
            .O(N__42041),
            .I(\pid_front.error_i_acumm_preregZ0Z_17 ));
    LocalMux I__6293 (
            .O(N__42038),
            .I(\pid_front.error_i_acumm_preregZ0Z_17 ));
    InMux I__6292 (
            .O(N__42033),
            .I(N__42027));
    InMux I__6291 (
            .O(N__42032),
            .I(N__42027));
    LocalMux I__6290 (
            .O(N__42027),
            .I(\pid_front.error_i_acumm_preregZ0Z_22 ));
    InMux I__6289 (
            .O(N__42024),
            .I(N__42018));
    InMux I__6288 (
            .O(N__42023),
            .I(N__42018));
    LocalMux I__6287 (
            .O(N__42018),
            .I(\pid_front.error_i_acumm_preregZ0Z_23 ));
    CascadeMux I__6286 (
            .O(N__42015),
            .I(N__42012));
    InMux I__6285 (
            .O(N__42012),
            .I(N__42006));
    InMux I__6284 (
            .O(N__42011),
            .I(N__42006));
    LocalMux I__6283 (
            .O(N__42006),
            .I(\pid_front.error_i_acumm_preregZ0Z_24 ));
    InMux I__6282 (
            .O(N__42003),
            .I(N__41999));
    InMux I__6281 (
            .O(N__42002),
            .I(N__41996));
    LocalMux I__6280 (
            .O(N__41999),
            .I(\pid_front.error_i_acumm_preregZ0Z_16 ));
    LocalMux I__6279 (
            .O(N__41996),
            .I(\pid_front.error_i_acumm_preregZ0Z_16 ));
    CascadeMux I__6278 (
            .O(N__41991),
            .I(N__41987));
    InMux I__6277 (
            .O(N__41990),
            .I(N__41982));
    InMux I__6276 (
            .O(N__41987),
            .I(N__41982));
    LocalMux I__6275 (
            .O(N__41982),
            .I(\pid_front.error_i_acumm_preregZ0Z_25 ));
    InMux I__6274 (
            .O(N__41979),
            .I(N__41975));
    InMux I__6273 (
            .O(N__41978),
            .I(N__41972));
    LocalMux I__6272 (
            .O(N__41975),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    LocalMux I__6271 (
            .O(N__41972),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    CascadeMux I__6270 (
            .O(N__41967),
            .I(\pid_front.un1_pid_prereg_0_19_cascade_ ));
    CascadeMux I__6269 (
            .O(N__41964),
            .I(N__41961));
    InMux I__6268 (
            .O(N__41961),
            .I(N__41952));
    InMux I__6267 (
            .O(N__41960),
            .I(N__41952));
    InMux I__6266 (
            .O(N__41959),
            .I(N__41952));
    LocalMux I__6265 (
            .O(N__41952),
            .I(\pid_front.un1_pid_prereg_0_17 ));
    CascadeMux I__6264 (
            .O(N__41949),
            .I(\pid_front.un1_pid_prereg_0_25_cascade_ ));
    InMux I__6263 (
            .O(N__41946),
            .I(N__41942));
    InMux I__6262 (
            .O(N__41945),
            .I(N__41939));
    LocalMux I__6261 (
            .O(N__41942),
            .I(\pid_front.un1_pid_prereg_0_24 ));
    LocalMux I__6260 (
            .O(N__41939),
            .I(\pid_front.un1_pid_prereg_0_24 ));
    CascadeMux I__6259 (
            .O(N__41934),
            .I(\pid_front.un1_pid_prereg_0_26_cascade_ ));
    CascadeMux I__6258 (
            .O(N__41931),
            .I(N__41928));
    InMux I__6257 (
            .O(N__41928),
            .I(N__41922));
    InMux I__6256 (
            .O(N__41927),
            .I(N__41922));
    LocalMux I__6255 (
            .O(N__41922),
            .I(\pid_front.un1_pid_prereg_0_26 ));
    InMux I__6254 (
            .O(N__41919),
            .I(N__41906));
    InMux I__6253 (
            .O(N__41918),
            .I(N__41906));
    InMux I__6252 (
            .O(N__41917),
            .I(N__41906));
    InMux I__6251 (
            .O(N__41916),
            .I(N__41906));
    InMux I__6250 (
            .O(N__41915),
            .I(N__41903));
    LocalMux I__6249 (
            .O(N__41906),
            .I(\pid_front.un1_pid_prereg_0_25 ));
    LocalMux I__6248 (
            .O(N__41903),
            .I(\pid_front.un1_pid_prereg_0_25 ));
    CascadeMux I__6247 (
            .O(N__41898),
            .I(N__41894));
    CascadeMux I__6246 (
            .O(N__41897),
            .I(N__41890));
    InMux I__6245 (
            .O(N__41894),
            .I(N__41887));
    InMux I__6244 (
            .O(N__41893),
            .I(N__41882));
    InMux I__6243 (
            .O(N__41890),
            .I(N__41882));
    LocalMux I__6242 (
            .O(N__41887),
            .I(N__41879));
    LocalMux I__6241 (
            .O(N__41882),
            .I(N__41876));
    Odrv4 I__6240 (
            .O(N__41879),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    Odrv4 I__6239 (
            .O(N__41876),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    InMux I__6238 (
            .O(N__41871),
            .I(N__41866));
    InMux I__6237 (
            .O(N__41870),
            .I(N__41861));
    InMux I__6236 (
            .O(N__41869),
            .I(N__41861));
    LocalMux I__6235 (
            .O(N__41866),
            .I(N__41858));
    LocalMux I__6234 (
            .O(N__41861),
            .I(N__41855));
    Odrv4 I__6233 (
            .O(N__41858),
            .I(\pid_front.error_i_acumm_preregZ0Z_13 ));
    Odrv4 I__6232 (
            .O(N__41855),
            .I(\pid_front.error_i_acumm_preregZ0Z_13 ));
    CascadeMux I__6231 (
            .O(N__41850),
            .I(N__41845));
    CascadeMux I__6230 (
            .O(N__41849),
            .I(N__41841));
    InMux I__6229 (
            .O(N__41848),
            .I(N__41826));
    InMux I__6228 (
            .O(N__41845),
            .I(N__41826));
    InMux I__6227 (
            .O(N__41844),
            .I(N__41826));
    InMux I__6226 (
            .O(N__41841),
            .I(N__41826));
    InMux I__6225 (
            .O(N__41840),
            .I(N__41826));
    InMux I__6224 (
            .O(N__41839),
            .I(N__41826));
    LocalMux I__6223 (
            .O(N__41826),
            .I(\pid_front.error_i_acumm_2_sqmuxa_1 ));
    CascadeMux I__6222 (
            .O(N__41823),
            .I(N__41820));
    InMux I__6221 (
            .O(N__41820),
            .I(N__41817));
    LocalMux I__6220 (
            .O(N__41817),
            .I(N__41814));
    Span4Mux_v I__6219 (
            .O(N__41814),
            .I(N__41809));
    InMux I__6218 (
            .O(N__41813),
            .I(N__41804));
    InMux I__6217 (
            .O(N__41812),
            .I(N__41804));
    Odrv4 I__6216 (
            .O(N__41809),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__6215 (
            .O(N__41804),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__6214 (
            .O(N__41799),
            .I(\pid_front.un1_pid_prereg_0_24_cascade_ ));
    CascadeMux I__6213 (
            .O(N__41796),
            .I(\pid_front.un1_pid_prereg_0_16_cascade_ ));
    InMux I__6212 (
            .O(N__41793),
            .I(N__41787));
    InMux I__6211 (
            .O(N__41792),
            .I(N__41787));
    LocalMux I__6210 (
            .O(N__41787),
            .I(\pid_front.un1_pid_prereg_0_16 ));
    InMux I__6209 (
            .O(N__41784),
            .I(N__41775));
    InMux I__6208 (
            .O(N__41783),
            .I(N__41775));
    InMux I__6207 (
            .O(N__41782),
            .I(N__41775));
    LocalMux I__6206 (
            .O(N__41775),
            .I(\pid_front.error_i_acumm_3_sqmuxa ));
    InMux I__6205 (
            .O(N__41772),
            .I(N__41769));
    LocalMux I__6204 (
            .O(N__41769),
            .I(N__41766));
    Span4Mux_v I__6203 (
            .O(N__41766),
            .I(N__41761));
    InMux I__6202 (
            .O(N__41765),
            .I(N__41756));
    InMux I__6201 (
            .O(N__41764),
            .I(N__41756));
    Odrv4 I__6200 (
            .O(N__41761),
            .I(\pid_front.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__6199 (
            .O(N__41756),
            .I(\pid_front.error_i_acumm_preregZ0Z_9 ));
    InMux I__6198 (
            .O(N__41751),
            .I(N__41748));
    LocalMux I__6197 (
            .O(N__41748),
            .I(N__41744));
    InMux I__6196 (
            .O(N__41747),
            .I(N__41741));
    Odrv4 I__6195 (
            .O(N__41744),
            .I(\pid_front.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__6194 (
            .O(N__41741),
            .I(\pid_front.error_i_acumm_preregZ0Z_1 ));
    InMux I__6193 (
            .O(N__41736),
            .I(N__41733));
    LocalMux I__6192 (
            .O(N__41733),
            .I(N__41729));
    CascadeMux I__6191 (
            .O(N__41732),
            .I(N__41726));
    Span4Mux_v I__6190 (
            .O(N__41729),
            .I(N__41723));
    InMux I__6189 (
            .O(N__41726),
            .I(N__41720));
    Odrv4 I__6188 (
            .O(N__41723),
            .I(\pid_front.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__6187 (
            .O(N__41720),
            .I(\pid_front.error_i_acumm_preregZ0Z_2 ));
    InMux I__6186 (
            .O(N__41715),
            .I(N__41712));
    LocalMux I__6185 (
            .O(N__41712),
            .I(N__41709));
    Odrv4 I__6184 (
            .O(N__41709),
            .I(\pid_front.error_i_acumm16lto27_13 ));
    InMux I__6183 (
            .O(N__41706),
            .I(N__41703));
    LocalMux I__6182 (
            .O(N__41703),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ));
    CascadeMux I__6181 (
            .O(N__41700),
            .I(\pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ));
    CascadeMux I__6180 (
            .O(N__41697),
            .I(\pid_front.error_i_acumm_2_sqmuxa_cascade_ ));
    CascadeMux I__6179 (
            .O(N__41694),
            .I(N__41690));
    InMux I__6178 (
            .O(N__41693),
            .I(N__41686));
    InMux I__6177 (
            .O(N__41690),
            .I(N__41681));
    InMux I__6176 (
            .O(N__41689),
            .I(N__41681));
    LocalMux I__6175 (
            .O(N__41686),
            .I(N__41678));
    LocalMux I__6174 (
            .O(N__41681),
            .I(N__41675));
    Odrv12 I__6173 (
            .O(N__41678),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    Odrv4 I__6172 (
            .O(N__41675),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    CascadeMux I__6171 (
            .O(N__41670),
            .I(N__41667));
    InMux I__6170 (
            .O(N__41667),
            .I(N__41662));
    InMux I__6169 (
            .O(N__41666),
            .I(N__41657));
    InMux I__6168 (
            .O(N__41665),
            .I(N__41657));
    LocalMux I__6167 (
            .O(N__41662),
            .I(N__41654));
    LocalMux I__6166 (
            .O(N__41657),
            .I(N__41651));
    Odrv12 I__6165 (
            .O(N__41654),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    Odrv4 I__6164 (
            .O(N__41651),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    InMux I__6163 (
            .O(N__41646),
            .I(N__41641));
    InMux I__6162 (
            .O(N__41645),
            .I(N__41638));
    InMux I__6161 (
            .O(N__41644),
            .I(N__41635));
    LocalMux I__6160 (
            .O(N__41641),
            .I(N__41632));
    LocalMux I__6159 (
            .O(N__41638),
            .I(N__41627));
    LocalMux I__6158 (
            .O(N__41635),
            .I(N__41627));
    Odrv12 I__6157 (
            .O(N__41632),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    Odrv4 I__6156 (
            .O(N__41627),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    CascadeMux I__6155 (
            .O(N__41622),
            .I(\pid_front.un1_pid_prereg_79_cascade_ ));
    CascadeMux I__6154 (
            .O(N__41619),
            .I(N__41616));
    InMux I__6153 (
            .O(N__41616),
            .I(N__41610));
    InMux I__6152 (
            .O(N__41615),
            .I(N__41605));
    InMux I__6151 (
            .O(N__41614),
            .I(N__41605));
    InMux I__6150 (
            .O(N__41613),
            .I(N__41602));
    LocalMux I__6149 (
            .O(N__41610),
            .I(\pid_front.error_d_regZ0Z_7 ));
    LocalMux I__6148 (
            .O(N__41605),
            .I(\pid_front.error_d_regZ0Z_7 ));
    LocalMux I__6147 (
            .O(N__41602),
            .I(\pid_front.error_d_regZ0Z_7 ));
    InMux I__6146 (
            .O(N__41595),
            .I(N__41590));
    InMux I__6145 (
            .O(N__41594),
            .I(N__41585));
    InMux I__6144 (
            .O(N__41593),
            .I(N__41585));
    LocalMux I__6143 (
            .O(N__41590),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    LocalMux I__6142 (
            .O(N__41585),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    InMux I__6141 (
            .O(N__41580),
            .I(N__41577));
    LocalMux I__6140 (
            .O(N__41577),
            .I(N__41574));
    Span4Mux_h I__6139 (
            .O(N__41574),
            .I(N__41569));
    InMux I__6138 (
            .O(N__41573),
            .I(N__41564));
    InMux I__6137 (
            .O(N__41572),
            .I(N__41564));
    Odrv4 I__6136 (
            .O(N__41569),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__6135 (
            .O(N__41564),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    CascadeMux I__6134 (
            .O(N__41559),
            .I(\pid_front.error_i_acumm_3_sqmuxa_cascade_ ));
    InMux I__6133 (
            .O(N__41556),
            .I(N__41553));
    LocalMux I__6132 (
            .O(N__41553),
            .I(N__41548));
    InMux I__6131 (
            .O(N__41552),
            .I(N__41545));
    InMux I__6130 (
            .O(N__41551),
            .I(N__41542));
    Span4Mux_h I__6129 (
            .O(N__41548),
            .I(N__41539));
    LocalMux I__6128 (
            .O(N__41545),
            .I(N__41534));
    LocalMux I__6127 (
            .O(N__41542),
            .I(N__41534));
    Odrv4 I__6126 (
            .O(N__41539),
            .I(\pid_front.error_i_acumm_preregZ0Z_8 ));
    Odrv4 I__6125 (
            .O(N__41534),
            .I(\pid_front.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__6124 (
            .O(N__41529),
            .I(\pid_front.N_1698_i_cascade_ ));
    InMux I__6123 (
            .O(N__41526),
            .I(N__41523));
    LocalMux I__6122 (
            .O(N__41523),
            .I(N__41520));
    Span4Mux_h I__6121 (
            .O(N__41520),
            .I(N__41517));
    Odrv4 I__6120 (
            .O(N__41517),
            .I(\pid_front.error_d_reg_prev_esr_RNIUO6U_0Z0Z_12 ));
    CascadeMux I__6119 (
            .O(N__41514),
            .I(\pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13_cascade_ ));
    InMux I__6118 (
            .O(N__41511),
            .I(N__41508));
    LocalMux I__6117 (
            .O(N__41508),
            .I(\pid_front.error_p_reg_esr_RNIROQ33Z0Z_12 ));
    InMux I__6116 (
            .O(N__41505),
            .I(N__41499));
    InMux I__6115 (
            .O(N__41504),
            .I(N__41499));
    LocalMux I__6114 (
            .O(N__41499),
            .I(N__41496));
    Sp12to4 I__6113 (
            .O(N__41496),
            .I(N__41493));
    Odrv12 I__6112 (
            .O(N__41493),
            .I(\pid_front.error_p_regZ0Z_14 ));
    InMux I__6111 (
            .O(N__41490),
            .I(N__41484));
    InMux I__6110 (
            .O(N__41489),
            .I(N__41484));
    LocalMux I__6109 (
            .O(N__41484),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    InMux I__6108 (
            .O(N__41481),
            .I(N__41478));
    LocalMux I__6107 (
            .O(N__41478),
            .I(\pid_front.N_1674_i ));
    InMux I__6106 (
            .O(N__41475),
            .I(N__41471));
    InMux I__6105 (
            .O(N__41474),
            .I(N__41468));
    LocalMux I__6104 (
            .O(N__41471),
            .I(N__41465));
    LocalMux I__6103 (
            .O(N__41468),
            .I(N__41462));
    Span4Mux_h I__6102 (
            .O(N__41465),
            .I(N__41459));
    Span4Mux_h I__6101 (
            .O(N__41462),
            .I(N__41456));
    Span4Mux_h I__6100 (
            .O(N__41459),
            .I(N__41453));
    Span4Mux_h I__6099 (
            .O(N__41456),
            .I(N__41450));
    Odrv4 I__6098 (
            .O(N__41453),
            .I(\pid_front.error_p_regZ0Z_8 ));
    Odrv4 I__6097 (
            .O(N__41450),
            .I(\pid_front.error_p_regZ0Z_8 ));
    CascadeMux I__6096 (
            .O(N__41445),
            .I(\pid_front.N_1674_i_cascade_ ));
    InMux I__6095 (
            .O(N__41442),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    CascadeMux I__6094 (
            .O(N__41439),
            .I(N__41436));
    InMux I__6093 (
            .O(N__41436),
            .I(N__41433));
    LocalMux I__6092 (
            .O(N__41433),
            .I(N__41429));
    InMux I__6091 (
            .O(N__41432),
            .I(N__41424));
    Span4Mux_h I__6090 (
            .O(N__41429),
            .I(N__41421));
    InMux I__6089 (
            .O(N__41428),
            .I(N__41416));
    InMux I__6088 (
            .O(N__41427),
            .I(N__41416));
    LocalMux I__6087 (
            .O(N__41424),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    Odrv4 I__6086 (
            .O(N__41421),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__6085 (
            .O(N__41416),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    InMux I__6084 (
            .O(N__41409),
            .I(N__41402));
    InMux I__6083 (
            .O(N__41408),
            .I(N__41402));
    InMux I__6082 (
            .O(N__41407),
            .I(N__41399));
    LocalMux I__6081 (
            .O(N__41402),
            .I(\pid_front.pid_preregZ0Z_14 ));
    LocalMux I__6080 (
            .O(N__41399),
            .I(\pid_front.pid_preregZ0Z_14 ));
    CascadeMux I__6079 (
            .O(N__41394),
            .I(\pid_front.pid_prereg_esr_RNIQ6EVZ0Z_17_cascade_ ));
    CascadeMux I__6078 (
            .O(N__41391),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0_cascade_ ));
    InMux I__6077 (
            .O(N__41388),
            .I(N__41384));
    InMux I__6076 (
            .O(N__41387),
            .I(N__41381));
    LocalMux I__6075 (
            .O(N__41384),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    LocalMux I__6074 (
            .O(N__41381),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    InMux I__6073 (
            .O(N__41376),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__6072 (
            .O(N__41373),
            .I(N__41369));
    InMux I__6071 (
            .O(N__41372),
            .I(N__41366));
    LocalMux I__6070 (
            .O(N__41369),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__6069 (
            .O(N__41366),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__6068 (
            .O(N__41361),
            .I(bfn_9_14_0_));
    InMux I__6067 (
            .O(N__41358),
            .I(N__41354));
    InMux I__6066 (
            .O(N__41357),
            .I(N__41351));
    LocalMux I__6065 (
            .O(N__41354),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__6064 (
            .O(N__41351),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__6063 (
            .O(N__41346),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    CascadeMux I__6062 (
            .O(N__41343),
            .I(N__41339));
    InMux I__6061 (
            .O(N__41342),
            .I(N__41335));
    InMux I__6060 (
            .O(N__41339),
            .I(N__41330));
    InMux I__6059 (
            .O(N__41338),
            .I(N__41330));
    LocalMux I__6058 (
            .O(N__41335),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__6057 (
            .O(N__41330),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__6056 (
            .O(N__41325),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__6055 (
            .O(N__41322),
            .I(N__41316));
    InMux I__6054 (
            .O(N__41321),
            .I(N__41309));
    InMux I__6053 (
            .O(N__41320),
            .I(N__41309));
    InMux I__6052 (
            .O(N__41319),
            .I(N__41309));
    LocalMux I__6051 (
            .O(N__41316),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__6050 (
            .O(N__41309),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__6049 (
            .O(N__41304),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    CascadeMux I__6048 (
            .O(N__41301),
            .I(N__41296));
    InMux I__6047 (
            .O(N__41300),
            .I(N__41292));
    InMux I__6046 (
            .O(N__41299),
            .I(N__41285));
    InMux I__6045 (
            .O(N__41296),
            .I(N__41285));
    InMux I__6044 (
            .O(N__41295),
            .I(N__41285));
    LocalMux I__6043 (
            .O(N__41292),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__6042 (
            .O(N__41285),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__6041 (
            .O(N__41280),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    InMux I__6040 (
            .O(N__41277),
            .I(N__41273));
    InMux I__6039 (
            .O(N__41276),
            .I(N__41269));
    LocalMux I__6038 (
            .O(N__41273),
            .I(N__41266));
    InMux I__6037 (
            .O(N__41272),
            .I(N__41263));
    LocalMux I__6036 (
            .O(N__41269),
            .I(N__41258));
    Span4Mux_v I__6035 (
            .O(N__41266),
            .I(N__41258));
    LocalMux I__6034 (
            .O(N__41263),
            .I(N__41255));
    Sp12to4 I__6033 (
            .O(N__41258),
            .I(N__41251));
    Span4Mux_h I__6032 (
            .O(N__41255),
            .I(N__41248));
    InMux I__6031 (
            .O(N__41254),
            .I(N__41245));
    Odrv12 I__6030 (
            .O(N__41251),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    Odrv4 I__6029 (
            .O(N__41248),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__6028 (
            .O(N__41245),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__6027 (
            .O(N__41238),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__6026 (
            .O(N__41235),
            .I(N__41232));
    LocalMux I__6025 (
            .O(N__41232),
            .I(N__41228));
    InMux I__6024 (
            .O(N__41231),
            .I(N__41223));
    Span4Mux_h I__6023 (
            .O(N__41228),
            .I(N__41220));
    InMux I__6022 (
            .O(N__41227),
            .I(N__41215));
    InMux I__6021 (
            .O(N__41226),
            .I(N__41215));
    LocalMux I__6020 (
            .O(N__41223),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    Odrv4 I__6019 (
            .O(N__41220),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__6018 (
            .O(N__41215),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__6017 (
            .O(N__41208),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__6016 (
            .O(N__41205),
            .I(N__41201));
    InMux I__6015 (
            .O(N__41204),
            .I(N__41198));
    LocalMux I__6014 (
            .O(N__41201),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    LocalMux I__6013 (
            .O(N__41198),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    CascadeMux I__6012 (
            .O(N__41193),
            .I(N__41189));
    CascadeMux I__6011 (
            .O(N__41192),
            .I(N__41185));
    InMux I__6010 (
            .O(N__41189),
            .I(N__41181));
    InMux I__6009 (
            .O(N__41188),
            .I(N__41178));
    InMux I__6008 (
            .O(N__41185),
            .I(N__41175));
    InMux I__6007 (
            .O(N__41184),
            .I(N__41172));
    LocalMux I__6006 (
            .O(N__41181),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__6005 (
            .O(N__41178),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__6004 (
            .O(N__41175),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__6003 (
            .O(N__41172),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    CascadeMux I__6002 (
            .O(N__41163),
            .I(N__41159));
    InMux I__6001 (
            .O(N__41162),
            .I(N__41156));
    InMux I__6000 (
            .O(N__41159),
            .I(N__41153));
    LocalMux I__5999 (
            .O(N__41156),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__5998 (
            .O(N__41153),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__5997 (
            .O(N__41148),
            .I(N__41145));
    LocalMux I__5996 (
            .O(N__41145),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__5995 (
            .O(N__41142),
            .I(N__41139));
    LocalMux I__5994 (
            .O(N__41139),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__5993 (
            .O(N__41136),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__5992 (
            .O(N__41133),
            .I(N__41130));
    LocalMux I__5991 (
            .O(N__41130),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__5990 (
            .O(N__41127),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__5989 (
            .O(N__41124),
            .I(N__41121));
    LocalMux I__5988 (
            .O(N__41121),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__5987 (
            .O(N__41118),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__5986 (
            .O(N__41115),
            .I(N__41111));
    InMux I__5985 (
            .O(N__41114),
            .I(N__41108));
    LocalMux I__5984 (
            .O(N__41111),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    LocalMux I__5983 (
            .O(N__41108),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__5982 (
            .O(N__41103),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__5981 (
            .O(N__41100),
            .I(N__41096));
    InMux I__5980 (
            .O(N__41099),
            .I(N__41093));
    LocalMux I__5979 (
            .O(N__41096),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    LocalMux I__5978 (
            .O(N__41093),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    InMux I__5977 (
            .O(N__41088),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__5976 (
            .O(N__41085),
            .I(N__41081));
    InMux I__5975 (
            .O(N__41084),
            .I(N__41078));
    LocalMux I__5974 (
            .O(N__41081),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    LocalMux I__5973 (
            .O(N__41078),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__5972 (
            .O(N__41073),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    CascadeMux I__5971 (
            .O(N__41070),
            .I(N__41067));
    InMux I__5970 (
            .O(N__41067),
            .I(N__41064));
    LocalMux I__5969 (
            .O(N__41064),
            .I(N__41060));
    InMux I__5968 (
            .O(N__41063),
            .I(N__41057));
    Span4Mux_h I__5967 (
            .O(N__41060),
            .I(N__41054));
    LocalMux I__5966 (
            .O(N__41057),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__5965 (
            .O(N__41054),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__5964 (
            .O(N__41049),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__5963 (
            .O(N__41046),
            .I(N__41042));
    InMux I__5962 (
            .O(N__41045),
            .I(N__41039));
    LocalMux I__5961 (
            .O(N__41042),
            .I(N__41036));
    LocalMux I__5960 (
            .O(N__41039),
            .I(\reset_module_System.countZ0Z_19 ));
    Odrv4 I__5959 (
            .O(N__41036),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__5958 (
            .O(N__41031),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__5957 (
            .O(N__41028),
            .I(N__41025));
    InMux I__5956 (
            .O(N__41025),
            .I(N__41021));
    InMux I__5955 (
            .O(N__41024),
            .I(N__41018));
    LocalMux I__5954 (
            .O(N__41021),
            .I(N__41015));
    LocalMux I__5953 (
            .O(N__41018),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__5952 (
            .O(N__41015),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__5951 (
            .O(N__41010),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__5950 (
            .O(N__41007),
            .I(\reset_module_System.count_1_cry_20 ));
    CascadeMux I__5949 (
            .O(N__41004),
            .I(N__41001));
    InMux I__5948 (
            .O(N__41001),
            .I(N__40997));
    InMux I__5947 (
            .O(N__41000),
            .I(N__40994));
    LocalMux I__5946 (
            .O(N__40997),
            .I(N__40991));
    LocalMux I__5945 (
            .O(N__40994),
            .I(\reset_module_System.countZ0Z_21 ));
    Odrv4 I__5944 (
            .O(N__40991),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__5943 (
            .O(N__40986),
            .I(N__40983));
    LocalMux I__5942 (
            .O(N__40983),
            .I(N__40979));
    InMux I__5941 (
            .O(N__40982),
            .I(N__40976));
    Sp12to4 I__5940 (
            .O(N__40979),
            .I(N__40973));
    LocalMux I__5939 (
            .O(N__40976),
            .I(\reset_module_System.countZ0Z_10 ));
    Odrv12 I__5938 (
            .O(N__40973),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__5937 (
            .O(N__40968),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__5936 (
            .O(N__40965),
            .I(N__40962));
    LocalMux I__5935 (
            .O(N__40962),
            .I(N__40958));
    InMux I__5934 (
            .O(N__40961),
            .I(N__40955));
    Span4Mux_v I__5933 (
            .O(N__40958),
            .I(N__40952));
    LocalMux I__5932 (
            .O(N__40955),
            .I(\reset_module_System.countZ0Z_11 ));
    Odrv4 I__5931 (
            .O(N__40952),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__5930 (
            .O(N__40947),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__5929 (
            .O(N__40944),
            .I(N__40940));
    InMux I__5928 (
            .O(N__40943),
            .I(N__40937));
    LocalMux I__5927 (
            .O(N__40940),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__5926 (
            .O(N__40937),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__5925 (
            .O(N__40932),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__5924 (
            .O(N__40929),
            .I(N__40926));
    LocalMux I__5923 (
            .O(N__40926),
            .I(N__40922));
    InMux I__5922 (
            .O(N__40925),
            .I(N__40919));
    Odrv4 I__5921 (
            .O(N__40922),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__5920 (
            .O(N__40919),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__5919 (
            .O(N__40914),
            .I(\reset_module_System.count_1_cry_12 ));
    CascadeMux I__5918 (
            .O(N__40911),
            .I(N__40907));
    InMux I__5917 (
            .O(N__40910),
            .I(N__40904));
    InMux I__5916 (
            .O(N__40907),
            .I(N__40901));
    LocalMux I__5915 (
            .O(N__40904),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__5914 (
            .O(N__40901),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__5913 (
            .O(N__40896),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__5912 (
            .O(N__40893),
            .I(N__40890));
    LocalMux I__5911 (
            .O(N__40890),
            .I(N__40886));
    InMux I__5910 (
            .O(N__40889),
            .I(N__40883));
    Odrv4 I__5909 (
            .O(N__40886),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__5908 (
            .O(N__40883),
            .I(\reset_module_System.countZ0Z_15 ));
    InMux I__5907 (
            .O(N__40878),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__5906 (
            .O(N__40875),
            .I(N__40872));
    LocalMux I__5905 (
            .O(N__40872),
            .I(N__40868));
    InMux I__5904 (
            .O(N__40871),
            .I(N__40865));
    Odrv4 I__5903 (
            .O(N__40868),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__5902 (
            .O(N__40865),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__5901 (
            .O(N__40860),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__5900 (
            .O(N__40857),
            .I(N__40853));
    InMux I__5899 (
            .O(N__40856),
            .I(N__40850));
    LocalMux I__5898 (
            .O(N__40853),
            .I(N__40847));
    LocalMux I__5897 (
            .O(N__40850),
            .I(\reset_module_System.countZ0Z_17 ));
    Odrv4 I__5896 (
            .O(N__40847),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__5895 (
            .O(N__40842),
            .I(bfn_9_10_0_));
    InMux I__5894 (
            .O(N__40839),
            .I(N__40835));
    InMux I__5893 (
            .O(N__40838),
            .I(N__40832));
    LocalMux I__5892 (
            .O(N__40835),
            .I(N__40828));
    LocalMux I__5891 (
            .O(N__40832),
            .I(N__40825));
    InMux I__5890 (
            .O(N__40831),
            .I(N__40822));
    Span4Mux_h I__5889 (
            .O(N__40828),
            .I(N__40819));
    Odrv4 I__5888 (
            .O(N__40825),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__5887 (
            .O(N__40822),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__5886 (
            .O(N__40819),
            .I(\reset_module_System.countZ0Z_1 ));
    CascadeMux I__5885 (
            .O(N__40812),
            .I(N__40806));
    InMux I__5884 (
            .O(N__40811),
            .I(N__40803));
    InMux I__5883 (
            .O(N__40810),
            .I(N__40798));
    InMux I__5882 (
            .O(N__40809),
            .I(N__40798));
    InMux I__5881 (
            .O(N__40806),
            .I(N__40795));
    LocalMux I__5880 (
            .O(N__40803),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5879 (
            .O(N__40798),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5878 (
            .O(N__40795),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__5877 (
            .O(N__40788),
            .I(N__40784));
    InMux I__5876 (
            .O(N__40787),
            .I(N__40781));
    LocalMux I__5875 (
            .O(N__40784),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__5874 (
            .O(N__40781),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__5873 (
            .O(N__40776),
            .I(N__40773));
    LocalMux I__5872 (
            .O(N__40773),
            .I(\reset_module_System.count_1_2 ));
    InMux I__5871 (
            .O(N__40770),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__5870 (
            .O(N__40767),
            .I(N__40763));
    InMux I__5869 (
            .O(N__40766),
            .I(N__40760));
    LocalMux I__5868 (
            .O(N__40763),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__5867 (
            .O(N__40760),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__5866 (
            .O(N__40755),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__5865 (
            .O(N__40752),
            .I(N__40748));
    InMux I__5864 (
            .O(N__40751),
            .I(N__40745));
    LocalMux I__5863 (
            .O(N__40748),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__5862 (
            .O(N__40745),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__5861 (
            .O(N__40740),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__5860 (
            .O(N__40737),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__5859 (
            .O(N__40734),
            .I(N__40730));
    InMux I__5858 (
            .O(N__40733),
            .I(N__40727));
    LocalMux I__5857 (
            .O(N__40730),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__5856 (
            .O(N__40727),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__5855 (
            .O(N__40722),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__5854 (
            .O(N__40719),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__5853 (
            .O(N__40716),
            .I(\reset_module_System.count_1_cry_7 ));
    InMux I__5852 (
            .O(N__40713),
            .I(bfn_9_9_0_));
    InMux I__5851 (
            .O(N__40710),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__5850 (
            .O(N__40707),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    SRMux I__5849 (
            .O(N__40704),
            .I(N__40700));
    SRMux I__5848 (
            .O(N__40703),
            .I(N__40697));
    LocalMux I__5847 (
            .O(N__40700),
            .I(N__40694));
    LocalMux I__5846 (
            .O(N__40697),
            .I(N__40691));
    Odrv4 I__5845 (
            .O(N__40694),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    Odrv4 I__5844 (
            .O(N__40691),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    InMux I__5843 (
            .O(N__40686),
            .I(N__40683));
    LocalMux I__5842 (
            .O(N__40683),
            .I(N__40680));
    Odrv4 I__5841 (
            .O(N__40680),
            .I(\reset_module_System.count_1_1 ));
    CascadeMux I__5840 (
            .O(N__40677),
            .I(N__40673));
    InMux I__5839 (
            .O(N__40676),
            .I(N__40668));
    InMux I__5838 (
            .O(N__40673),
            .I(N__40665));
    InMux I__5837 (
            .O(N__40672),
            .I(N__40660));
    InMux I__5836 (
            .O(N__40671),
            .I(N__40660));
    LocalMux I__5835 (
            .O(N__40668),
            .I(N__40657));
    LocalMux I__5834 (
            .O(N__40665),
            .I(N__40654));
    LocalMux I__5833 (
            .O(N__40660),
            .I(N__40651));
    Span4Mux_s2_v I__5832 (
            .O(N__40657),
            .I(N__40648));
    Span4Mux_h I__5831 (
            .O(N__40654),
            .I(N__40641));
    Span4Mux_v I__5830 (
            .O(N__40651),
            .I(N__40641));
    Span4Mux_v I__5829 (
            .O(N__40648),
            .I(N__40641));
    Odrv4 I__5828 (
            .O(N__40641),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__5827 (
            .O(N__40638),
            .I(N__40633));
    InMux I__5826 (
            .O(N__40637),
            .I(N__40630));
    InMux I__5825 (
            .O(N__40636),
            .I(N__40625));
    InMux I__5824 (
            .O(N__40633),
            .I(N__40625));
    LocalMux I__5823 (
            .O(N__40630),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__5822 (
            .O(N__40625),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    CascadeMux I__5821 (
            .O(N__40620),
            .I(\uart_drone.N_126_li_cascade_ ));
    CascadeMux I__5820 (
            .O(N__40617),
            .I(\uart_drone.N_143_cascade_ ));
    InMux I__5819 (
            .O(N__40614),
            .I(N__40611));
    LocalMux I__5818 (
            .O(N__40611),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__5817 (
            .O(N__40608),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__5816 (
            .O(N__40605),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__5815 (
            .O(N__40602),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__5814 (
            .O(N__40599),
            .I(bfn_9_6_0_));
    InMux I__5813 (
            .O(N__40596),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__5812 (
            .O(N__40593),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__5811 (
            .O(N__40590),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__5810 (
            .O(N__40587),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__5809 (
            .O(N__40584),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__5808 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__5807 (
            .O(N__40578),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__5806 (
            .O(N__40575),
            .I(N__40572));
    LocalMux I__5805 (
            .O(N__40572),
            .I(N__40569));
    Odrv4 I__5804 (
            .O(N__40569),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    InMux I__5803 (
            .O(N__40566),
            .I(N__40563));
    LocalMux I__5802 (
            .O(N__40563),
            .I(N__40560));
    Span4Mux_h I__5801 (
            .O(N__40560),
            .I(N__40557));
    Odrv4 I__5800 (
            .O(N__40557),
            .I(uart_input_drone_c));
    InMux I__5799 (
            .O(N__40554),
            .I(N__40551));
    LocalMux I__5798 (
            .O(N__40551),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__5797 (
            .O(N__40548),
            .I(N__40545));
    LocalMux I__5796 (
            .O(N__40545),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__5795 (
            .O(N__40542),
            .I(N__40539));
    LocalMux I__5794 (
            .O(N__40539),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__5793 (
            .O(N__40536),
            .I(N__40533));
    LocalMux I__5792 (
            .O(N__40533),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__5791 (
            .O(N__40530),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__5790 (
            .O(N__40527),
            .I(N__40524));
    LocalMux I__5789 (
            .O(N__40524),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__5788 (
            .O(N__40521),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__5787 (
            .O(N__40518),
            .I(N__40515));
    LocalMux I__5786 (
            .O(N__40515),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__5785 (
            .O(N__40512),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__5784 (
            .O(N__40509),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    CascadeMux I__5783 (
            .O(N__40506),
            .I(N__40502));
    InMux I__5782 (
            .O(N__40505),
            .I(N__40499));
    InMux I__5781 (
            .O(N__40502),
            .I(N__40496));
    LocalMux I__5780 (
            .O(N__40499),
            .I(\pid_front.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__5779 (
            .O(N__40496),
            .I(\pid_front.error_i_acumm_preregZ0Z_14 ));
    InMux I__5778 (
            .O(N__40491),
            .I(N__40488));
    LocalMux I__5777 (
            .O(N__40488),
            .I(N__40484));
    InMux I__5776 (
            .O(N__40487),
            .I(N__40481));
    Odrv4 I__5775 (
            .O(N__40484),
            .I(\pid_front.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__5774 (
            .O(N__40481),
            .I(\pid_front.error_i_acumm_preregZ0Z_20 ));
    InMux I__5773 (
            .O(N__40476),
            .I(N__40472));
    InMux I__5772 (
            .O(N__40475),
            .I(N__40469));
    LocalMux I__5771 (
            .O(N__40472),
            .I(\pid_front.error_i_acumm_preregZ0Z_15 ));
    LocalMux I__5770 (
            .O(N__40469),
            .I(\pid_front.error_i_acumm_preregZ0Z_15 ));
    InMux I__5769 (
            .O(N__40464),
            .I(N__40460));
    InMux I__5768 (
            .O(N__40463),
            .I(N__40457));
    LocalMux I__5767 (
            .O(N__40460),
            .I(drone_H_disp_side_3));
    LocalMux I__5766 (
            .O(N__40457),
            .I(drone_H_disp_side_3));
    CEMux I__5765 (
            .O(N__40452),
            .I(N__40449));
    LocalMux I__5764 (
            .O(N__40449),
            .I(N__40445));
    CEMux I__5763 (
            .O(N__40448),
            .I(N__40442));
    Span4Mux_v I__5762 (
            .O(N__40445),
            .I(N__40439));
    LocalMux I__5761 (
            .O(N__40442),
            .I(N__40436));
    Odrv4 I__5760 (
            .O(N__40439),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    Odrv4 I__5759 (
            .O(N__40436),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__5758 (
            .O(N__40431),
            .I(N__40428));
    LocalMux I__5757 (
            .O(N__40428),
            .I(N__40425));
    Odrv12 I__5756 (
            .O(N__40425),
            .I(uart_input_pc_c));
    InMux I__5755 (
            .O(N__40422),
            .I(N__40419));
    LocalMux I__5754 (
            .O(N__40419),
            .I(N__40416));
    Odrv4 I__5753 (
            .O(N__40416),
            .I(\pid_front.error_i_acumm16lto27_10 ));
    CascadeMux I__5752 (
            .O(N__40413),
            .I(\pid_front.un10lto27_8_cascade_ ));
    InMux I__5751 (
            .O(N__40410),
            .I(N__40404));
    InMux I__5750 (
            .O(N__40409),
            .I(N__40404));
    LocalMux I__5749 (
            .O(N__40404),
            .I(\pid_front.error_i_acumm_preregZ0Z_26 ));
    CascadeMux I__5748 (
            .O(N__40401),
            .I(\pid_front.un10lto27_9_cascade_ ));
    InMux I__5747 (
            .O(N__40398),
            .I(N__40395));
    LocalMux I__5746 (
            .O(N__40395),
            .I(\pid_front.un10lto27_11 ));
    InMux I__5745 (
            .O(N__40392),
            .I(N__40389));
    LocalMux I__5744 (
            .O(N__40389),
            .I(\pid_front.un10lto27_10 ));
    InMux I__5743 (
            .O(N__40386),
            .I(N__40382));
    InMux I__5742 (
            .O(N__40385),
            .I(N__40379));
    LocalMux I__5741 (
            .O(N__40382),
            .I(\pid_front.error_i_acumm_preregZ0Z_18 ));
    LocalMux I__5740 (
            .O(N__40379),
            .I(\pid_front.error_i_acumm_preregZ0Z_18 ));
    InMux I__5739 (
            .O(N__40374),
            .I(N__40370));
    InMux I__5738 (
            .O(N__40373),
            .I(N__40367));
    LocalMux I__5737 (
            .O(N__40370),
            .I(\pid_front.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__5736 (
            .O(N__40367),
            .I(\pid_front.error_i_acumm_preregZ0Z_19 ));
    InMux I__5735 (
            .O(N__40362),
            .I(N__40359));
    LocalMux I__5734 (
            .O(N__40359),
            .I(N__40356));
    Odrv4 I__5733 (
            .O(N__40356),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ));
    CascadeMux I__5732 (
            .O(N__40353),
            .I(\pid_front.error_i_acumm16lt9_0_cascade_ ));
    InMux I__5731 (
            .O(N__40350),
            .I(N__40347));
    LocalMux I__5730 (
            .O(N__40347),
            .I(\pid_front.un10lt9_1 ));
    CascadeMux I__5729 (
            .O(N__40344),
            .I(\pid_front.un10lt9_cascade_ ));
    InMux I__5728 (
            .O(N__40341),
            .I(N__40338));
    LocalMux I__5727 (
            .O(N__40338),
            .I(\pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ));
    CascadeMux I__5726 (
            .O(N__40335),
            .I(\pid_front.error_i_acumm16lto27_7_cascade_ ));
    InMux I__5725 (
            .O(N__40332),
            .I(N__40329));
    LocalMux I__5724 (
            .O(N__40329),
            .I(\pid_front.error_i_acumm16lto27_8 ));
    InMux I__5723 (
            .O(N__40326),
            .I(N__40323));
    LocalMux I__5722 (
            .O(N__40323),
            .I(\pid_front.error_i_acumm16lto27_9 ));
    InMux I__5721 (
            .O(N__40320),
            .I(N__40314));
    InMux I__5720 (
            .O(N__40319),
            .I(N__40309));
    InMux I__5719 (
            .O(N__40318),
            .I(N__40309));
    InMux I__5718 (
            .O(N__40317),
            .I(N__40306));
    LocalMux I__5717 (
            .O(N__40314),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    LocalMux I__5716 (
            .O(N__40309),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    LocalMux I__5715 (
            .O(N__40306),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    InMux I__5714 (
            .O(N__40299),
            .I(N__40293));
    InMux I__5713 (
            .O(N__40298),
            .I(N__40293));
    LocalMux I__5712 (
            .O(N__40293),
            .I(N__40287));
    InMux I__5711 (
            .O(N__40292),
            .I(N__40280));
    InMux I__5710 (
            .O(N__40291),
            .I(N__40280));
    InMux I__5709 (
            .O(N__40290),
            .I(N__40280));
    Odrv4 I__5708 (
            .O(N__40287),
            .I(\pid_front.error_d_regZ0Z_5 ));
    LocalMux I__5707 (
            .O(N__40280),
            .I(\pid_front.error_d_regZ0Z_5 ));
    CascadeMux I__5706 (
            .O(N__40275),
            .I(N__40271));
    InMux I__5705 (
            .O(N__40274),
            .I(N__40266));
    InMux I__5704 (
            .O(N__40271),
            .I(N__40266));
    LocalMux I__5703 (
            .O(N__40266),
            .I(N__40263));
    Span4Mux_h I__5702 (
            .O(N__40263),
            .I(N__40260));
    Span4Mux_h I__5701 (
            .O(N__40260),
            .I(N__40257));
    Odrv4 I__5700 (
            .O(N__40257),
            .I(\pid_front.error_p_regZ0Z_5 ));
    InMux I__5699 (
            .O(N__40254),
            .I(N__40251));
    LocalMux I__5698 (
            .O(N__40251),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ));
    CascadeMux I__5697 (
            .O(N__40248),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ));
    InMux I__5696 (
            .O(N__40245),
            .I(N__40242));
    LocalMux I__5695 (
            .O(N__40242),
            .I(N__40238));
    InMux I__5694 (
            .O(N__40241),
            .I(N__40235));
    Span4Mux_v I__5693 (
            .O(N__40238),
            .I(N__40230));
    LocalMux I__5692 (
            .O(N__40235),
            .I(N__40230));
    Span4Mux_v I__5691 (
            .O(N__40230),
            .I(N__40227));
    Odrv4 I__5690 (
            .O(N__40227),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__5689 (
            .O(N__40224),
            .I(N__40218));
    InMux I__5688 (
            .O(N__40223),
            .I(N__40215));
    InMux I__5687 (
            .O(N__40222),
            .I(N__40210));
    InMux I__5686 (
            .O(N__40221),
            .I(N__40210));
    LocalMux I__5685 (
            .O(N__40218),
            .I(N__40199));
    LocalMux I__5684 (
            .O(N__40215),
            .I(N__40194));
    LocalMux I__5683 (
            .O(N__40210),
            .I(N__40194));
    InMux I__5682 (
            .O(N__40209),
            .I(N__40179));
    InMux I__5681 (
            .O(N__40208),
            .I(N__40179));
    InMux I__5680 (
            .O(N__40207),
            .I(N__40179));
    InMux I__5679 (
            .O(N__40206),
            .I(N__40179));
    InMux I__5678 (
            .O(N__40205),
            .I(N__40179));
    InMux I__5677 (
            .O(N__40204),
            .I(N__40179));
    InMux I__5676 (
            .O(N__40203),
            .I(N__40179));
    InMux I__5675 (
            .O(N__40202),
            .I(N__40174));
    Span12Mux_v I__5674 (
            .O(N__40199),
            .I(N__40167));
    Sp12to4 I__5673 (
            .O(N__40194),
            .I(N__40167));
    LocalMux I__5672 (
            .O(N__40179),
            .I(N__40167));
    InMux I__5671 (
            .O(N__40178),
            .I(N__40162));
    InMux I__5670 (
            .O(N__40177),
            .I(N__40162));
    LocalMux I__5669 (
            .O(N__40174),
            .I(\Commands_frame_decoder.N_402 ));
    Odrv12 I__5668 (
            .O(N__40167),
            .I(\Commands_frame_decoder.N_402 ));
    LocalMux I__5667 (
            .O(N__40162),
            .I(\Commands_frame_decoder.N_402 ));
    InMux I__5666 (
            .O(N__40155),
            .I(N__40151));
    InMux I__5665 (
            .O(N__40154),
            .I(N__40148));
    LocalMux I__5664 (
            .O(N__40151),
            .I(N__40145));
    LocalMux I__5663 (
            .O(N__40148),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    Odrv12 I__5662 (
            .O(N__40145),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__5661 (
            .O(N__40140),
            .I(N__40136));
    InMux I__5660 (
            .O(N__40139),
            .I(N__40133));
    LocalMux I__5659 (
            .O(N__40136),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    LocalMux I__5658 (
            .O(N__40133),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    CascadeMux I__5657 (
            .O(N__40128),
            .I(\pid_front.un10lt9_1_cascade_ ));
    InMux I__5656 (
            .O(N__40125),
            .I(N__40122));
    LocalMux I__5655 (
            .O(N__40122),
            .I(N__40119));
    Span12Mux_v I__5654 (
            .O(N__40119),
            .I(N__40116));
    Span12Mux_h I__5653 (
            .O(N__40116),
            .I(N__40113));
    Odrv12 I__5652 (
            .O(N__40113),
            .I(\pid_front.O_9 ));
    InMux I__5651 (
            .O(N__40110),
            .I(N__40107));
    LocalMux I__5650 (
            .O(N__40107),
            .I(N__40104));
    Span4Mux_v I__5649 (
            .O(N__40104),
            .I(N__40101));
    Span4Mux_h I__5648 (
            .O(N__40101),
            .I(N__40098));
    Odrv4 I__5647 (
            .O(N__40098),
            .I(\pid_front.O_0_13 ));
    InMux I__5646 (
            .O(N__40095),
            .I(N__40092));
    LocalMux I__5645 (
            .O(N__40092),
            .I(N__40089));
    Span4Mux_h I__5644 (
            .O(N__40089),
            .I(N__40086));
    Span4Mux_h I__5643 (
            .O(N__40086),
            .I(N__40083));
    Odrv4 I__5642 (
            .O(N__40083),
            .I(\pid_front.O_0_14 ));
    InMux I__5641 (
            .O(N__40080),
            .I(N__40077));
    LocalMux I__5640 (
            .O(N__40077),
            .I(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ));
    CascadeMux I__5639 (
            .O(N__40074),
            .I(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ));
    CascadeMux I__5638 (
            .O(N__40071),
            .I(N__40068));
    InMux I__5637 (
            .O(N__40068),
            .I(N__40062));
    InMux I__5636 (
            .O(N__40067),
            .I(N__40062));
    LocalMux I__5635 (
            .O(N__40062),
            .I(N__40059));
    Span4Mux_h I__5634 (
            .O(N__40059),
            .I(N__40056));
    Span4Mux_h I__5633 (
            .O(N__40056),
            .I(N__40053));
    Odrv4 I__5632 (
            .O(N__40053),
            .I(\pid_front.error_p_regZ0Z_4 ));
    InMux I__5631 (
            .O(N__40050),
            .I(N__40044));
    InMux I__5630 (
            .O(N__40049),
            .I(N__40044));
    LocalMux I__5629 (
            .O(N__40044),
            .I(\pid_front.error_d_reg_prevZ0Z_4 ));
    CascadeMux I__5628 (
            .O(N__40041),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ));
    InMux I__5627 (
            .O(N__40038),
            .I(N__40032));
    InMux I__5626 (
            .O(N__40037),
            .I(N__40032));
    LocalMux I__5625 (
            .O(N__40032),
            .I(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ));
    CascadeMux I__5624 (
            .O(N__40029),
            .I(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8_cascade_ ));
    InMux I__5623 (
            .O(N__40026),
            .I(N__40023));
    LocalMux I__5622 (
            .O(N__40023),
            .I(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ));
    InMux I__5621 (
            .O(N__40020),
            .I(N__40017));
    LocalMux I__5620 (
            .O(N__40017),
            .I(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ));
    CascadeMux I__5619 (
            .O(N__40014),
            .I(N__40011));
    InMux I__5618 (
            .O(N__40011),
            .I(N__40005));
    InMux I__5617 (
            .O(N__40010),
            .I(N__40005));
    LocalMux I__5616 (
            .O(N__40005),
            .I(N__40002));
    Odrv4 I__5615 (
            .O(N__40002),
            .I(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ));
    CascadeMux I__5614 (
            .O(N__39999),
            .I(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ));
    InMux I__5613 (
            .O(N__39996),
            .I(N__39993));
    LocalMux I__5612 (
            .O(N__39993),
            .I(\pid_front.N_1668_i ));
    InMux I__5611 (
            .O(N__39990),
            .I(N__39984));
    InMux I__5610 (
            .O(N__39989),
            .I(N__39984));
    LocalMux I__5609 (
            .O(N__39984),
            .I(N__39981));
    Span4Mux_v I__5608 (
            .O(N__39981),
            .I(N__39978));
    Span4Mux_h I__5607 (
            .O(N__39978),
            .I(N__39975));
    Odrv4 I__5606 (
            .O(N__39975),
            .I(\pid_front.error_p_regZ0Z_7 ));
    CascadeMux I__5605 (
            .O(N__39972),
            .I(N__39969));
    InMux I__5604 (
            .O(N__39969),
            .I(N__39963));
    InMux I__5603 (
            .O(N__39968),
            .I(N__39963));
    LocalMux I__5602 (
            .O(N__39963),
            .I(N__39959));
    InMux I__5601 (
            .O(N__39962),
            .I(N__39956));
    Odrv4 I__5600 (
            .O(N__39959),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    LocalMux I__5599 (
            .O(N__39956),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    CascadeMux I__5598 (
            .O(N__39951),
            .I(\pid_front.N_1668_i_cascade_ ));
    InMux I__5597 (
            .O(N__39948),
            .I(N__39942));
    InMux I__5596 (
            .O(N__39947),
            .I(N__39942));
    LocalMux I__5595 (
            .O(N__39942),
            .I(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ));
    InMux I__5594 (
            .O(N__39939),
            .I(N__39936));
    LocalMux I__5593 (
            .O(N__39936),
            .I(N__39933));
    Span4Mux_v I__5592 (
            .O(N__39933),
            .I(N__39930));
    Span4Mux_h I__5591 (
            .O(N__39930),
            .I(N__39927));
    Span4Mux_h I__5590 (
            .O(N__39927),
            .I(N__39924));
    Span4Mux_h I__5589 (
            .O(N__39924),
            .I(N__39921));
    Span4Mux_h I__5588 (
            .O(N__39921),
            .I(N__39918));
    Odrv4 I__5587 (
            .O(N__39918),
            .I(\pid_front.O_7 ));
    InMux I__5586 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__5585 (
            .O(N__39912),
            .I(N__39909));
    Sp12to4 I__5584 (
            .O(N__39909),
            .I(N__39906));
    Span12Mux_v I__5583 (
            .O(N__39906),
            .I(N__39903));
    Span12Mux_h I__5582 (
            .O(N__39903),
            .I(N__39900));
    Odrv12 I__5581 (
            .O(N__39900),
            .I(\pid_front.O_8 ));
    InMux I__5580 (
            .O(N__39897),
            .I(N__39889));
    InMux I__5579 (
            .O(N__39896),
            .I(N__39889));
    InMux I__5578 (
            .O(N__39895),
            .I(N__39884));
    InMux I__5577 (
            .O(N__39894),
            .I(N__39884));
    LocalMux I__5576 (
            .O(N__39889),
            .I(\pid_front.error_d_regZ0Z_6 ));
    LocalMux I__5575 (
            .O(N__39884),
            .I(\pid_front.error_d_regZ0Z_6 ));
    InMux I__5574 (
            .O(N__39879),
            .I(N__39876));
    LocalMux I__5573 (
            .O(N__39876),
            .I(N__39873));
    Span4Mux_v I__5572 (
            .O(N__39873),
            .I(N__39870));
    Span4Mux_h I__5571 (
            .O(N__39870),
            .I(N__39867));
    Odrv4 I__5570 (
            .O(N__39867),
            .I(\dron_frame_decoder_1.state_ns_i_i_a2_1_0 ));
    CascadeMux I__5569 (
            .O(N__39864),
            .I(\dron_frame_decoder_1.N_186_cascade_ ));
    InMux I__5568 (
            .O(N__39861),
            .I(N__39857));
    InMux I__5567 (
            .O(N__39860),
            .I(N__39854));
    LocalMux I__5566 (
            .O(N__39857),
            .I(\dron_frame_decoder_1.N_127_mux ));
    LocalMux I__5565 (
            .O(N__39854),
            .I(\dron_frame_decoder_1.N_127_mux ));
    InMux I__5564 (
            .O(N__39849),
            .I(N__39846));
    LocalMux I__5563 (
            .O(N__39846),
            .I(\dron_frame_decoder_1.state_ns_i_i_0_0 ));
    InMux I__5562 (
            .O(N__39843),
            .I(N__39840));
    LocalMux I__5561 (
            .O(N__39840),
            .I(N__39837));
    Odrv12 I__5560 (
            .O(N__39837),
            .I(\reset_module_System.reset6_3 ));
    InMux I__5559 (
            .O(N__39834),
            .I(N__39831));
    LocalMux I__5558 (
            .O(N__39831),
            .I(\dron_frame_decoder_1.drone_H_disp_front_9 ));
    InMux I__5557 (
            .O(N__39828),
            .I(N__39825));
    LocalMux I__5556 (
            .O(N__39825),
            .I(N__39822));
    Span4Mux_v I__5555 (
            .O(N__39822),
            .I(N__39819));
    Span4Mux_h I__5554 (
            .O(N__39819),
            .I(N__39816));
    Span4Mux_v I__5553 (
            .O(N__39816),
            .I(N__39813));
    Odrv4 I__5552 (
            .O(N__39813),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    CascadeMux I__5551 (
            .O(N__39810),
            .I(N__39807));
    InMux I__5550 (
            .O(N__39807),
            .I(N__39803));
    InMux I__5549 (
            .O(N__39806),
            .I(N__39800));
    LocalMux I__5548 (
            .O(N__39803),
            .I(N__39795));
    LocalMux I__5547 (
            .O(N__39800),
            .I(N__39795));
    Span4Mux_h I__5546 (
            .O(N__39795),
            .I(N__39792));
    Span4Mux_v I__5545 (
            .O(N__39792),
            .I(N__39789));
    Odrv4 I__5544 (
            .O(N__39789),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    CascadeMux I__5543 (
            .O(N__39786),
            .I(\dron_frame_decoder_1.WDT10_0_icf1_1_cascade_ ));
    InMux I__5542 (
            .O(N__39783),
            .I(N__39780));
    LocalMux I__5541 (
            .O(N__39780),
            .I(\dron_frame_decoder_1.WDT10_0_icf1 ));
    CascadeMux I__5540 (
            .O(N__39777),
            .I(\dron_frame_decoder_1.WDT10lto9_3_cascade_ ));
    InMux I__5539 (
            .O(N__39774),
            .I(N__39768));
    InMux I__5538 (
            .O(N__39773),
            .I(N__39768));
    LocalMux I__5537 (
            .O(N__39768),
            .I(\dron_frame_decoder_1.WDT10lt10 ));
    InMux I__5536 (
            .O(N__39765),
            .I(N__39762));
    LocalMux I__5535 (
            .O(N__39762),
            .I(\dron_frame_decoder_1.m34Z0Z_2 ));
    InMux I__5534 (
            .O(N__39759),
            .I(N__39756));
    LocalMux I__5533 (
            .O(N__39756),
            .I(\dron_frame_decoder_1.N_123_mux ));
    InMux I__5532 (
            .O(N__39753),
            .I(N__39748));
    InMux I__5531 (
            .O(N__39752),
            .I(N__39745));
    InMux I__5530 (
            .O(N__39751),
            .I(N__39742));
    LocalMux I__5529 (
            .O(N__39748),
            .I(N__39739));
    LocalMux I__5528 (
            .O(N__39745),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__5527 (
            .O(N__39742),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    Odrv12 I__5526 (
            .O(N__39739),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    CascadeMux I__5525 (
            .O(N__39732),
            .I(\dron_frame_decoder_1.N_123_mux_cascade_ ));
    InMux I__5524 (
            .O(N__39729),
            .I(N__39726));
    LocalMux I__5523 (
            .O(N__39726),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_3Z0Z_1 ));
    CascadeMux I__5522 (
            .O(N__39723),
            .I(N__39719));
    InMux I__5521 (
            .O(N__39722),
            .I(N__39713));
    InMux I__5520 (
            .O(N__39719),
            .I(N__39713));
    InMux I__5519 (
            .O(N__39718),
            .I(N__39710));
    LocalMux I__5518 (
            .O(N__39713),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    LocalMux I__5517 (
            .O(N__39710),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    InMux I__5516 (
            .O(N__39705),
            .I(N__39698));
    InMux I__5515 (
            .O(N__39704),
            .I(N__39698));
    InMux I__5514 (
            .O(N__39703),
            .I(N__39695));
    LocalMux I__5513 (
            .O(N__39698),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    LocalMux I__5512 (
            .O(N__39695),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    CascadeMux I__5511 (
            .O(N__39690),
            .I(N__39686));
    InMux I__5510 (
            .O(N__39689),
            .I(N__39681));
    InMux I__5509 (
            .O(N__39686),
            .I(N__39681));
    LocalMux I__5508 (
            .O(N__39681),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    InMux I__5507 (
            .O(N__39678),
            .I(N__39675));
    LocalMux I__5506 (
            .O(N__39675),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    CascadeMux I__5505 (
            .O(N__39672),
            .I(N__39669));
    InMux I__5504 (
            .O(N__39669),
            .I(N__39666));
    LocalMux I__5503 (
            .O(N__39666),
            .I(N__39662));
    CascadeMux I__5502 (
            .O(N__39665),
            .I(N__39658));
    Span4Mux_h I__5501 (
            .O(N__39662),
            .I(N__39655));
    InMux I__5500 (
            .O(N__39661),
            .I(N__39651));
    InMux I__5499 (
            .O(N__39658),
            .I(N__39648));
    Span4Mux_v I__5498 (
            .O(N__39655),
            .I(N__39645));
    InMux I__5497 (
            .O(N__39654),
            .I(N__39642));
    LocalMux I__5496 (
            .O(N__39651),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__5495 (
            .O(N__39648),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv4 I__5494 (
            .O(N__39645),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__5493 (
            .O(N__39642),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__5492 (
            .O(N__39633),
            .I(N__39630));
    LocalMux I__5491 (
            .O(N__39630),
            .I(N__39627));
    Odrv4 I__5490 (
            .O(N__39627),
            .I(\dron_frame_decoder_1.WDT10lt13 ));
    CascadeMux I__5489 (
            .O(N__39624),
            .I(\dron_frame_decoder_1.WDT10_0_icf0_1_cascade_ ));
    CascadeMux I__5488 (
            .O(N__39621),
            .I(\dron_frame_decoder_1.WDT10_0_icf0_cascade_ ));
    InMux I__5487 (
            .O(N__39618),
            .I(N__39615));
    LocalMux I__5486 (
            .O(N__39615),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    CascadeMux I__5485 (
            .O(N__39612),
            .I(N__39609));
    InMux I__5484 (
            .O(N__39609),
            .I(N__39605));
    CascadeMux I__5483 (
            .O(N__39608),
            .I(N__39602));
    LocalMux I__5482 (
            .O(N__39605),
            .I(N__39599));
    InMux I__5481 (
            .O(N__39602),
            .I(N__39596));
    Odrv4 I__5480 (
            .O(N__39599),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__5479 (
            .O(N__39596),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__5478 (
            .O(N__39591),
            .I(N__39580));
    InMux I__5477 (
            .O(N__39590),
            .I(N__39577));
    InMux I__5476 (
            .O(N__39589),
            .I(N__39572));
    InMux I__5475 (
            .O(N__39588),
            .I(N__39572));
    InMux I__5474 (
            .O(N__39587),
            .I(N__39569));
    InMux I__5473 (
            .O(N__39586),
            .I(N__39562));
    InMux I__5472 (
            .O(N__39585),
            .I(N__39562));
    InMux I__5471 (
            .O(N__39584),
            .I(N__39562));
    InMux I__5470 (
            .O(N__39583),
            .I(N__39559));
    LocalMux I__5469 (
            .O(N__39580),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5468 (
            .O(N__39577),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5467 (
            .O(N__39572),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5466 (
            .O(N__39569),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5465 (
            .O(N__39562),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5464 (
            .O(N__39559),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    CascadeMux I__5463 (
            .O(N__39546),
            .I(N__39539));
    CascadeMux I__5462 (
            .O(N__39545),
            .I(N__39534));
    CascadeMux I__5461 (
            .O(N__39544),
            .I(N__39530));
    InMux I__5460 (
            .O(N__39543),
            .I(N__39523));
    InMux I__5459 (
            .O(N__39542),
            .I(N__39523));
    InMux I__5458 (
            .O(N__39539),
            .I(N__39518));
    InMux I__5457 (
            .O(N__39538),
            .I(N__39518));
    InMux I__5456 (
            .O(N__39537),
            .I(N__39507));
    InMux I__5455 (
            .O(N__39534),
            .I(N__39507));
    InMux I__5454 (
            .O(N__39533),
            .I(N__39507));
    InMux I__5453 (
            .O(N__39530),
            .I(N__39507));
    InMux I__5452 (
            .O(N__39529),
            .I(N__39507));
    InMux I__5451 (
            .O(N__39528),
            .I(N__39504));
    LocalMux I__5450 (
            .O(N__39523),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5449 (
            .O(N__39518),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5448 (
            .O(N__39507),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5447 (
            .O(N__39504),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__5446 (
            .O(N__39495),
            .I(N__39480));
    InMux I__5445 (
            .O(N__39494),
            .I(N__39480));
    InMux I__5444 (
            .O(N__39493),
            .I(N__39475));
    InMux I__5443 (
            .O(N__39492),
            .I(N__39475));
    InMux I__5442 (
            .O(N__39491),
            .I(N__39462));
    InMux I__5441 (
            .O(N__39490),
            .I(N__39462));
    InMux I__5440 (
            .O(N__39489),
            .I(N__39462));
    InMux I__5439 (
            .O(N__39488),
            .I(N__39462));
    InMux I__5438 (
            .O(N__39487),
            .I(N__39462));
    InMux I__5437 (
            .O(N__39486),
            .I(N__39462));
    InMux I__5436 (
            .O(N__39485),
            .I(N__39459));
    LocalMux I__5435 (
            .O(N__39480),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5434 (
            .O(N__39475),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5433 (
            .O(N__39462),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5432 (
            .O(N__39459),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CascadeMux I__5431 (
            .O(N__39450),
            .I(N__39447));
    InMux I__5430 (
            .O(N__39447),
            .I(N__39444));
    LocalMux I__5429 (
            .O(N__39444),
            .I(\uart_pc.data_Auxce_0_6 ));
    CascadeMux I__5428 (
            .O(N__39441),
            .I(N__39438));
    InMux I__5427 (
            .O(N__39438),
            .I(N__39435));
    LocalMux I__5426 (
            .O(N__39435),
            .I(N__39431));
    InMux I__5425 (
            .O(N__39434),
            .I(N__39428));
    Odrv4 I__5424 (
            .O(N__39431),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__5423 (
            .O(N__39428),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    CascadeMux I__5422 (
            .O(N__39423),
            .I(N__39416));
    CascadeMux I__5421 (
            .O(N__39422),
            .I(N__39413));
    CascadeMux I__5420 (
            .O(N__39421),
            .I(N__39410));
    IoInMux I__5419 (
            .O(N__39420),
            .I(N__39402));
    InMux I__5418 (
            .O(N__39419),
            .I(N__39396));
    InMux I__5417 (
            .O(N__39416),
            .I(N__39396));
    InMux I__5416 (
            .O(N__39413),
            .I(N__39387));
    InMux I__5415 (
            .O(N__39410),
            .I(N__39387));
    InMux I__5414 (
            .O(N__39409),
            .I(N__39387));
    InMux I__5413 (
            .O(N__39408),
            .I(N__39387));
    InMux I__5412 (
            .O(N__39407),
            .I(N__39382));
    InMux I__5411 (
            .O(N__39406),
            .I(N__39382));
    InMux I__5410 (
            .O(N__39405),
            .I(N__39379));
    LocalMux I__5409 (
            .O(N__39402),
            .I(N__39373));
    InMux I__5408 (
            .O(N__39401),
            .I(N__39370));
    LocalMux I__5407 (
            .O(N__39396),
            .I(N__39367));
    LocalMux I__5406 (
            .O(N__39387),
            .I(N__39362));
    LocalMux I__5405 (
            .O(N__39382),
            .I(N__39362));
    LocalMux I__5404 (
            .O(N__39379),
            .I(N__39359));
    InMux I__5403 (
            .O(N__39378),
            .I(N__39352));
    InMux I__5402 (
            .O(N__39377),
            .I(N__39352));
    InMux I__5401 (
            .O(N__39376),
            .I(N__39352));
    Span4Mux_s3_v I__5400 (
            .O(N__39373),
            .I(N__39349));
    LocalMux I__5399 (
            .O(N__39370),
            .I(N__39346));
    Span4Mux_v I__5398 (
            .O(N__39367),
            .I(N__39341));
    Span4Mux_v I__5397 (
            .O(N__39362),
            .I(N__39341));
    Span4Mux_v I__5396 (
            .O(N__39359),
            .I(N__39336));
    LocalMux I__5395 (
            .O(N__39352),
            .I(N__39336));
    Sp12to4 I__5394 (
            .O(N__39349),
            .I(N__39333));
    Span4Mux_v I__5393 (
            .O(N__39346),
            .I(N__39328));
    Span4Mux_v I__5392 (
            .O(N__39341),
            .I(N__39328));
    Span4Mux_v I__5391 (
            .O(N__39336),
            .I(N__39325));
    Odrv12 I__5390 (
            .O(N__39333),
            .I(debug_CH2_18A_c));
    Odrv4 I__5389 (
            .O(N__39328),
            .I(debug_CH2_18A_c));
    Odrv4 I__5388 (
            .O(N__39325),
            .I(debug_CH2_18A_c));
    InMux I__5387 (
            .O(N__39318),
            .I(N__39306));
    InMux I__5386 (
            .O(N__39317),
            .I(N__39306));
    InMux I__5385 (
            .O(N__39316),
            .I(N__39293));
    InMux I__5384 (
            .O(N__39315),
            .I(N__39293));
    InMux I__5383 (
            .O(N__39314),
            .I(N__39293));
    InMux I__5382 (
            .O(N__39313),
            .I(N__39293));
    InMux I__5381 (
            .O(N__39312),
            .I(N__39293));
    InMux I__5380 (
            .O(N__39311),
            .I(N__39293));
    LocalMux I__5379 (
            .O(N__39306),
            .I(N__39288));
    LocalMux I__5378 (
            .O(N__39293),
            .I(N__39288));
    Span4Mux_v I__5377 (
            .O(N__39288),
            .I(N__39285));
    Odrv4 I__5376 (
            .O(N__39285),
            .I(\uart_pc.un1_state_2_0 ));
    InMux I__5375 (
            .O(N__39282),
            .I(N__39277));
    InMux I__5374 (
            .O(N__39281),
            .I(N__39274));
    InMux I__5373 (
            .O(N__39280),
            .I(N__39271));
    LocalMux I__5372 (
            .O(N__39277),
            .I(N__39268));
    LocalMux I__5371 (
            .O(N__39274),
            .I(N__39265));
    LocalMux I__5370 (
            .O(N__39271),
            .I(\uart_pc.N_152 ));
    Odrv4 I__5369 (
            .O(N__39268),
            .I(\uart_pc.N_152 ));
    Odrv4 I__5368 (
            .O(N__39265),
            .I(\uart_pc.N_152 ));
    CascadeMux I__5367 (
            .O(N__39258),
            .I(N__39255));
    InMux I__5366 (
            .O(N__39255),
            .I(N__39251));
    CascadeMux I__5365 (
            .O(N__39254),
            .I(N__39248));
    LocalMux I__5364 (
            .O(N__39251),
            .I(N__39245));
    InMux I__5363 (
            .O(N__39248),
            .I(N__39242));
    Odrv4 I__5362 (
            .O(N__39245),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__5361 (
            .O(N__39242),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    SRMux I__5360 (
            .O(N__39237),
            .I(N__39233));
    SRMux I__5359 (
            .O(N__39236),
            .I(N__39230));
    LocalMux I__5358 (
            .O(N__39233),
            .I(N__39227));
    LocalMux I__5357 (
            .O(N__39230),
            .I(N__39224));
    Odrv12 I__5356 (
            .O(N__39227),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv4 I__5355 (
            .O(N__39224),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__5354 (
            .O(N__39219),
            .I(N__39215));
    InMux I__5353 (
            .O(N__39218),
            .I(N__39212));
    LocalMux I__5352 (
            .O(N__39215),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    LocalMux I__5351 (
            .O(N__39212),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    CascadeMux I__5350 (
            .O(N__39207),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    InMux I__5349 (
            .O(N__39204),
            .I(N__39188));
    InMux I__5348 (
            .O(N__39203),
            .I(N__39188));
    InMux I__5347 (
            .O(N__39202),
            .I(N__39188));
    InMux I__5346 (
            .O(N__39201),
            .I(N__39188));
    InMux I__5345 (
            .O(N__39200),
            .I(N__39181));
    InMux I__5344 (
            .O(N__39199),
            .I(N__39181));
    InMux I__5343 (
            .O(N__39198),
            .I(N__39181));
    InMux I__5342 (
            .O(N__39197),
            .I(N__39178));
    LocalMux I__5341 (
            .O(N__39188),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__5340 (
            .O(N__39181),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__5339 (
            .O(N__39178),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    InMux I__5338 (
            .O(N__39171),
            .I(N__39157));
    InMux I__5337 (
            .O(N__39170),
            .I(N__39157));
    InMux I__5336 (
            .O(N__39169),
            .I(N__39157));
    InMux I__5335 (
            .O(N__39168),
            .I(N__39157));
    InMux I__5334 (
            .O(N__39167),
            .I(N__39152));
    InMux I__5333 (
            .O(N__39166),
            .I(N__39152));
    LocalMux I__5332 (
            .O(N__39157),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__5331 (
            .O(N__39152),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__5330 (
            .O(N__39147),
            .I(N__39144));
    LocalMux I__5329 (
            .O(N__39144),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__5328 (
            .O(N__39141),
            .I(N__39138));
    InMux I__5327 (
            .O(N__39138),
            .I(N__39134));
    InMux I__5326 (
            .O(N__39137),
            .I(N__39131));
    LocalMux I__5325 (
            .O(N__39134),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__5324 (
            .O(N__39131),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    InMux I__5323 (
            .O(N__39126),
            .I(N__39123));
    LocalMux I__5322 (
            .O(N__39123),
            .I(\uart_pc.data_Auxce_0_1 ));
    CascadeMux I__5321 (
            .O(N__39120),
            .I(N__39117));
    InMux I__5320 (
            .O(N__39117),
            .I(N__39114));
    LocalMux I__5319 (
            .O(N__39114),
            .I(N__39110));
    InMux I__5318 (
            .O(N__39113),
            .I(N__39107));
    Odrv4 I__5317 (
            .O(N__39110),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__5316 (
            .O(N__39107),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__5315 (
            .O(N__39102),
            .I(N__39099));
    LocalMux I__5314 (
            .O(N__39099),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    CascadeMux I__5313 (
            .O(N__39096),
            .I(N__39092));
    CascadeMux I__5312 (
            .O(N__39095),
            .I(N__39089));
    InMux I__5311 (
            .O(N__39092),
            .I(N__39086));
    InMux I__5310 (
            .O(N__39089),
            .I(N__39083));
    LocalMux I__5309 (
            .O(N__39086),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__5308 (
            .O(N__39083),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    InMux I__5307 (
            .O(N__39078),
            .I(N__39075));
    LocalMux I__5306 (
            .O(N__39075),
            .I(\uart_pc.data_Auxce_0_3 ));
    InMux I__5305 (
            .O(N__39072),
            .I(N__39068));
    InMux I__5304 (
            .O(N__39071),
            .I(N__39065));
    LocalMux I__5303 (
            .O(N__39068),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__5302 (
            .O(N__39065),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    CascadeMux I__5301 (
            .O(N__39060),
            .I(\uart_pc.data_Auxce_0_5_cascade_ ));
    CascadeMux I__5300 (
            .O(N__39057),
            .I(N__39054));
    InMux I__5299 (
            .O(N__39054),
            .I(N__39050));
    InMux I__5298 (
            .O(N__39053),
            .I(N__39047));
    LocalMux I__5297 (
            .O(N__39050),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__5296 (
            .O(N__39047),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    InMux I__5295 (
            .O(N__39042),
            .I(N__39038));
    InMux I__5294 (
            .O(N__39041),
            .I(N__39034));
    LocalMux I__5293 (
            .O(N__39038),
            .I(N__39031));
    InMux I__5292 (
            .O(N__39037),
            .I(N__39028));
    LocalMux I__5291 (
            .O(N__39034),
            .I(\uart_pc.data_rdyc_1 ));
    Odrv4 I__5290 (
            .O(N__39031),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__5289 (
            .O(N__39028),
            .I(\uart_pc.data_rdyc_1 ));
    CascadeMux I__5288 (
            .O(N__39021),
            .I(\reset_module_System.reset6_17_cascade_ ));
    CascadeMux I__5287 (
            .O(N__39018),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__5286 (
            .O(N__39015),
            .I(N__39011));
    CascadeMux I__5285 (
            .O(N__39014),
            .I(N__39007));
    LocalMux I__5284 (
            .O(N__39011),
            .I(N__39003));
    InMux I__5283 (
            .O(N__39010),
            .I(N__39000));
    InMux I__5282 (
            .O(N__39007),
            .I(N__38997));
    InMux I__5281 (
            .O(N__39006),
            .I(N__38994));
    Span4Mux_s2_v I__5280 (
            .O(N__39003),
            .I(N__38991));
    LocalMux I__5279 (
            .O(N__39000),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5278 (
            .O(N__38997),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5277 (
            .O(N__38994),
            .I(\reset_module_System.reset6_14 ));
    Odrv4 I__5276 (
            .O(N__38991),
            .I(\reset_module_System.reset6_14 ));
    InMux I__5275 (
            .O(N__38982),
            .I(N__38979));
    LocalMux I__5274 (
            .O(N__38979),
            .I(N__38974));
    InMux I__5273 (
            .O(N__38978),
            .I(N__38971));
    InMux I__5272 (
            .O(N__38977),
            .I(N__38968));
    Span4Mux_s3_v I__5271 (
            .O(N__38974),
            .I(N__38965));
    LocalMux I__5270 (
            .O(N__38971),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__5269 (
            .O(N__38968),
            .I(\reset_module_System.reset6_19 ));
    Odrv4 I__5268 (
            .O(N__38965),
            .I(\reset_module_System.reset6_19 ));
    InMux I__5267 (
            .O(N__38958),
            .I(N__38955));
    LocalMux I__5266 (
            .O(N__38955),
            .I(\reset_module_System.reset6_11 ));
    InMux I__5265 (
            .O(N__38952),
            .I(N__38944));
    InMux I__5264 (
            .O(N__38951),
            .I(N__38944));
    InMux I__5263 (
            .O(N__38950),
            .I(N__38941));
    InMux I__5262 (
            .O(N__38949),
            .I(N__38938));
    LocalMux I__5261 (
            .O(N__38944),
            .I(N__38935));
    LocalMux I__5260 (
            .O(N__38941),
            .I(N__38932));
    LocalMux I__5259 (
            .O(N__38938),
            .I(N__38927));
    Span4Mux_v I__5258 (
            .O(N__38935),
            .I(N__38922));
    Span4Mux_v I__5257 (
            .O(N__38932),
            .I(N__38922));
    InMux I__5256 (
            .O(N__38931),
            .I(N__38917));
    InMux I__5255 (
            .O(N__38930),
            .I(N__38917));
    Odrv4 I__5254 (
            .O(N__38927),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv4 I__5253 (
            .O(N__38922),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5252 (
            .O(N__38917),
            .I(\uart_pc.stateZ0Z_4 ));
    InMux I__5251 (
            .O(N__38910),
            .I(N__38907));
    LocalMux I__5250 (
            .O(N__38907),
            .I(N__38898));
    InMux I__5249 (
            .O(N__38906),
            .I(N__38895));
    InMux I__5248 (
            .O(N__38905),
            .I(N__38892));
    InMux I__5247 (
            .O(N__38904),
            .I(N__38889));
    InMux I__5246 (
            .O(N__38903),
            .I(N__38886));
    InMux I__5245 (
            .O(N__38902),
            .I(N__38880));
    InMux I__5244 (
            .O(N__38901),
            .I(N__38880));
    Span4Mux_v I__5243 (
            .O(N__38898),
            .I(N__38875));
    LocalMux I__5242 (
            .O(N__38895),
            .I(N__38875));
    LocalMux I__5241 (
            .O(N__38892),
            .I(N__38868));
    LocalMux I__5240 (
            .O(N__38889),
            .I(N__38868));
    LocalMux I__5239 (
            .O(N__38886),
            .I(N__38868));
    InMux I__5238 (
            .O(N__38885),
            .I(N__38865));
    LocalMux I__5237 (
            .O(N__38880),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__5236 (
            .O(N__38875),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__5235 (
            .O(N__38868),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__5234 (
            .O(N__38865),
            .I(\uart_pc.stateZ0Z_3 ));
    InMux I__5233 (
            .O(N__38856),
            .I(N__38853));
    LocalMux I__5232 (
            .O(N__38853),
            .I(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ));
    InMux I__5231 (
            .O(N__38850),
            .I(N__38847));
    LocalMux I__5230 (
            .O(N__38847),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    InMux I__5229 (
            .O(N__38844),
            .I(N__38840));
    InMux I__5228 (
            .O(N__38843),
            .I(N__38837));
    LocalMux I__5227 (
            .O(N__38840),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__5226 (
            .O(N__38837),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    CascadeMux I__5225 (
            .O(N__38832),
            .I(N__38826));
    InMux I__5224 (
            .O(N__38831),
            .I(N__38821));
    InMux I__5223 (
            .O(N__38830),
            .I(N__38821));
    InMux I__5222 (
            .O(N__38829),
            .I(N__38816));
    InMux I__5221 (
            .O(N__38826),
            .I(N__38816));
    LocalMux I__5220 (
            .O(N__38821),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__5219 (
            .O(N__38816),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    InMux I__5218 (
            .O(N__38811),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__5217 (
            .O(N__38808),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__5216 (
            .O(N__38805),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__5215 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__5214 (
            .O(N__38799),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__5213 (
            .O(N__38796),
            .I(N__38793));
    LocalMux I__5212 (
            .O(N__38793),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    InMux I__5211 (
            .O(N__38790),
            .I(N__38787));
    LocalMux I__5210 (
            .O(N__38787),
            .I(N__38784));
    Span4Mux_v I__5209 (
            .O(N__38784),
            .I(N__38781));
    Span4Mux_h I__5208 (
            .O(N__38781),
            .I(N__38778));
    Odrv4 I__5207 (
            .O(N__38778),
            .I(alt_kp_5));
    CEMux I__5206 (
            .O(N__38775),
            .I(N__38770));
    CEMux I__5205 (
            .O(N__38774),
            .I(N__38767));
    CEMux I__5204 (
            .O(N__38773),
            .I(N__38764));
    LocalMux I__5203 (
            .O(N__38770),
            .I(N__38760));
    LocalMux I__5202 (
            .O(N__38767),
            .I(N__38757));
    LocalMux I__5201 (
            .O(N__38764),
            .I(N__38754));
    CEMux I__5200 (
            .O(N__38763),
            .I(N__38751));
    Span4Mux_v I__5199 (
            .O(N__38760),
            .I(N__38741));
    Span4Mux_v I__5198 (
            .O(N__38757),
            .I(N__38741));
    Span4Mux_s3_h I__5197 (
            .O(N__38754),
            .I(N__38741));
    LocalMux I__5196 (
            .O(N__38751),
            .I(N__38741));
    CEMux I__5195 (
            .O(N__38750),
            .I(N__38738));
    Span4Mux_v I__5194 (
            .O(N__38741),
            .I(N__38735));
    LocalMux I__5193 (
            .O(N__38738),
            .I(N__38732));
    Span4Mux_h I__5192 (
            .O(N__38735),
            .I(N__38729));
    Span4Mux_v I__5191 (
            .O(N__38732),
            .I(N__38726));
    Sp12to4 I__5190 (
            .O(N__38729),
            .I(N__38723));
    Span4Mux_v I__5189 (
            .O(N__38726),
            .I(N__38720));
    Odrv12 I__5188 (
            .O(N__38723),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    Odrv4 I__5187 (
            .O(N__38720),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    InMux I__5186 (
            .O(N__38715),
            .I(N__38709));
    InMux I__5185 (
            .O(N__38714),
            .I(N__38709));
    LocalMux I__5184 (
            .O(N__38709),
            .I(\Commands_frame_decoder.N_364_0 ));
    InMux I__5183 (
            .O(N__38706),
            .I(N__38703));
    LocalMux I__5182 (
            .O(N__38703),
            .I(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4 ));
    CascadeMux I__5181 (
            .O(N__38700),
            .I(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ));
    InMux I__5180 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__5179 (
            .O(N__38694),
            .I(N__38691));
    Odrv4 I__5178 (
            .O(N__38691),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    CascadeMux I__5177 (
            .O(N__38688),
            .I(\Commands_frame_decoder.WDT8lt14_0_cascade_ ));
    InMux I__5176 (
            .O(N__38685),
            .I(N__38682));
    LocalMux I__5175 (
            .O(N__38682),
            .I(N__38679));
    Span4Mux_s3_h I__5174 (
            .O(N__38679),
            .I(N__38676));
    Span4Mux_h I__5173 (
            .O(N__38676),
            .I(N__38673));
    Odrv4 I__5172 (
            .O(N__38673),
            .I(alt_kp_0));
    InMux I__5171 (
            .O(N__38670),
            .I(N__38667));
    LocalMux I__5170 (
            .O(N__38667),
            .I(\pid_front.N_1662_i ));
    CascadeMux I__5169 (
            .O(N__38664),
            .I(N__38661));
    InMux I__5168 (
            .O(N__38661),
            .I(N__38655));
    InMux I__5167 (
            .O(N__38660),
            .I(N__38655));
    LocalMux I__5166 (
            .O(N__38655),
            .I(N__38652));
    Span4Mux_h I__5165 (
            .O(N__38652),
            .I(N__38649));
    Span4Mux_h I__5164 (
            .O(N__38649),
            .I(N__38646));
    Odrv4 I__5163 (
            .O(N__38646),
            .I(\pid_front.error_p_regZ0Z_6 ));
    CascadeMux I__5162 (
            .O(N__38643),
            .I(\pid_front.N_1662_i_cascade_ ));
    CascadeMux I__5161 (
            .O(N__38640),
            .I(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ));
    InMux I__5160 (
            .O(N__38637),
            .I(N__38634));
    LocalMux I__5159 (
            .O(N__38634),
            .I(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ));
    CascadeMux I__5158 (
            .O(N__38631),
            .I(\pid_front.un1_pid_prereg_66_0_cascade_ ));
    CEMux I__5157 (
            .O(N__38628),
            .I(N__38625));
    LocalMux I__5156 (
            .O(N__38625),
            .I(N__38621));
    CEMux I__5155 (
            .O(N__38624),
            .I(N__38618));
    Span4Mux_v I__5154 (
            .O(N__38621),
            .I(N__38615));
    LocalMux I__5153 (
            .O(N__38618),
            .I(N__38612));
    Span4Mux_h I__5152 (
            .O(N__38615),
            .I(N__38609));
    Span4Mux_v I__5151 (
            .O(N__38612),
            .I(N__38606));
    Odrv4 I__5150 (
            .O(N__38609),
            .I(\dron_frame_decoder_1.N_371_0 ));
    Odrv4 I__5149 (
            .O(N__38606),
            .I(\dron_frame_decoder_1.N_371_0 ));
    CascadeMux I__5148 (
            .O(N__38601),
            .I(N__38597));
    CascadeMux I__5147 (
            .O(N__38600),
            .I(N__38594));
    InMux I__5146 (
            .O(N__38597),
            .I(N__38590));
    InMux I__5145 (
            .O(N__38594),
            .I(N__38585));
    InMux I__5144 (
            .O(N__38593),
            .I(N__38585));
    LocalMux I__5143 (
            .O(N__38590),
            .I(N__38582));
    LocalMux I__5142 (
            .O(N__38585),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    Odrv4 I__5141 (
            .O(N__38582),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    InMux I__5140 (
            .O(N__38577),
            .I(N__38574));
    LocalMux I__5139 (
            .O(N__38574),
            .I(N__38571));
    Span4Mux_h I__5138 (
            .O(N__38571),
            .I(N__38568));
    Odrv4 I__5137 (
            .O(N__38568),
            .I(\dron_frame_decoder_1.N_10_0 ));
    InMux I__5136 (
            .O(N__38565),
            .I(N__38562));
    LocalMux I__5135 (
            .O(N__38562),
            .I(N__38559));
    Span4Mux_v I__5134 (
            .O(N__38559),
            .I(N__38554));
    InMux I__5133 (
            .O(N__38558),
            .I(N__38549));
    InMux I__5132 (
            .O(N__38557),
            .I(N__38549));
    Odrv4 I__5131 (
            .O(N__38554),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    LocalMux I__5130 (
            .O(N__38549),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    InMux I__5129 (
            .O(N__38544),
            .I(N__38541));
    LocalMux I__5128 (
            .O(N__38541),
            .I(N__38538));
    Span4Mux_v I__5127 (
            .O(N__38538),
            .I(N__38531));
    InMux I__5126 (
            .O(N__38537),
            .I(N__38522));
    InMux I__5125 (
            .O(N__38536),
            .I(N__38522));
    InMux I__5124 (
            .O(N__38535),
            .I(N__38522));
    InMux I__5123 (
            .O(N__38534),
            .I(N__38522));
    Odrv4 I__5122 (
            .O(N__38531),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    LocalMux I__5121 (
            .O(N__38522),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    InMux I__5120 (
            .O(N__38517),
            .I(N__38514));
    LocalMux I__5119 (
            .O(N__38514),
            .I(N__38510));
    CascadeMux I__5118 (
            .O(N__38513),
            .I(N__38507));
    Span4Mux_h I__5117 (
            .O(N__38510),
            .I(N__38503));
    InMux I__5116 (
            .O(N__38507),
            .I(N__38500));
    InMux I__5115 (
            .O(N__38506),
            .I(N__38497));
    Odrv4 I__5114 (
            .O(N__38503),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    LocalMux I__5113 (
            .O(N__38500),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    LocalMux I__5112 (
            .O(N__38497),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    SRMux I__5111 (
            .O(N__38490),
            .I(N__38485));
    SRMux I__5110 (
            .O(N__38489),
            .I(N__38482));
    SRMux I__5109 (
            .O(N__38488),
            .I(N__38478));
    LocalMux I__5108 (
            .O(N__38485),
            .I(N__38473));
    LocalMux I__5107 (
            .O(N__38482),
            .I(N__38473));
    SRMux I__5106 (
            .O(N__38481),
            .I(N__38470));
    LocalMux I__5105 (
            .O(N__38478),
            .I(N__38467));
    Span4Mux_v I__5104 (
            .O(N__38473),
            .I(N__38462));
    LocalMux I__5103 (
            .O(N__38470),
            .I(N__38462));
    Span4Mux_h I__5102 (
            .O(N__38467),
            .I(N__38458));
    Span4Mux_v I__5101 (
            .O(N__38462),
            .I(N__38455));
    InMux I__5100 (
            .O(N__38461),
            .I(N__38452));
    Odrv4 I__5099 (
            .O(N__38458),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__5098 (
            .O(N__38455),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__5097 (
            .O(N__38452),
            .I(\pid_alt.un1_reset_0_i ));
    InMux I__5096 (
            .O(N__38445),
            .I(N__38442));
    LocalMux I__5095 (
            .O(N__38442),
            .I(N__38439));
    Span12Mux_h I__5094 (
            .O(N__38439),
            .I(N__38436));
    Odrv12 I__5093 (
            .O(N__38436),
            .I(\pid_front.O_0_3 ));
    InMux I__5092 (
            .O(N__38433),
            .I(N__38430));
    LocalMux I__5091 (
            .O(N__38430),
            .I(N__38427));
    Span4Mux_h I__5090 (
            .O(N__38427),
            .I(N__38424));
    Span4Mux_h I__5089 (
            .O(N__38424),
            .I(N__38421));
    Odrv4 I__5088 (
            .O(N__38421),
            .I(\pid_front.O_0_6 ));
    CascadeMux I__5087 (
            .O(N__38418),
            .I(\dron_frame_decoder_1.WDT10_0_cascade_ ));
    InMux I__5086 (
            .O(N__38415),
            .I(N__38411));
    InMux I__5085 (
            .O(N__38414),
            .I(N__38408));
    LocalMux I__5084 (
            .O(N__38411),
            .I(N__38405));
    LocalMux I__5083 (
            .O(N__38408),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    Odrv12 I__5082 (
            .O(N__38405),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    InMux I__5081 (
            .O(N__38400),
            .I(N__38397));
    LocalMux I__5080 (
            .O(N__38397),
            .I(N__38394));
    Span4Mux_v I__5079 (
            .O(N__38394),
            .I(N__38391));
    Span4Mux_v I__5078 (
            .O(N__38391),
            .I(N__38388));
    Odrv4 I__5077 (
            .O(N__38388),
            .I(\Commands_frame_decoder.source_CH1data_1_sqmuxa ));
    CascadeMux I__5076 (
            .O(N__38385),
            .I(\Commands_frame_decoder.source_CH1data_1_sqmuxa_cascade_ ));
    InMux I__5075 (
            .O(N__38382),
            .I(N__38376));
    InMux I__5074 (
            .O(N__38381),
            .I(N__38376));
    LocalMux I__5073 (
            .O(N__38376),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    CascadeMux I__5072 (
            .O(N__38373),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ));
    InMux I__5071 (
            .O(N__38370),
            .I(N__38366));
    InMux I__5070 (
            .O(N__38369),
            .I(N__38363));
    LocalMux I__5069 (
            .O(N__38366),
            .I(N__38360));
    LocalMux I__5068 (
            .O(N__38363),
            .I(N__38357));
    Span4Mux_v I__5067 (
            .O(N__38360),
            .I(N__38354));
    Span4Mux_v I__5066 (
            .O(N__38357),
            .I(N__38351));
    Span4Mux_h I__5065 (
            .O(N__38354),
            .I(N__38348));
    Span4Mux_h I__5064 (
            .O(N__38351),
            .I(N__38345));
    Span4Mux_h I__5063 (
            .O(N__38348),
            .I(N__38342));
    Span4Mux_h I__5062 (
            .O(N__38345),
            .I(N__38336));
    Span4Mux_h I__5061 (
            .O(N__38342),
            .I(N__38336));
    InMux I__5060 (
            .O(N__38341),
            .I(N__38333));
    Span4Mux_h I__5059 (
            .O(N__38336),
            .I(N__38330));
    LocalMux I__5058 (
            .O(N__38333),
            .I(xy_kp_4));
    Odrv4 I__5057 (
            .O(N__38330),
            .I(xy_kp_4));
    CEMux I__5056 (
            .O(N__38325),
            .I(N__38322));
    LocalMux I__5055 (
            .O(N__38322),
            .I(N__38319));
    Span4Mux_s3_h I__5054 (
            .O(N__38319),
            .I(N__38316));
    Span4Mux_h I__5053 (
            .O(N__38316),
            .I(N__38313));
    Odrv4 I__5052 (
            .O(N__38313),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    CEMux I__5051 (
            .O(N__38310),
            .I(N__38305));
    CEMux I__5050 (
            .O(N__38309),
            .I(N__38302));
    CEMux I__5049 (
            .O(N__38308),
            .I(N__38299));
    LocalMux I__5048 (
            .O(N__38305),
            .I(N__38296));
    LocalMux I__5047 (
            .O(N__38302),
            .I(N__38293));
    LocalMux I__5046 (
            .O(N__38299),
            .I(N__38290));
    Span4Mux_v I__5045 (
            .O(N__38296),
            .I(N__38285));
    Span4Mux_s3_h I__5044 (
            .O(N__38293),
            .I(N__38285));
    Span4Mux_v I__5043 (
            .O(N__38290),
            .I(N__38282));
    Span4Mux_v I__5042 (
            .O(N__38285),
            .I(N__38279));
    Span4Mux_h I__5041 (
            .O(N__38282),
            .I(N__38276));
    Span4Mux_h I__5040 (
            .O(N__38279),
            .I(N__38273));
    Odrv4 I__5039 (
            .O(N__38276),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    Odrv4 I__5038 (
            .O(N__38273),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    CascadeMux I__5037 (
            .O(N__38268),
            .I(\uart_pc.N_152_cascade_ ));
    CascadeMux I__5036 (
            .O(N__38265),
            .I(\uart_pc.CO0_cascade_ ));
    CascadeMux I__5035 (
            .O(N__38262),
            .I(N__38258));
    InMux I__5034 (
            .O(N__38261),
            .I(N__38250));
    InMux I__5033 (
            .O(N__38258),
            .I(N__38250));
    InMux I__5032 (
            .O(N__38257),
            .I(N__38250));
    LocalMux I__5031 (
            .O(N__38250),
            .I(N__38246));
    InMux I__5030 (
            .O(N__38249),
            .I(N__38243));
    Odrv4 I__5029 (
            .O(N__38246),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__5028 (
            .O(N__38243),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__5027 (
            .O(N__38238),
            .I(N__38232));
    InMux I__5026 (
            .O(N__38237),
            .I(N__38232));
    LocalMux I__5025 (
            .O(N__38232),
            .I(\uart_pc.un1_state_7_0 ));
    CascadeMux I__5024 (
            .O(N__38229),
            .I(N__38226));
    InMux I__5023 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__5022 (
            .O(N__38223),
            .I(N__38219));
    InMux I__5021 (
            .O(N__38222),
            .I(N__38216));
    Odrv12 I__5020 (
            .O(N__38219),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__5019 (
            .O(N__38216),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__5018 (
            .O(N__38211),
            .I(N__38206));
    InMux I__5017 (
            .O(N__38210),
            .I(N__38199));
    InMux I__5016 (
            .O(N__38209),
            .I(N__38199));
    InMux I__5015 (
            .O(N__38206),
            .I(N__38199));
    LocalMux I__5014 (
            .O(N__38199),
            .I(\uart_pc.stateZ0Z_1 ));
    InMux I__5013 (
            .O(N__38196),
            .I(N__38193));
    LocalMux I__5012 (
            .O(N__38193),
            .I(N__38189));
    InMux I__5011 (
            .O(N__38192),
            .I(N__38185));
    Span4Mux_h I__5010 (
            .O(N__38189),
            .I(N__38182));
    InMux I__5009 (
            .O(N__38188),
            .I(N__38179));
    LocalMux I__5008 (
            .O(N__38185),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    Odrv4 I__5007 (
            .O(N__38182),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__5006 (
            .O(N__38179),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    CascadeMux I__5005 (
            .O(N__38172),
            .I(\uart_pc.data_rdyc_1_cascade_ ));
    CascadeMux I__5004 (
            .O(N__38169),
            .I(N__38164));
    CascadeMux I__5003 (
            .O(N__38168),
            .I(N__38161));
    InMux I__5002 (
            .O(N__38167),
            .I(N__38152));
    InMux I__5001 (
            .O(N__38164),
            .I(N__38152));
    InMux I__5000 (
            .O(N__38161),
            .I(N__38152));
    InMux I__4999 (
            .O(N__38160),
            .I(N__38149));
    InMux I__4998 (
            .O(N__38159),
            .I(N__38146));
    LocalMux I__4997 (
            .O(N__38152),
            .I(N__38140));
    LocalMux I__4996 (
            .O(N__38149),
            .I(N__38135));
    LocalMux I__4995 (
            .O(N__38146),
            .I(N__38135));
    InMux I__4994 (
            .O(N__38145),
            .I(N__38130));
    InMux I__4993 (
            .O(N__38144),
            .I(N__38130));
    InMux I__4992 (
            .O(N__38143),
            .I(N__38127));
    Span4Mux_h I__4991 (
            .O(N__38140),
            .I(N__38124));
    Odrv4 I__4990 (
            .O(N__38135),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4989 (
            .O(N__38130),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__4988 (
            .O(N__38127),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__4987 (
            .O(N__38124),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__4986 (
            .O(N__38115),
            .I(N__38104));
    InMux I__4985 (
            .O(N__38114),
            .I(N__38104));
    InMux I__4984 (
            .O(N__38113),
            .I(N__38104));
    InMux I__4983 (
            .O(N__38112),
            .I(N__38096));
    InMux I__4982 (
            .O(N__38111),
            .I(N__38096));
    LocalMux I__4981 (
            .O(N__38104),
            .I(N__38092));
    InMux I__4980 (
            .O(N__38103),
            .I(N__38089));
    InMux I__4979 (
            .O(N__38102),
            .I(N__38084));
    InMux I__4978 (
            .O(N__38101),
            .I(N__38084));
    LocalMux I__4977 (
            .O(N__38096),
            .I(N__38081));
    InMux I__4976 (
            .O(N__38095),
            .I(N__38078));
    Span4Mux_v I__4975 (
            .O(N__38092),
            .I(N__38075));
    LocalMux I__4974 (
            .O(N__38089),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4973 (
            .O(N__38084),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__4972 (
            .O(N__38081),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__4971 (
            .O(N__38078),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__4970 (
            .O(N__38075),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__4969 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__4968 (
            .O(N__38061),
            .I(N__38058));
    Span4Mux_v I__4967 (
            .O(N__38058),
            .I(N__38055));
    Odrv4 I__4966 (
            .O(N__38055),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ));
    InMux I__4965 (
            .O(N__38052),
            .I(N__38049));
    LocalMux I__4964 (
            .O(N__38049),
            .I(N__38046));
    Odrv12 I__4963 (
            .O(N__38046),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ));
    CascadeMux I__4962 (
            .O(N__38043),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ));
    CascadeMux I__4961 (
            .O(N__38040),
            .I(N__38037));
    InMux I__4960 (
            .O(N__38037),
            .I(N__38034));
    LocalMux I__4959 (
            .O(N__38034),
            .I(N__38027));
    InMux I__4958 (
            .O(N__38033),
            .I(N__38024));
    InMux I__4957 (
            .O(N__38032),
            .I(N__38017));
    InMux I__4956 (
            .O(N__38031),
            .I(N__38017));
    InMux I__4955 (
            .O(N__38030),
            .I(N__38017));
    Span4Mux_h I__4954 (
            .O(N__38027),
            .I(N__38014));
    LocalMux I__4953 (
            .O(N__38024),
            .I(\uart_pc.N_143 ));
    LocalMux I__4952 (
            .O(N__38017),
            .I(\uart_pc.N_143 ));
    Odrv4 I__4951 (
            .O(N__38014),
            .I(\uart_pc.N_143 ));
    InMux I__4950 (
            .O(N__38007),
            .I(N__38001));
    InMux I__4949 (
            .O(N__38006),
            .I(N__38001));
    LocalMux I__4948 (
            .O(N__38001),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__4947 (
            .O(N__37998),
            .I(\uart_pc.N_145_cascade_ ));
    CascadeMux I__4946 (
            .O(N__37995),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    CascadeMux I__4945 (
            .O(N__37992),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__4944 (
            .O(N__37989),
            .I(N__37985));
    CascadeMux I__4943 (
            .O(N__37988),
            .I(N__37981));
    InMux I__4942 (
            .O(N__37985),
            .I(N__37977));
    InMux I__4941 (
            .O(N__37984),
            .I(N__37974));
    InMux I__4940 (
            .O(N__37981),
            .I(N__37971));
    InMux I__4939 (
            .O(N__37980),
            .I(N__37968));
    LocalMux I__4938 (
            .O(N__37977),
            .I(N__37965));
    LocalMux I__4937 (
            .O(N__37974),
            .I(N__37960));
    LocalMux I__4936 (
            .O(N__37971),
            .I(N__37960));
    LocalMux I__4935 (
            .O(N__37968),
            .I(N__37955));
    Span4Mux_v I__4934 (
            .O(N__37965),
            .I(N__37955));
    Odrv4 I__4933 (
            .O(N__37960),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__4932 (
            .O(N__37955),
            .I(\uart_pc.stateZ0Z_2 ));
    CascadeMux I__4931 (
            .O(N__37950),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1_0_cascade_ ));
    InMux I__4930 (
            .O(N__37947),
            .I(N__37944));
    LocalMux I__4929 (
            .O(N__37944),
            .I(\Commands_frame_decoder.N_405 ));
    InMux I__4928 (
            .O(N__37941),
            .I(N__37937));
    InMux I__4927 (
            .O(N__37940),
            .I(N__37934));
    LocalMux I__4926 (
            .O(N__37937),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    LocalMux I__4925 (
            .O(N__37934),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    CascadeMux I__4924 (
            .O(N__37929),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ));
    CascadeMux I__4923 (
            .O(N__37926),
            .I(\Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ));
    CascadeMux I__4922 (
            .O(N__37923),
            .I(N__37919));
    InMux I__4921 (
            .O(N__37922),
            .I(N__37914));
    InMux I__4920 (
            .O(N__37919),
            .I(N__37910));
    InMux I__4919 (
            .O(N__37918),
            .I(N__37905));
    InMux I__4918 (
            .O(N__37917),
            .I(N__37905));
    LocalMux I__4917 (
            .O(N__37914),
            .I(N__37902));
    InMux I__4916 (
            .O(N__37913),
            .I(N__37899));
    LocalMux I__4915 (
            .O(N__37910),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__4914 (
            .O(N__37905),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    Odrv4 I__4913 (
            .O(N__37902),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__4912 (
            .O(N__37899),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    CascadeMux I__4911 (
            .O(N__37890),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ));
    InMux I__4910 (
            .O(N__37887),
            .I(N__37880));
    InMux I__4909 (
            .O(N__37886),
            .I(N__37880));
    InMux I__4908 (
            .O(N__37885),
            .I(N__37877));
    LocalMux I__4907 (
            .O(N__37880),
            .I(\Commands_frame_decoder.N_409 ));
    LocalMux I__4906 (
            .O(N__37877),
            .I(\Commands_frame_decoder.N_409 ));
    CascadeMux I__4905 (
            .O(N__37872),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_3_2_cascade_ ));
    InMux I__4904 (
            .O(N__37869),
            .I(N__37866));
    LocalMux I__4903 (
            .O(N__37866),
            .I(N__37862));
    InMux I__4902 (
            .O(N__37865),
            .I(N__37859));
    Odrv4 I__4901 (
            .O(N__37862),
            .I(\Commands_frame_decoder.N_371 ));
    LocalMux I__4900 (
            .O(N__37859),
            .I(\Commands_frame_decoder.N_371 ));
    InMux I__4899 (
            .O(N__37854),
            .I(N__37848));
    InMux I__4898 (
            .O(N__37853),
            .I(N__37848));
    LocalMux I__4897 (
            .O(N__37848),
            .I(N__37843));
    InMux I__4896 (
            .O(N__37847),
            .I(N__37838));
    InMux I__4895 (
            .O(N__37846),
            .I(N__37838));
    Span4Mux_h I__4894 (
            .O(N__37843),
            .I(N__37835));
    LocalMux I__4893 (
            .O(N__37838),
            .I(N__37832));
    Odrv4 I__4892 (
            .O(N__37835),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    Odrv4 I__4891 (
            .O(N__37832),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    InMux I__4890 (
            .O(N__37827),
            .I(N__37824));
    LocalMux I__4889 (
            .O(N__37824),
            .I(N__37820));
    InMux I__4888 (
            .O(N__37823),
            .I(N__37817));
    Span12Mux_s5_h I__4887 (
            .O(N__37820),
            .I(N__37814));
    LocalMux I__4886 (
            .O(N__37817),
            .I(alt_kp_4));
    Odrv12 I__4885 (
            .O(N__37814),
            .I(alt_kp_4));
    CascadeMux I__4884 (
            .O(N__37809),
            .I(\Commands_frame_decoder.N_369_2_cascade_ ));
    CascadeMux I__4883 (
            .O(N__37806),
            .I(\Commands_frame_decoder.N_370_cascade_ ));
    InMux I__4882 (
            .O(N__37803),
            .I(N__37800));
    LocalMux I__4881 (
            .O(N__37800),
            .I(\Commands_frame_decoder.N_369_2 ));
    CascadeMux I__4880 (
            .O(N__37797),
            .I(N__37794));
    InMux I__4879 (
            .O(N__37794),
            .I(N__37791));
    LocalMux I__4878 (
            .O(N__37791),
            .I(N__37787));
    CascadeMux I__4877 (
            .O(N__37790),
            .I(N__37784));
    Span4Mux_h I__4876 (
            .O(N__37787),
            .I(N__37780));
    InMux I__4875 (
            .O(N__37784),
            .I(N__37775));
    InMux I__4874 (
            .O(N__37783),
            .I(N__37775));
    Odrv4 I__4873 (
            .O(N__37780),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    LocalMux I__4872 (
            .O(N__37775),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    InMux I__4871 (
            .O(N__37770),
            .I(N__37767));
    LocalMux I__4870 (
            .O(N__37767),
            .I(\Commands_frame_decoder.state_ns_i_0_0 ));
    CascadeMux I__4869 (
            .O(N__37764),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ));
    InMux I__4868 (
            .O(N__37761),
            .I(N__37754));
    InMux I__4867 (
            .O(N__37760),
            .I(N__37754));
    InMux I__4866 (
            .O(N__37759),
            .I(N__37751));
    LocalMux I__4865 (
            .O(N__37754),
            .I(N__37748));
    LocalMux I__4864 (
            .O(N__37751),
            .I(N__37745));
    Span4Mux_h I__4863 (
            .O(N__37748),
            .I(N__37742));
    Odrv12 I__4862 (
            .O(N__37745),
            .I(\pid_alt.un2_pid_prereg_cry_14_c_RNINTBA ));
    Odrv4 I__4861 (
            .O(N__37742),
            .I(\pid_alt.un2_pid_prereg_cry_14_c_RNINTBA ));
    CascadeMux I__4860 (
            .O(N__37737),
            .I(N__37733));
    InMux I__4859 (
            .O(N__37736),
            .I(N__37730));
    InMux I__4858 (
            .O(N__37733),
            .I(N__37727));
    LocalMux I__4857 (
            .O(N__37730),
            .I(N__37724));
    LocalMux I__4856 (
            .O(N__37727),
            .I(N__37721));
    Odrv4 I__4855 (
            .O(N__37724),
            .I(\pid_alt.error_d_reg_prev_esr_RNICEFN1Z0Z_14 ));
    Odrv4 I__4854 (
            .O(N__37721),
            .I(\pid_alt.error_d_reg_prev_esr_RNICEFN1Z0Z_14 ));
    InMux I__4853 (
            .O(N__37716),
            .I(N__37712));
    InMux I__4852 (
            .O(N__37715),
            .I(N__37709));
    LocalMux I__4851 (
            .O(N__37712),
            .I(N__37704));
    LocalMux I__4850 (
            .O(N__37709),
            .I(N__37704));
    Span4Mux_h I__4849 (
            .O(N__37704),
            .I(N__37701));
    Span4Mux_v I__4848 (
            .O(N__37701),
            .I(N__37698));
    Span4Mux_s2_h I__4847 (
            .O(N__37698),
            .I(N__37695));
    Odrv4 I__4846 (
            .O(N__37695),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__4845 (
            .O(N__37692),
            .I(N__37689));
    LocalMux I__4844 (
            .O(N__37689),
            .I(N__37685));
    InMux I__4843 (
            .O(N__37688),
            .I(N__37682));
    Span4Mux_v I__4842 (
            .O(N__37685),
            .I(N__37679));
    LocalMux I__4841 (
            .O(N__37682),
            .I(N__37676));
    Span4Mux_v I__4840 (
            .O(N__37679),
            .I(N__37673));
    Odrv12 I__4839 (
            .O(N__37676),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    Odrv4 I__4838 (
            .O(N__37673),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    InMux I__4837 (
            .O(N__37668),
            .I(N__37664));
    InMux I__4836 (
            .O(N__37667),
            .I(N__37661));
    LocalMux I__4835 (
            .O(N__37664),
            .I(N__37657));
    LocalMux I__4834 (
            .O(N__37661),
            .I(N__37654));
    InMux I__4833 (
            .O(N__37660),
            .I(N__37651));
    Span4Mux_v I__4832 (
            .O(N__37657),
            .I(N__37648));
    Sp12to4 I__4831 (
            .O(N__37654),
            .I(N__37645));
    LocalMux I__4830 (
            .O(N__37651),
            .I(N__37640));
    Span4Mux_v I__4829 (
            .O(N__37648),
            .I(N__37640));
    Span12Mux_v I__4828 (
            .O(N__37645),
            .I(N__37637));
    Odrv4 I__4827 (
            .O(N__37640),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    Odrv12 I__4826 (
            .O(N__37637),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__4825 (
            .O(N__37632),
            .I(N__37626));
    InMux I__4824 (
            .O(N__37631),
            .I(N__37626));
    LocalMux I__4823 (
            .O(N__37626),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    InMux I__4822 (
            .O(N__37623),
            .I(N__37617));
    InMux I__4821 (
            .O(N__37622),
            .I(N__37617));
    LocalMux I__4820 (
            .O(N__37617),
            .I(N__37614));
    Span4Mux_v I__4819 (
            .O(N__37614),
            .I(N__37611));
    Span4Mux_h I__4818 (
            .O(N__37611),
            .I(N__37608));
    Odrv4 I__4817 (
            .O(N__37608),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    InMux I__4816 (
            .O(N__37605),
            .I(N__37602));
    LocalMux I__4815 (
            .O(N__37602),
            .I(N__37598));
    CascadeMux I__4814 (
            .O(N__37601),
            .I(N__37595));
    Span4Mux_v I__4813 (
            .O(N__37598),
            .I(N__37592));
    InMux I__4812 (
            .O(N__37595),
            .I(N__37589));
    Odrv4 I__4811 (
            .O(N__37592),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG0FQ1Z0Z_12 ));
    LocalMux I__4810 (
            .O(N__37589),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG0FQ1Z0Z_12 ));
    CascadeMux I__4809 (
            .O(N__37584),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__4808 (
            .O(N__37581),
            .I(N__37578));
    LocalMux I__4807 (
            .O(N__37578),
            .I(N__37575));
    Span4Mux_v I__4806 (
            .O(N__37575),
            .I(N__37572));
    Odrv4 I__4805 (
            .O(N__37572),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK5TH3Z0Z_13 ));
    InMux I__4804 (
            .O(N__37569),
            .I(N__37560));
    InMux I__4803 (
            .O(N__37568),
            .I(N__37560));
    InMux I__4802 (
            .O(N__37567),
            .I(N__37560));
    LocalMux I__4801 (
            .O(N__37560),
            .I(N__37557));
    Span4Mux_v I__4800 (
            .O(N__37557),
            .I(N__37554));
    Span4Mux_v I__4799 (
            .O(N__37554),
            .I(N__37551));
    Span4Mux_h I__4798 (
            .O(N__37551),
            .I(N__37548));
    Odrv4 I__4797 (
            .O(N__37548),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    CascadeMux I__4796 (
            .O(N__37545),
            .I(N__37542));
    InMux I__4795 (
            .O(N__37542),
            .I(N__37536));
    InMux I__4794 (
            .O(N__37541),
            .I(N__37536));
    LocalMux I__4793 (
            .O(N__37536),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    CEMux I__4792 (
            .O(N__37533),
            .I(N__37479));
    CEMux I__4791 (
            .O(N__37532),
            .I(N__37479));
    CEMux I__4790 (
            .O(N__37531),
            .I(N__37479));
    CEMux I__4789 (
            .O(N__37530),
            .I(N__37479));
    CEMux I__4788 (
            .O(N__37529),
            .I(N__37479));
    CEMux I__4787 (
            .O(N__37528),
            .I(N__37479));
    CEMux I__4786 (
            .O(N__37527),
            .I(N__37479));
    CEMux I__4785 (
            .O(N__37526),
            .I(N__37479));
    CEMux I__4784 (
            .O(N__37525),
            .I(N__37479));
    CEMux I__4783 (
            .O(N__37524),
            .I(N__37479));
    CEMux I__4782 (
            .O(N__37523),
            .I(N__37479));
    CEMux I__4781 (
            .O(N__37522),
            .I(N__37479));
    CEMux I__4780 (
            .O(N__37521),
            .I(N__37479));
    CEMux I__4779 (
            .O(N__37520),
            .I(N__37479));
    CEMux I__4778 (
            .O(N__37519),
            .I(N__37479));
    CEMux I__4777 (
            .O(N__37518),
            .I(N__37479));
    CEMux I__4776 (
            .O(N__37517),
            .I(N__37479));
    CEMux I__4775 (
            .O(N__37516),
            .I(N__37479));
    GlobalMux I__4774 (
            .O(N__37479),
            .I(N__37476));
    gio2CtrlBuf I__4773 (
            .O(N__37476),
            .I(\pid_alt.state_0_g_0 ));
    InMux I__4772 (
            .O(N__37473),
            .I(N__37470));
    LocalMux I__4771 (
            .O(N__37470),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    InMux I__4770 (
            .O(N__37467),
            .I(N__37461));
    InMux I__4769 (
            .O(N__37466),
            .I(N__37461));
    LocalMux I__4768 (
            .O(N__37461),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__4767 (
            .O(N__37458),
            .I(N__37453));
    InMux I__4766 (
            .O(N__37457),
            .I(N__37448));
    InMux I__4765 (
            .O(N__37456),
            .I(N__37448));
    LocalMux I__4764 (
            .O(N__37453),
            .I(N__37445));
    LocalMux I__4763 (
            .O(N__37448),
            .I(N__37442));
    Span4Mux_v I__4762 (
            .O(N__37445),
            .I(N__37439));
    Span4Mux_h I__4761 (
            .O(N__37442),
            .I(N__37436));
    Odrv4 I__4760 (
            .O(N__37439),
            .I(\pid_alt.un2_pid_prereg_cry_13_c_RNILQAA ));
    Odrv4 I__4759 (
            .O(N__37436),
            .I(\pid_alt.un2_pid_prereg_cry_13_c_RNILQAA ));
    CascadeMux I__4758 (
            .O(N__37431),
            .I(N__37427));
    CascadeMux I__4757 (
            .O(N__37430),
            .I(N__37424));
    InMux I__4756 (
            .O(N__37427),
            .I(N__37421));
    InMux I__4755 (
            .O(N__37424),
            .I(N__37418));
    LocalMux I__4754 (
            .O(N__37421),
            .I(N__37415));
    LocalMux I__4753 (
            .O(N__37418),
            .I(\pid_alt.error_d_reg_prev_esr_RNI45EN1Z0Z_13 ));
    Odrv4 I__4752 (
            .O(N__37415),
            .I(\pid_alt.error_d_reg_prev_esr_RNI45EN1Z0Z_13 ));
    CEMux I__4751 (
            .O(N__37410),
            .I(N__37406));
    CEMux I__4750 (
            .O(N__37409),
            .I(N__37403));
    LocalMux I__4749 (
            .O(N__37406),
            .I(N__37400));
    LocalMux I__4748 (
            .O(N__37403),
            .I(N__37397));
    Span4Mux_h I__4747 (
            .O(N__37400),
            .I(N__37394));
    Span4Mux_h I__4746 (
            .O(N__37397),
            .I(N__37391));
    Span4Mux_h I__4745 (
            .O(N__37394),
            .I(N__37388));
    Odrv4 I__4744 (
            .O(N__37391),
            .I(\Commands_frame_decoder.source_CH1data_1_sqmuxa_0 ));
    Odrv4 I__4743 (
            .O(N__37388),
            .I(\Commands_frame_decoder.source_CH1data_1_sqmuxa_0 ));
    InMux I__4742 (
            .O(N__37383),
            .I(N__37378));
    InMux I__4741 (
            .O(N__37382),
            .I(N__37375));
    InMux I__4740 (
            .O(N__37381),
            .I(N__37372));
    LocalMux I__4739 (
            .O(N__37378),
            .I(N__37369));
    LocalMux I__4738 (
            .O(N__37375),
            .I(N__37366));
    LocalMux I__4737 (
            .O(N__37372),
            .I(\pid_alt.N_90 ));
    Odrv4 I__4736 (
            .O(N__37369),
            .I(\pid_alt.N_90 ));
    Odrv4 I__4735 (
            .O(N__37366),
            .I(\pid_alt.N_90 ));
    CascadeMux I__4734 (
            .O(N__37359),
            .I(N__37355));
    InMux I__4733 (
            .O(N__37358),
            .I(N__37350));
    InMux I__4732 (
            .O(N__37355),
            .I(N__37350));
    LocalMux I__4731 (
            .O(N__37350),
            .I(N__37347));
    Span4Mux_v I__4730 (
            .O(N__37347),
            .I(N__37341));
    InMux I__4729 (
            .O(N__37346),
            .I(N__37338));
    InMux I__4728 (
            .O(N__37345),
            .I(N__37335));
    InMux I__4727 (
            .O(N__37344),
            .I(N__37332));
    Odrv4 I__4726 (
            .O(N__37341),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    LocalMux I__4725 (
            .O(N__37338),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    LocalMux I__4724 (
            .O(N__37335),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    LocalMux I__4723 (
            .O(N__37332),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    CascadeMux I__4722 (
            .O(N__37323),
            .I(\pid_alt.source_pid_9_0_0_4_cascade_ ));
    InMux I__4721 (
            .O(N__37320),
            .I(N__37314));
    InMux I__4720 (
            .O(N__37319),
            .I(N__37314));
    LocalMux I__4719 (
            .O(N__37314),
            .I(N__37311));
    Odrv4 I__4718 (
            .O(N__37311),
            .I(\pid_alt.N_44 ));
    InMux I__4717 (
            .O(N__37308),
            .I(N__37305));
    LocalMux I__4716 (
            .O(N__37305),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__4715 (
            .O(N__37302),
            .I(N__37299));
    LocalMux I__4714 (
            .O(N__37299),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    CascadeMux I__4713 (
            .O(N__37296),
            .I(N__37293));
    InMux I__4712 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__4711 (
            .O(N__37290),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    InMux I__4710 (
            .O(N__37287),
            .I(N__37284));
    LocalMux I__4709 (
            .O(N__37284),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    InMux I__4708 (
            .O(N__37281),
            .I(N__37278));
    LocalMux I__4707 (
            .O(N__37278),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__4706 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__4705 (
            .O(N__37272),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    CascadeMux I__4704 (
            .O(N__37269),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ));
    InMux I__4703 (
            .O(N__37266),
            .I(N__37263));
    LocalMux I__4702 (
            .O(N__37263),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ));
    InMux I__4701 (
            .O(N__37260),
            .I(N__37252));
    InMux I__4700 (
            .O(N__37259),
            .I(N__37249));
    InMux I__4699 (
            .O(N__37258),
            .I(N__37236));
    InMux I__4698 (
            .O(N__37257),
            .I(N__37236));
    InMux I__4697 (
            .O(N__37256),
            .I(N__37236));
    InMux I__4696 (
            .O(N__37255),
            .I(N__37236));
    LocalMux I__4695 (
            .O(N__37252),
            .I(N__37231));
    LocalMux I__4694 (
            .O(N__37249),
            .I(N__37231));
    InMux I__4693 (
            .O(N__37248),
            .I(N__37221));
    InMux I__4692 (
            .O(N__37247),
            .I(N__37221));
    InMux I__4691 (
            .O(N__37246),
            .I(N__37221));
    InMux I__4690 (
            .O(N__37245),
            .I(N__37221));
    LocalMux I__4689 (
            .O(N__37236),
            .I(N__37216));
    Span4Mux_h I__4688 (
            .O(N__37231),
            .I(N__37216));
    InMux I__4687 (
            .O(N__37230),
            .I(N__37213));
    LocalMux I__4686 (
            .O(N__37221),
            .I(\pid_alt.N_216 ));
    Odrv4 I__4685 (
            .O(N__37216),
            .I(\pid_alt.N_216 ));
    LocalMux I__4684 (
            .O(N__37213),
            .I(\pid_alt.N_216 ));
    InMux I__4683 (
            .O(N__37206),
            .I(N__37203));
    LocalMux I__4682 (
            .O(N__37203),
            .I(N__37196));
    InMux I__4681 (
            .O(N__37202),
            .I(N__37193));
    InMux I__4680 (
            .O(N__37201),
            .I(N__37189));
    InMux I__4679 (
            .O(N__37200),
            .I(N__37184));
    InMux I__4678 (
            .O(N__37199),
            .I(N__37184));
    Span4Mux_h I__4677 (
            .O(N__37196),
            .I(N__37181));
    LocalMux I__4676 (
            .O(N__37193),
            .I(N__37178));
    InMux I__4675 (
            .O(N__37192),
            .I(N__37175));
    LocalMux I__4674 (
            .O(N__37189),
            .I(N__37172));
    LocalMux I__4673 (
            .O(N__37184),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4672 (
            .O(N__37181),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4671 (
            .O(N__37178),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    LocalMux I__4670 (
            .O(N__37175),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__4669 (
            .O(N__37172),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    CascadeMux I__4668 (
            .O(N__37161),
            .I(N__37156));
    CascadeMux I__4667 (
            .O(N__37160),
            .I(N__37151));
    InMux I__4666 (
            .O(N__37159),
            .I(N__37139));
    InMux I__4665 (
            .O(N__37156),
            .I(N__37139));
    InMux I__4664 (
            .O(N__37155),
            .I(N__37139));
    InMux I__4663 (
            .O(N__37154),
            .I(N__37139));
    InMux I__4662 (
            .O(N__37151),
            .I(N__37136));
    CascadeMux I__4661 (
            .O(N__37150),
            .I(N__37133));
    CascadeMux I__4660 (
            .O(N__37149),
            .I(N__37130));
    CascadeMux I__4659 (
            .O(N__37148),
            .I(N__37127));
    LocalMux I__4658 (
            .O(N__37139),
            .I(N__37122));
    LocalMux I__4657 (
            .O(N__37136),
            .I(N__37119));
    InMux I__4656 (
            .O(N__37133),
            .I(N__37116));
    InMux I__4655 (
            .O(N__37130),
            .I(N__37107));
    InMux I__4654 (
            .O(N__37127),
            .I(N__37107));
    InMux I__4653 (
            .O(N__37126),
            .I(N__37107));
    InMux I__4652 (
            .O(N__37125),
            .I(N__37107));
    Span4Mux_v I__4651 (
            .O(N__37122),
            .I(N__37104));
    Span4Mux_h I__4650 (
            .O(N__37119),
            .I(N__37101));
    LocalMux I__4649 (
            .O(N__37116),
            .I(N__37098));
    LocalMux I__4648 (
            .O(N__37107),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__4647 (
            .O(N__37104),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__4646 (
            .O(N__37101),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv12 I__4645 (
            .O(N__37098),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    CascadeMux I__4644 (
            .O(N__37089),
            .I(\pid_alt.N_216_cascade_ ));
    InMux I__4643 (
            .O(N__37086),
            .I(N__37083));
    LocalMux I__4642 (
            .O(N__37083),
            .I(N__37078));
    InMux I__4641 (
            .O(N__37082),
            .I(N__37074));
    InMux I__4640 (
            .O(N__37081),
            .I(N__37071));
    Span4Mux_v I__4639 (
            .O(N__37078),
            .I(N__37068));
    InMux I__4638 (
            .O(N__37077),
            .I(N__37065));
    LocalMux I__4637 (
            .O(N__37074),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    LocalMux I__4636 (
            .O(N__37071),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__4635 (
            .O(N__37068),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    LocalMux I__4634 (
            .O(N__37065),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    CEMux I__4633 (
            .O(N__37056),
            .I(N__37052));
    CEMux I__4632 (
            .O(N__37055),
            .I(N__37049));
    LocalMux I__4631 (
            .O(N__37052),
            .I(N__37044));
    LocalMux I__4630 (
            .O(N__37049),
            .I(N__37044));
    Odrv4 I__4629 (
            .O(N__37044),
            .I(\pid_alt.N_76_i_1 ));
    InMux I__4628 (
            .O(N__37041),
            .I(N__37038));
    LocalMux I__4627 (
            .O(N__37038),
            .I(N__37033));
    CascadeMux I__4626 (
            .O(N__37037),
            .I(N__37030));
    CascadeMux I__4625 (
            .O(N__37036),
            .I(N__37025));
    Span4Mux_v I__4624 (
            .O(N__37033),
            .I(N__37022));
    InMux I__4623 (
            .O(N__37030),
            .I(N__37013));
    InMux I__4622 (
            .O(N__37029),
            .I(N__37013));
    InMux I__4621 (
            .O(N__37028),
            .I(N__37013));
    InMux I__4620 (
            .O(N__37025),
            .I(N__37013));
    Span4Mux_v I__4619 (
            .O(N__37022),
            .I(N__37009));
    LocalMux I__4618 (
            .O(N__37013),
            .I(N__37006));
    InMux I__4617 (
            .O(N__37012),
            .I(N__37003));
    Odrv4 I__4616 (
            .O(N__37009),
            .I(\pid_alt.error_i_acumm7lto4 ));
    Odrv4 I__4615 (
            .O(N__37006),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__4614 (
            .O(N__37003),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__4613 (
            .O(N__36996),
            .I(N__36993));
    LocalMux I__4612 (
            .O(N__36993),
            .I(N__36990));
    Span4Mux_v I__4611 (
            .O(N__36990),
            .I(N__36979));
    InMux I__4610 (
            .O(N__36989),
            .I(N__36966));
    InMux I__4609 (
            .O(N__36988),
            .I(N__36966));
    InMux I__4608 (
            .O(N__36987),
            .I(N__36966));
    InMux I__4607 (
            .O(N__36986),
            .I(N__36966));
    InMux I__4606 (
            .O(N__36985),
            .I(N__36966));
    InMux I__4605 (
            .O(N__36984),
            .I(N__36966));
    InMux I__4604 (
            .O(N__36983),
            .I(N__36961));
    InMux I__4603 (
            .O(N__36982),
            .I(N__36961));
    Span4Mux_v I__4602 (
            .O(N__36979),
            .I(N__36958));
    LocalMux I__4601 (
            .O(N__36966),
            .I(N__36953));
    LocalMux I__4600 (
            .O(N__36961),
            .I(N__36953));
    Odrv4 I__4599 (
            .O(N__36958),
            .I(\pid_alt.N_93 ));
    Odrv4 I__4598 (
            .O(N__36953),
            .I(\pid_alt.N_93 ));
    InMux I__4597 (
            .O(N__36948),
            .I(N__36945));
    LocalMux I__4596 (
            .O(N__36945),
            .I(N__36942));
    Span4Mux_h I__4595 (
            .O(N__36942),
            .I(N__36939));
    Odrv4 I__4594 (
            .O(N__36939),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    CEMux I__4593 (
            .O(N__36936),
            .I(N__36932));
    CEMux I__4592 (
            .O(N__36935),
            .I(N__36929));
    LocalMux I__4591 (
            .O(N__36932),
            .I(N__36926));
    LocalMux I__4590 (
            .O(N__36929),
            .I(N__36923));
    Span4Mux_v I__4589 (
            .O(N__36926),
            .I(N__36919));
    Span4Mux_h I__4588 (
            .O(N__36923),
            .I(N__36916));
    CEMux I__4587 (
            .O(N__36922),
            .I(N__36913));
    Odrv4 I__4586 (
            .O(N__36919),
            .I(\pid_alt.N_76_i_0 ));
    Odrv4 I__4585 (
            .O(N__36916),
            .I(\pid_alt.N_76_i_0 ));
    LocalMux I__4584 (
            .O(N__36913),
            .I(\pid_alt.N_76_i_0 ));
    InMux I__4583 (
            .O(N__36906),
            .I(N__36903));
    LocalMux I__4582 (
            .O(N__36903),
            .I(N__36900));
    Odrv4 I__4581 (
            .O(N__36900),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGJTE3Z0Z_14 ));
    InMux I__4580 (
            .O(N__36897),
            .I(N__36894));
    LocalMux I__4579 (
            .O(N__36894),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    InMux I__4578 (
            .O(N__36891),
            .I(N__36888));
    LocalMux I__4577 (
            .O(N__36888),
            .I(N__36883));
    InMux I__4576 (
            .O(N__36887),
            .I(N__36878));
    InMux I__4575 (
            .O(N__36886),
            .I(N__36878));
    Odrv4 I__4574 (
            .O(N__36883),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    LocalMux I__4573 (
            .O(N__36878),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    InMux I__4572 (
            .O(N__36873),
            .I(N__36869));
    CascadeMux I__4571 (
            .O(N__36872),
            .I(N__36866));
    LocalMux I__4570 (
            .O(N__36869),
            .I(N__36862));
    InMux I__4569 (
            .O(N__36866),
            .I(N__36857));
    InMux I__4568 (
            .O(N__36865),
            .I(N__36857));
    Odrv4 I__4567 (
            .O(N__36862),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    LocalMux I__4566 (
            .O(N__36857),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    InMux I__4565 (
            .O(N__36852),
            .I(N__36848));
    CascadeMux I__4564 (
            .O(N__36851),
            .I(N__36844));
    LocalMux I__4563 (
            .O(N__36848),
            .I(N__36841));
    InMux I__4562 (
            .O(N__36847),
            .I(N__36836));
    InMux I__4561 (
            .O(N__36844),
            .I(N__36836));
    Odrv4 I__4560 (
            .O(N__36841),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    LocalMux I__4559 (
            .O(N__36836),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    InMux I__4558 (
            .O(N__36831),
            .I(N__36826));
    InMux I__4557 (
            .O(N__36830),
            .I(N__36821));
    InMux I__4556 (
            .O(N__36829),
            .I(N__36821));
    LocalMux I__4555 (
            .O(N__36826),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    LocalMux I__4554 (
            .O(N__36821),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__4553 (
            .O(N__36816),
            .I(N__36813));
    LocalMux I__4552 (
            .O(N__36813),
            .I(N__36810));
    Span4Mux_h I__4551 (
            .O(N__36810),
            .I(N__36805));
    InMux I__4550 (
            .O(N__36809),
            .I(N__36800));
    InMux I__4549 (
            .O(N__36808),
            .I(N__36800));
    Odrv4 I__4548 (
            .O(N__36805),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    LocalMux I__4547 (
            .O(N__36800),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    CascadeMux I__4546 (
            .O(N__36795),
            .I(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ));
    CascadeMux I__4545 (
            .O(N__36792),
            .I(\pid_alt.N_90_cascade_ ));
    InMux I__4544 (
            .O(N__36789),
            .I(N__36783));
    InMux I__4543 (
            .O(N__36788),
            .I(N__36783));
    LocalMux I__4542 (
            .O(N__36783),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    CascadeMux I__4541 (
            .O(N__36780),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ));
    InMux I__4540 (
            .O(N__36777),
            .I(N__36773));
    InMux I__4539 (
            .O(N__36776),
            .I(N__36770));
    LocalMux I__4538 (
            .O(N__36773),
            .I(\pid_alt.N_43 ));
    LocalMux I__4537 (
            .O(N__36770),
            .I(\pid_alt.N_43 ));
    InMux I__4536 (
            .O(N__36765),
            .I(N__36762));
    LocalMux I__4535 (
            .O(N__36762),
            .I(N__36759));
    Odrv4 I__4534 (
            .O(N__36759),
            .I(\pid_alt.N_48 ));
    InMux I__4533 (
            .O(N__36756),
            .I(N__36753));
    LocalMux I__4532 (
            .O(N__36753),
            .I(N__36750));
    Span4Mux_v I__4531 (
            .O(N__36750),
            .I(N__36746));
    InMux I__4530 (
            .O(N__36749),
            .I(N__36743));
    Odrv4 I__4529 (
            .O(N__36746),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    LocalMux I__4528 (
            .O(N__36743),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__4527 (
            .O(N__36738),
            .I(N__36735));
    LocalMux I__4526 (
            .O(N__36735),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    InMux I__4525 (
            .O(N__36732),
            .I(N__36729));
    LocalMux I__4524 (
            .O(N__36729),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    CascadeMux I__4523 (
            .O(N__36726),
            .I(N__36723));
    InMux I__4522 (
            .O(N__36723),
            .I(N__36720));
    LocalMux I__4521 (
            .O(N__36720),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__4520 (
            .O(N__36717),
            .I(N__36714));
    LocalMux I__4519 (
            .O(N__36714),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    CascadeMux I__4518 (
            .O(N__36711),
            .I(\pid_alt.N_44_cascade_ ));
    CascadeMux I__4517 (
            .O(N__36708),
            .I(\pid_alt.N_46_cascade_ ));
    InMux I__4516 (
            .O(N__36705),
            .I(N__36701));
    InMux I__4515 (
            .O(N__36704),
            .I(N__36698));
    LocalMux I__4514 (
            .O(N__36701),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    LocalMux I__4513 (
            .O(N__36698),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__4512 (
            .O(N__36693),
            .I(N__36689));
    InMux I__4511 (
            .O(N__36692),
            .I(N__36686));
    LocalMux I__4510 (
            .O(N__36689),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    LocalMux I__4509 (
            .O(N__36686),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    CascadeMux I__4508 (
            .O(N__36681),
            .I(N__36677));
    InMux I__4507 (
            .O(N__36680),
            .I(N__36672));
    InMux I__4506 (
            .O(N__36677),
            .I(N__36672));
    LocalMux I__4505 (
            .O(N__36672),
            .I(N__36669));
    Odrv4 I__4504 (
            .O(N__36669),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    CascadeMux I__4503 (
            .O(N__36666),
            .I(N__36662));
    CascadeMux I__4502 (
            .O(N__36665),
            .I(N__36659));
    InMux I__4501 (
            .O(N__36662),
            .I(N__36655));
    InMux I__4500 (
            .O(N__36659),
            .I(N__36650));
    InMux I__4499 (
            .O(N__36658),
            .I(N__36650));
    LocalMux I__4498 (
            .O(N__36655),
            .I(\pid_alt.N_46 ));
    LocalMux I__4497 (
            .O(N__36650),
            .I(\pid_alt.N_46 ));
    InMux I__4496 (
            .O(N__36645),
            .I(N__36639));
    InMux I__4495 (
            .O(N__36644),
            .I(N__36639));
    LocalMux I__4494 (
            .O(N__36639),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    InMux I__4493 (
            .O(N__36636),
            .I(N__36633));
    LocalMux I__4492 (
            .O(N__36633),
            .I(N__36630));
    Span12Mux_s5_v I__4491 (
            .O(N__36630),
            .I(N__36627));
    Odrv12 I__4490 (
            .O(N__36627),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    CascadeMux I__4489 (
            .O(N__36624),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ));
    InMux I__4488 (
            .O(N__36621),
            .I(N__36618));
    LocalMux I__4487 (
            .O(N__36618),
            .I(N__36615));
    Odrv4 I__4486 (
            .O(N__36615),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ));
    InMux I__4485 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__4484 (
            .O(N__36609),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ));
    CascadeMux I__4483 (
            .O(N__36606),
            .I(N__36603));
    InMux I__4482 (
            .O(N__36603),
            .I(N__36599));
    InMux I__4481 (
            .O(N__36602),
            .I(N__36596));
    LocalMux I__4480 (
            .O(N__36599),
            .I(N__36593));
    LocalMux I__4479 (
            .O(N__36596),
            .I(\uart_pc.N_126_li ));
    Odrv4 I__4478 (
            .O(N__36593),
            .I(\uart_pc.N_126_li ));
    CascadeMux I__4477 (
            .O(N__36588),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__4476 (
            .O(N__36585),
            .I(\pid_alt.source_pid_9_0_tz_6_cascade_ ));
    InMux I__4475 (
            .O(N__36582),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__4474 (
            .O(N__36579),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    CascadeMux I__4473 (
            .O(N__36576),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ));
    InMux I__4472 (
            .O(N__36573),
            .I(N__36570));
    LocalMux I__4471 (
            .O(N__36570),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    CascadeMux I__4470 (
            .O(N__36567),
            .I(\uart_pc.timer_Count_0_sqmuxa_cascade_ ));
    InMux I__4469 (
            .O(N__36564),
            .I(N__36561));
    LocalMux I__4468 (
            .O(N__36561),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    CascadeMux I__4467 (
            .O(N__36558),
            .I(N__36552));
    InMux I__4466 (
            .O(N__36557),
            .I(N__36547));
    InMux I__4465 (
            .O(N__36556),
            .I(N__36547));
    InMux I__4464 (
            .O(N__36555),
            .I(N__36542));
    InMux I__4463 (
            .O(N__36552),
            .I(N__36542));
    LocalMux I__4462 (
            .O(N__36547),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4461 (
            .O(N__36542),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__4460 (
            .O(N__36537),
            .I(N__36534));
    LocalMux I__4459 (
            .O(N__36534),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    CascadeMux I__4458 (
            .O(N__36531),
            .I(\uart_pc.N_126_li_cascade_ ));
    IoInMux I__4457 (
            .O(N__36528),
            .I(N__36525));
    LocalMux I__4456 (
            .O(N__36525),
            .I(N__36522));
    Span4Mux_s3_v I__4455 (
            .O(N__36522),
            .I(N__36519));
    Span4Mux_h I__4454 (
            .O(N__36519),
            .I(N__36516));
    Span4Mux_h I__4453 (
            .O(N__36516),
            .I(N__36513));
    Span4Mux_h I__4452 (
            .O(N__36513),
            .I(N__36510));
    Odrv4 I__4451 (
            .O(N__36510),
            .I(\pid_alt.N_579_0 ));
    CascadeMux I__4450 (
            .O(N__36507),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ));
    CascadeMux I__4449 (
            .O(N__36504),
            .I(\uart_pc.N_143_cascade_ ));
    InMux I__4448 (
            .O(N__36501),
            .I(N__36497));
    InMux I__4447 (
            .O(N__36500),
            .I(N__36494));
    LocalMux I__4446 (
            .O(N__36497),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__4445 (
            .O(N__36494),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    CascadeMux I__4444 (
            .O(N__36489),
            .I(N__36483));
    InMux I__4443 (
            .O(N__36488),
            .I(N__36480));
    InMux I__4442 (
            .O(N__36487),
            .I(N__36477));
    InMux I__4441 (
            .O(N__36486),
            .I(N__36472));
    InMux I__4440 (
            .O(N__36483),
            .I(N__36472));
    LocalMux I__4439 (
            .O(N__36480),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4438 (
            .O(N__36477),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4437 (
            .O(N__36472),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__4436 (
            .O(N__36465),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    CascadeMux I__4435 (
            .O(N__36462),
            .I(N__36459));
    InMux I__4434 (
            .O(N__36459),
            .I(N__36456));
    LocalMux I__4433 (
            .O(N__36456),
            .I(N__36451));
    InMux I__4432 (
            .O(N__36455),
            .I(N__36446));
    InMux I__4431 (
            .O(N__36454),
            .I(N__36446));
    Odrv4 I__4430 (
            .O(N__36451),
            .I(drone_altitude_1));
    LocalMux I__4429 (
            .O(N__36446),
            .I(drone_altitude_1));
    InMux I__4428 (
            .O(N__36441),
            .I(N__36438));
    LocalMux I__4427 (
            .O(N__36438),
            .I(N__36435));
    Span4Mux_v I__4426 (
            .O(N__36435),
            .I(N__36432));
    Span4Mux_s1_h I__4425 (
            .O(N__36432),
            .I(N__36429));
    Odrv4 I__4424 (
            .O(N__36429),
            .I(\pid_alt.error_axbZ0Z_1 ));
    InMux I__4423 (
            .O(N__36426),
            .I(N__36420));
    InMux I__4422 (
            .O(N__36425),
            .I(N__36420));
    LocalMux I__4421 (
            .O(N__36420),
            .I(drone_H_disp_side_1));
    InMux I__4420 (
            .O(N__36417),
            .I(N__36412));
    InMux I__4419 (
            .O(N__36416),
            .I(N__36407));
    InMux I__4418 (
            .O(N__36415),
            .I(N__36407));
    LocalMux I__4417 (
            .O(N__36412),
            .I(drone_altitude_9));
    LocalMux I__4416 (
            .O(N__36407),
            .I(drone_altitude_9));
    InMux I__4415 (
            .O(N__36402),
            .I(N__36399));
    LocalMux I__4414 (
            .O(N__36399),
            .I(N__36396));
    Span4Mux_h I__4413 (
            .O(N__36396),
            .I(N__36393));
    Odrv4 I__4412 (
            .O(N__36393),
            .I(drone_altitude_i_9));
    InMux I__4411 (
            .O(N__36390),
            .I(N__36387));
    LocalMux I__4410 (
            .O(N__36387),
            .I(N__36384));
    Span4Mux_v I__4409 (
            .O(N__36384),
            .I(N__36381));
    Span4Mux_h I__4408 (
            .O(N__36381),
            .I(N__36378));
    Odrv4 I__4407 (
            .O(N__36378),
            .I(\pid_alt.O_5_5 ));
    InMux I__4406 (
            .O(N__36375),
            .I(N__36366));
    InMux I__4405 (
            .O(N__36374),
            .I(N__36366));
    InMux I__4404 (
            .O(N__36373),
            .I(N__36366));
    LocalMux I__4403 (
            .O(N__36366),
            .I(N__36363));
    Odrv4 I__4402 (
            .O(N__36363),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    InMux I__4401 (
            .O(N__36360),
            .I(N__36357));
    LocalMux I__4400 (
            .O(N__36357),
            .I(N__36354));
    Span4Mux_h I__4399 (
            .O(N__36354),
            .I(N__36351));
    Odrv4 I__4398 (
            .O(N__36351),
            .I(\pid_alt.O_5_7 ));
    InMux I__4397 (
            .O(N__36348),
            .I(N__36342));
    InMux I__4396 (
            .O(N__36347),
            .I(N__36342));
    LocalMux I__4395 (
            .O(N__36342),
            .I(N__36339));
    Odrv4 I__4394 (
            .O(N__36339),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__4393 (
            .O(N__36336),
            .I(N__36333));
    LocalMux I__4392 (
            .O(N__36333),
            .I(N__36330));
    Span4Mux_h I__4391 (
            .O(N__36330),
            .I(N__36327));
    Odrv4 I__4390 (
            .O(N__36327),
            .I(\pid_alt.O_5_6 ));
    InMux I__4389 (
            .O(N__36324),
            .I(N__36320));
    InMux I__4388 (
            .O(N__36323),
            .I(N__36317));
    LocalMux I__4387 (
            .O(N__36320),
            .I(N__36314));
    LocalMux I__4386 (
            .O(N__36317),
            .I(N__36311));
    Odrv12 I__4385 (
            .O(N__36314),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    Odrv4 I__4384 (
            .O(N__36311),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    InMux I__4383 (
            .O(N__36306),
            .I(N__36303));
    LocalMux I__4382 (
            .O(N__36303),
            .I(N__36300));
    Span4Mux_h I__4381 (
            .O(N__36300),
            .I(N__36297));
    Odrv4 I__4380 (
            .O(N__36297),
            .I(\pid_alt.O_5_13 ));
    InMux I__4379 (
            .O(N__36294),
            .I(N__36288));
    InMux I__4378 (
            .O(N__36293),
            .I(N__36288));
    LocalMux I__4377 (
            .O(N__36288),
            .I(N__36285));
    Odrv12 I__4376 (
            .O(N__36285),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    CEMux I__4375 (
            .O(N__36282),
            .I(N__36237));
    CEMux I__4374 (
            .O(N__36281),
            .I(N__36237));
    CEMux I__4373 (
            .O(N__36280),
            .I(N__36237));
    CEMux I__4372 (
            .O(N__36279),
            .I(N__36237));
    CEMux I__4371 (
            .O(N__36278),
            .I(N__36237));
    CEMux I__4370 (
            .O(N__36277),
            .I(N__36237));
    CEMux I__4369 (
            .O(N__36276),
            .I(N__36237));
    CEMux I__4368 (
            .O(N__36275),
            .I(N__36237));
    CEMux I__4367 (
            .O(N__36274),
            .I(N__36237));
    CEMux I__4366 (
            .O(N__36273),
            .I(N__36237));
    CEMux I__4365 (
            .O(N__36272),
            .I(N__36237));
    CEMux I__4364 (
            .O(N__36271),
            .I(N__36237));
    CEMux I__4363 (
            .O(N__36270),
            .I(N__36237));
    CEMux I__4362 (
            .O(N__36269),
            .I(N__36237));
    CEMux I__4361 (
            .O(N__36268),
            .I(N__36237));
    GlobalMux I__4360 (
            .O(N__36237),
            .I(N__36234));
    gio2CtrlBuf I__4359 (
            .O(N__36234),
            .I(\pid_alt.N_579_0_g ));
    CascadeMux I__4358 (
            .O(N__36231),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1_cascade_ ));
    InMux I__4357 (
            .O(N__36228),
            .I(N__36222));
    InMux I__4356 (
            .O(N__36227),
            .I(N__36222));
    LocalMux I__4355 (
            .O(N__36222),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ));
    InMux I__4354 (
            .O(N__36219),
            .I(N__36216));
    LocalMux I__4353 (
            .O(N__36216),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ));
    InMux I__4352 (
            .O(N__36213),
            .I(N__36201));
    InMux I__4351 (
            .O(N__36212),
            .I(N__36201));
    InMux I__4350 (
            .O(N__36211),
            .I(N__36201));
    InMux I__4349 (
            .O(N__36210),
            .I(N__36201));
    LocalMux I__4348 (
            .O(N__36201),
            .I(N__36198));
    Span12Mux_v I__4347 (
            .O(N__36198),
            .I(N__36195));
    Odrv12 I__4346 (
            .O(N__36195),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__4345 (
            .O(N__36192),
            .I(N__36187));
    InMux I__4344 (
            .O(N__36191),
            .I(N__36182));
    InMux I__4343 (
            .O(N__36190),
            .I(N__36182));
    LocalMux I__4342 (
            .O(N__36187),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__4341 (
            .O(N__36182),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__4340 (
            .O(N__36177),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ));
    InMux I__4339 (
            .O(N__36174),
            .I(N__36168));
    InMux I__4338 (
            .O(N__36173),
            .I(N__36168));
    LocalMux I__4337 (
            .O(N__36168),
            .I(N__36165));
    Odrv12 I__4336 (
            .O(N__36165),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ));
    InMux I__4335 (
            .O(N__36162),
            .I(N__36158));
    InMux I__4334 (
            .O(N__36161),
            .I(N__36154));
    LocalMux I__4333 (
            .O(N__36158),
            .I(N__36151));
    InMux I__4332 (
            .O(N__36157),
            .I(N__36148));
    LocalMux I__4331 (
            .O(N__36154),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    Odrv4 I__4330 (
            .O(N__36151),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    LocalMux I__4329 (
            .O(N__36148),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    CascadeMux I__4328 (
            .O(N__36141),
            .I(\pid_alt.un1_pid_prereg_16_0_cascade_ ));
    InMux I__4327 (
            .O(N__36138),
            .I(N__36134));
    CascadeMux I__4326 (
            .O(N__36137),
            .I(N__36131));
    LocalMux I__4325 (
            .O(N__36134),
            .I(N__36128));
    InMux I__4324 (
            .O(N__36131),
            .I(N__36124));
    Span4Mux_v I__4323 (
            .O(N__36128),
            .I(N__36121));
    InMux I__4322 (
            .O(N__36127),
            .I(N__36118));
    LocalMux I__4321 (
            .O(N__36124),
            .I(N__36115));
    Span4Mux_v I__4320 (
            .O(N__36121),
            .I(N__36112));
    LocalMux I__4319 (
            .O(N__36118),
            .I(N__36109));
    Span4Mux_h I__4318 (
            .O(N__36115),
            .I(N__36106));
    Odrv4 I__4317 (
            .O(N__36112),
            .I(\pid_alt.un2_pid_prereg_cry_1_c_RNIHS3R ));
    Odrv4 I__4316 (
            .O(N__36109),
            .I(\pid_alt.un2_pid_prereg_cry_1_c_RNIHS3R ));
    Odrv4 I__4315 (
            .O(N__36106),
            .I(\pid_alt.un2_pid_prereg_cry_1_c_RNIHS3R ));
    InMux I__4314 (
            .O(N__36099),
            .I(N__36096));
    LocalMux I__4313 (
            .O(N__36096),
            .I(N__36093));
    Sp12to4 I__4312 (
            .O(N__36093),
            .I(N__36090));
    Odrv12 I__4311 (
            .O(N__36090),
            .I(\pid_alt.error_d_reg_prev_esr_RNI32PN4Z0Z_1 ));
    InMux I__4310 (
            .O(N__36087),
            .I(N__36080));
    InMux I__4309 (
            .O(N__36086),
            .I(N__36080));
    InMux I__4308 (
            .O(N__36085),
            .I(N__36077));
    LocalMux I__4307 (
            .O(N__36080),
            .I(N__36074));
    LocalMux I__4306 (
            .O(N__36077),
            .I(N__36071));
    Span12Mux_s6_h I__4305 (
            .O(N__36074),
            .I(N__36068));
    Span12Mux_h I__4304 (
            .O(N__36071),
            .I(N__36065));
    Span12Mux_v I__4303 (
            .O(N__36068),
            .I(N__36062));
    Odrv12 I__4302 (
            .O(N__36065),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    Odrv12 I__4301 (
            .O(N__36062),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    InMux I__4300 (
            .O(N__36057),
            .I(N__36053));
    InMux I__4299 (
            .O(N__36056),
            .I(N__36050));
    LocalMux I__4298 (
            .O(N__36053),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__4297 (
            .O(N__36050),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    CascadeMux I__4296 (
            .O(N__36045),
            .I(N__36042));
    InMux I__4295 (
            .O(N__36042),
            .I(N__36039));
    LocalMux I__4294 (
            .O(N__36039),
            .I(N__36035));
    CascadeMux I__4293 (
            .O(N__36038),
            .I(N__36031));
    Span4Mux_v I__4292 (
            .O(N__36035),
            .I(N__36028));
    InMux I__4291 (
            .O(N__36034),
            .I(N__36025));
    InMux I__4290 (
            .O(N__36031),
            .I(N__36022));
    Span4Mux_v I__4289 (
            .O(N__36028),
            .I(N__36019));
    LocalMux I__4288 (
            .O(N__36025),
            .I(N__36016));
    LocalMux I__4287 (
            .O(N__36022),
            .I(N__36013));
    Sp12to4 I__4286 (
            .O(N__36019),
            .I(N__36010));
    Span4Mux_v I__4285 (
            .O(N__36016),
            .I(N__36005));
    Span4Mux_h I__4284 (
            .O(N__36013),
            .I(N__36005));
    Odrv12 I__4283 (
            .O(N__36010),
            .I(\pid_alt.un2_pid_prereg_cry_2_c_RNIK05R ));
    Odrv4 I__4282 (
            .O(N__36005),
            .I(\pid_alt.un2_pid_prereg_cry_2_c_RNIK05R ));
    InMux I__4281 (
            .O(N__36000),
            .I(N__35997));
    LocalMux I__4280 (
            .O(N__35997),
            .I(N__35994));
    Odrv12 I__4279 (
            .O(N__35994),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9F5Q6Z0Z_2 ));
    InMux I__4278 (
            .O(N__35991),
            .I(N__35988));
    LocalMux I__4277 (
            .O(N__35988),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ));
    CascadeMux I__4276 (
            .O(N__35985),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2_cascade_ ));
    InMux I__4275 (
            .O(N__35982),
            .I(N__35979));
    LocalMux I__4274 (
            .O(N__35979),
            .I(N__35975));
    InMux I__4273 (
            .O(N__35978),
            .I(N__35972));
    Sp12to4 I__4272 (
            .O(N__35975),
            .I(N__35967));
    LocalMux I__4271 (
            .O(N__35972),
            .I(N__35967));
    Odrv12 I__4270 (
            .O(N__35967),
            .I(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ));
    InMux I__4269 (
            .O(N__35964),
            .I(N__35958));
    InMux I__4268 (
            .O(N__35963),
            .I(N__35958));
    LocalMux I__4267 (
            .O(N__35958),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    InMux I__4266 (
            .O(N__35955),
            .I(N__35946));
    InMux I__4265 (
            .O(N__35954),
            .I(N__35946));
    InMux I__4264 (
            .O(N__35953),
            .I(N__35946));
    LocalMux I__4263 (
            .O(N__35946),
            .I(N__35943));
    Sp12to4 I__4262 (
            .O(N__35943),
            .I(N__35940));
    Span12Mux_v I__4261 (
            .O(N__35940),
            .I(N__35937));
    Odrv12 I__4260 (
            .O(N__35937),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    InMux I__4259 (
            .O(N__35934),
            .I(N__35928));
    InMux I__4258 (
            .O(N__35933),
            .I(N__35928));
    LocalMux I__4257 (
            .O(N__35928),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__4256 (
            .O(N__35925),
            .I(N__35919));
    InMux I__4255 (
            .O(N__35924),
            .I(N__35919));
    LocalMux I__4254 (
            .O(N__35919),
            .I(N__35916));
    Span4Mux_v I__4253 (
            .O(N__35916),
            .I(N__35913));
    Odrv4 I__4252 (
            .O(N__35913),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    CascadeMux I__4251 (
            .O(N__35910),
            .I(N__35906));
    CascadeMux I__4250 (
            .O(N__35909),
            .I(N__35903));
    InMux I__4249 (
            .O(N__35906),
            .I(N__35900));
    InMux I__4248 (
            .O(N__35903),
            .I(N__35897));
    LocalMux I__4247 (
            .O(N__35900),
            .I(N__35894));
    LocalMux I__4246 (
            .O(N__35897),
            .I(N__35891));
    Span4Mux_v I__4245 (
            .O(N__35894),
            .I(N__35888));
    Span4Mux_h I__4244 (
            .O(N__35891),
            .I(N__35885));
    Odrv4 I__4243 (
            .O(N__35888),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIKNU2Z0Z_6 ));
    Odrv4 I__4242 (
            .O(N__35885),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIKNU2Z0Z_6 ));
    InMux I__4241 (
            .O(N__35880),
            .I(N__35877));
    LocalMux I__4240 (
            .O(N__35877),
            .I(N__35874));
    Span4Mux_v I__4239 (
            .O(N__35874),
            .I(N__35871));
    Odrv4 I__4238 (
            .O(N__35871),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDJGT5Z0Z_7 ));
    InMux I__4237 (
            .O(N__35868),
            .I(N__35861));
    InMux I__4236 (
            .O(N__35867),
            .I(N__35861));
    InMux I__4235 (
            .O(N__35866),
            .I(N__35858));
    LocalMux I__4234 (
            .O(N__35861),
            .I(N__35855));
    LocalMux I__4233 (
            .O(N__35858),
            .I(N__35852));
    Span4Mux_v I__4232 (
            .O(N__35855),
            .I(N__35849));
    Odrv4 I__4231 (
            .O(N__35852),
            .I(\pid_alt.un2_pid_prereg_cry_7_c_RNIQMCS ));
    Odrv4 I__4230 (
            .O(N__35849),
            .I(\pid_alt.un2_pid_prereg_cry_7_c_RNIQMCS ));
    CascadeMux I__4229 (
            .O(N__35844),
            .I(N__35841));
    InMux I__4228 (
            .O(N__35841),
            .I(N__35835));
    InMux I__4227 (
            .O(N__35840),
            .I(N__35835));
    LocalMux I__4226 (
            .O(N__35835),
            .I(N__35832));
    Odrv4 I__4225 (
            .O(N__35832),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    InMux I__4224 (
            .O(N__35829),
            .I(N__35823));
    InMux I__4223 (
            .O(N__35828),
            .I(N__35823));
    LocalMux I__4222 (
            .O(N__35823),
            .I(N__35820));
    Odrv4 I__4221 (
            .O(N__35820),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    CascadeMux I__4220 (
            .O(N__35817),
            .I(N__35814));
    InMux I__4219 (
            .O(N__35814),
            .I(N__35811));
    LocalMux I__4218 (
            .O(N__35811),
            .I(N__35807));
    InMux I__4217 (
            .O(N__35810),
            .I(N__35804));
    Span4Mux_v I__4216 (
            .O(N__35807),
            .I(N__35801));
    LocalMux I__4215 (
            .O(N__35804),
            .I(\pid_alt.error_d_reg_prev_esr_RNIRUOU2Z0Z_7 ));
    Odrv4 I__4214 (
            .O(N__35801),
            .I(\pid_alt.error_d_reg_prev_esr_RNIRUOU2Z0Z_7 ));
    InMux I__4213 (
            .O(N__35796),
            .I(N__35790));
    InMux I__4212 (
            .O(N__35795),
            .I(N__35790));
    LocalMux I__4211 (
            .O(N__35790),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    InMux I__4210 (
            .O(N__35787),
            .I(N__35781));
    InMux I__4209 (
            .O(N__35786),
            .I(N__35781));
    LocalMux I__4208 (
            .O(N__35781),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__4207 (
            .O(N__35778),
            .I(N__35769));
    InMux I__4206 (
            .O(N__35777),
            .I(N__35769));
    InMux I__4205 (
            .O(N__35776),
            .I(N__35769));
    LocalMux I__4204 (
            .O(N__35769),
            .I(N__35766));
    Span4Mux_v I__4203 (
            .O(N__35766),
            .I(N__35763));
    Span4Mux_v I__4202 (
            .O(N__35763),
            .I(N__35760));
    Span4Mux_h I__4201 (
            .O(N__35760),
            .I(N__35757));
    Odrv4 I__4200 (
            .O(N__35757),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    InMux I__4199 (
            .O(N__35754),
            .I(N__35748));
    InMux I__4198 (
            .O(N__35753),
            .I(N__35748));
    LocalMux I__4197 (
            .O(N__35748),
            .I(N__35745));
    Odrv4 I__4196 (
            .O(N__35745),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    InMux I__4195 (
            .O(N__35742),
            .I(N__35738));
    InMux I__4194 (
            .O(N__35741),
            .I(N__35735));
    LocalMux I__4193 (
            .O(N__35738),
            .I(N__35732));
    LocalMux I__4192 (
            .O(N__35735),
            .I(N__35729));
    Span4Mux_h I__4191 (
            .O(N__35732),
            .I(N__35726));
    Span4Mux_h I__4190 (
            .O(N__35729),
            .I(N__35721));
    Span4Mux_v I__4189 (
            .O(N__35726),
            .I(N__35721));
    Span4Mux_v I__4188 (
            .O(N__35721),
            .I(N__35718));
    Odrv4 I__4187 (
            .O(N__35718),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__4186 (
            .O(N__35715),
            .I(N__35709));
    InMux I__4185 (
            .O(N__35714),
            .I(N__35709));
    LocalMux I__4184 (
            .O(N__35709),
            .I(N__35705));
    InMux I__4183 (
            .O(N__35708),
            .I(N__35702));
    Span4Mux_v I__4182 (
            .O(N__35705),
            .I(N__35697));
    LocalMux I__4181 (
            .O(N__35702),
            .I(N__35697));
    Span4Mux_h I__4180 (
            .O(N__35697),
            .I(N__35694));
    Span4Mux_v I__4179 (
            .O(N__35694),
            .I(N__35691));
    Odrv4 I__4178 (
            .O(N__35691),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__4177 (
            .O(N__35688),
            .I(N__35685));
    LocalMux I__4176 (
            .O(N__35685),
            .I(N__35681));
    InMux I__4175 (
            .O(N__35684),
            .I(N__35678));
    Span4Mux_h I__4174 (
            .O(N__35681),
            .I(N__35675));
    LocalMux I__4173 (
            .O(N__35678),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__4172 (
            .O(N__35675),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__4171 (
            .O(N__35670),
            .I(N__35666));
    InMux I__4170 (
            .O(N__35669),
            .I(N__35663));
    LocalMux I__4169 (
            .O(N__35666),
            .I(N__35660));
    LocalMux I__4168 (
            .O(N__35663),
            .I(N__35657));
    Span4Mux_v I__4167 (
            .O(N__35660),
            .I(N__35652));
    Span4Mux_v I__4166 (
            .O(N__35657),
            .I(N__35652));
    Span4Mux_v I__4165 (
            .O(N__35652),
            .I(N__35649));
    Odrv4 I__4164 (
            .O(N__35649),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    InMux I__4163 (
            .O(N__35646),
            .I(N__35640));
    InMux I__4162 (
            .O(N__35645),
            .I(N__35640));
    LocalMux I__4161 (
            .O(N__35640),
            .I(N__35637));
    Span4Mux_h I__4160 (
            .O(N__35637),
            .I(N__35634));
    Odrv4 I__4159 (
            .O(N__35634),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    InMux I__4158 (
            .O(N__35631),
            .I(N__35624));
    InMux I__4157 (
            .O(N__35630),
            .I(N__35624));
    InMux I__4156 (
            .O(N__35629),
            .I(N__35621));
    LocalMux I__4155 (
            .O(N__35624),
            .I(N__35616));
    LocalMux I__4154 (
            .O(N__35621),
            .I(N__35616));
    Span4Mux_v I__4153 (
            .O(N__35616),
            .I(N__35613));
    Span4Mux_v I__4152 (
            .O(N__35613),
            .I(N__35610));
    Span4Mux_v I__4151 (
            .O(N__35610),
            .I(N__35607));
    Odrv4 I__4150 (
            .O(N__35607),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    InMux I__4149 (
            .O(N__35604),
            .I(N__35600));
    InMux I__4148 (
            .O(N__35603),
            .I(N__35597));
    LocalMux I__4147 (
            .O(N__35600),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    LocalMux I__4146 (
            .O(N__35597),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    CascadeMux I__4145 (
            .O(N__35592),
            .I(N__35589));
    InMux I__4144 (
            .O(N__35589),
            .I(N__35585));
    InMux I__4143 (
            .O(N__35588),
            .I(N__35582));
    LocalMux I__4142 (
            .O(N__35585),
            .I(N__35579));
    LocalMux I__4141 (
            .O(N__35582),
            .I(N__35576));
    Span4Mux_h I__4140 (
            .O(N__35579),
            .I(N__35573));
    Odrv4 I__4139 (
            .O(N__35576),
            .I(\pid_alt.error_d_reg_prev_esr_RNI06021Z0Z_20 ));
    Odrv4 I__4138 (
            .O(N__35573),
            .I(\pid_alt.error_d_reg_prev_esr_RNI06021Z0Z_20 ));
    CascadeMux I__4137 (
            .O(N__35568),
            .I(N__35565));
    InMux I__4136 (
            .O(N__35565),
            .I(N__35562));
    LocalMux I__4135 (
            .O(N__35562),
            .I(N__35559));
    Odrv4 I__4134 (
            .O(N__35559),
            .I(\pid_alt.error_d_reg_prev_esr_RNI06021_2Z0Z_20 ));
    InMux I__4133 (
            .O(N__35556),
            .I(bfn_4_14_0_));
    InMux I__4132 (
            .O(N__35553),
            .I(N__35550));
    LocalMux I__4131 (
            .O(N__35550),
            .I(N__35547));
    Span4Mux_h I__4130 (
            .O(N__35547),
            .I(N__35544));
    Odrv4 I__4129 (
            .O(N__35544),
            .I(\pid_alt.un1_pid_prereg_0_axb_24 ));
    InMux I__4128 (
            .O(N__35541),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    CascadeMux I__4127 (
            .O(N__35538),
            .I(N__35533));
    InMux I__4126 (
            .O(N__35537),
            .I(N__35530));
    InMux I__4125 (
            .O(N__35536),
            .I(N__35527));
    InMux I__4124 (
            .O(N__35533),
            .I(N__35524));
    LocalMux I__4123 (
            .O(N__35530),
            .I(N__35521));
    LocalMux I__4122 (
            .O(N__35527),
            .I(N__35516));
    LocalMux I__4121 (
            .O(N__35524),
            .I(N__35516));
    Span4Mux_v I__4120 (
            .O(N__35521),
            .I(N__35511));
    Span4Mux_v I__4119 (
            .O(N__35516),
            .I(N__35511));
    Odrv4 I__4118 (
            .O(N__35511),
            .I(\pid_alt.un2_pid_prereg_cry_0_c_RNIEO2R ));
    CascadeMux I__4117 (
            .O(N__35508),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ));
    InMux I__4116 (
            .O(N__35505),
            .I(N__35502));
    LocalMux I__4115 (
            .O(N__35502),
            .I(N__35499));
    Odrv12 I__4114 (
            .O(N__35499),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3RCL2Z0Z_1 ));
    InMux I__4113 (
            .O(N__35496),
            .I(N__35493));
    LocalMux I__4112 (
            .O(N__35493),
            .I(N__35490));
    Span12Mux_h I__4111 (
            .O(N__35490),
            .I(N__35487));
    Odrv12 I__4110 (
            .O(N__35487),
            .I(\pid_alt.O_5_4 ));
    InMux I__4109 (
            .O(N__35484),
            .I(N__35481));
    LocalMux I__4108 (
            .O(N__35481),
            .I(N__35477));
    CascadeMux I__4107 (
            .O(N__35480),
            .I(N__35474));
    Span4Mux_v I__4106 (
            .O(N__35477),
            .I(N__35471));
    InMux I__4105 (
            .O(N__35474),
            .I(N__35468));
    Span4Mux_v I__4104 (
            .O(N__35471),
            .I(N__35465));
    LocalMux I__4103 (
            .O(N__35468),
            .I(N__35462));
    Span4Mux_h I__4102 (
            .O(N__35465),
            .I(N__35457));
    Span4Mux_v I__4101 (
            .O(N__35462),
            .I(N__35457));
    Odrv4 I__4100 (
            .O(N__35457),
            .I(\pid_alt.un1_pid_prereg_0 ));
    InMux I__4099 (
            .O(N__35454),
            .I(N__35448));
    InMux I__4098 (
            .O(N__35453),
            .I(N__35448));
    LocalMux I__4097 (
            .O(N__35448),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__4096 (
            .O(N__35445),
            .I(N__35442));
    LocalMux I__4095 (
            .O(N__35442),
            .I(N__35439));
    Span4Mux_v I__4094 (
            .O(N__35439),
            .I(N__35436));
    Odrv4 I__4093 (
            .O(N__35436),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    InMux I__4092 (
            .O(N__35433),
            .I(N__35430));
    LocalMux I__4091 (
            .O(N__35430),
            .I(N__35427));
    Span4Mux_v I__4090 (
            .O(N__35427),
            .I(N__35424));
    Span4Mux_h I__4089 (
            .O(N__35424),
            .I(N__35421));
    Span4Mux_v I__4088 (
            .O(N__35421),
            .I(N__35418));
    Odrv4 I__4087 (
            .O(N__35418),
            .I(\pid_alt.O_3_4 ));
    InMux I__4086 (
            .O(N__35415),
            .I(N__35412));
    LocalMux I__4085 (
            .O(N__35412),
            .I(N__35409));
    Span4Mux_v I__4084 (
            .O(N__35409),
            .I(N__35404));
    InMux I__4083 (
            .O(N__35408),
            .I(N__35399));
    InMux I__4082 (
            .O(N__35407),
            .I(N__35399));
    Odrv4 I__4081 (
            .O(N__35404),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    LocalMux I__4080 (
            .O(N__35399),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    InMux I__4079 (
            .O(N__35394),
            .I(N__35390));
    InMux I__4078 (
            .O(N__35393),
            .I(N__35387));
    LocalMux I__4077 (
            .O(N__35390),
            .I(N__35384));
    LocalMux I__4076 (
            .O(N__35387),
            .I(N__35381));
    Span4Mux_v I__4075 (
            .O(N__35384),
            .I(N__35376));
    Span4Mux_v I__4074 (
            .O(N__35381),
            .I(N__35376));
    Span4Mux_v I__4073 (
            .O(N__35376),
            .I(N__35373));
    Odrv4 I__4072 (
            .O(N__35373),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    InMux I__4071 (
            .O(N__35370),
            .I(N__35366));
    InMux I__4070 (
            .O(N__35369),
            .I(N__35363));
    LocalMux I__4069 (
            .O(N__35366),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    LocalMux I__4068 (
            .O(N__35363),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__4067 (
            .O(N__35358),
            .I(N__35351));
    InMux I__4066 (
            .O(N__35357),
            .I(N__35351));
    InMux I__4065 (
            .O(N__35356),
            .I(N__35348));
    LocalMux I__4064 (
            .O(N__35351),
            .I(N__35343));
    LocalMux I__4063 (
            .O(N__35348),
            .I(N__35343));
    Span4Mux_h I__4062 (
            .O(N__35343),
            .I(N__35340));
    Span4Mux_v I__4061 (
            .O(N__35340),
            .I(N__35337));
    Span4Mux_v I__4060 (
            .O(N__35337),
            .I(N__35334));
    Odrv4 I__4059 (
            .O(N__35334),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    InMux I__4058 (
            .O(N__35331),
            .I(N__35328));
    LocalMux I__4057 (
            .O(N__35328),
            .I(N__35324));
    InMux I__4056 (
            .O(N__35327),
            .I(N__35321));
    Span4Mux_h I__4055 (
            .O(N__35324),
            .I(N__35318));
    LocalMux I__4054 (
            .O(N__35321),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    Odrv4 I__4053 (
            .O(N__35318),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__4052 (
            .O(N__35313),
            .I(bfn_4_13_0_));
    InMux I__4051 (
            .O(N__35310),
            .I(N__35307));
    LocalMux I__4050 (
            .O(N__35307),
            .I(N__35304));
    Span4Mux_h I__4049 (
            .O(N__35304),
            .I(N__35301));
    Odrv4 I__4048 (
            .O(N__35301),
            .I(\pid_alt.error_d_reg_prev_esr_RNI060F3Z0Z_15 ));
    InMux I__4047 (
            .O(N__35298),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__4046 (
            .O(N__35295),
            .I(N__35292));
    LocalMux I__4045 (
            .O(N__35292),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGO2F3Z0Z_16 ));
    CascadeMux I__4044 (
            .O(N__35289),
            .I(N__35286));
    InMux I__4043 (
            .O(N__35286),
            .I(N__35282));
    InMux I__4042 (
            .O(N__35285),
            .I(N__35279));
    LocalMux I__4041 (
            .O(N__35282),
            .I(N__35276));
    LocalMux I__4040 (
            .O(N__35279),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKNGN1Z0Z_15 ));
    Odrv4 I__4039 (
            .O(N__35276),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKNGN1Z0Z_15 ));
    InMux I__4038 (
            .O(N__35271),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__4037 (
            .O(N__35268),
            .I(N__35265));
    LocalMux I__4036 (
            .O(N__35265),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0B5F3Z0Z_17 ));
    CascadeMux I__4035 (
            .O(N__35262),
            .I(N__35258));
    CascadeMux I__4034 (
            .O(N__35261),
            .I(N__35255));
    InMux I__4033 (
            .O(N__35258),
            .I(N__35252));
    InMux I__4032 (
            .O(N__35255),
            .I(N__35249));
    LocalMux I__4031 (
            .O(N__35252),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0IN1Z0Z_16 ));
    LocalMux I__4030 (
            .O(N__35249),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0IN1Z0Z_16 ));
    InMux I__4029 (
            .O(N__35244),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__4028 (
            .O(N__35241),
            .I(N__35238));
    LocalMux I__4027 (
            .O(N__35238),
            .I(N__35235));
    Odrv4 I__4026 (
            .O(N__35235),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGT7F3Z0Z_18 ));
    InMux I__4025 (
            .O(N__35232),
            .I(N__35228));
    CascadeMux I__4024 (
            .O(N__35231),
            .I(N__35225));
    LocalMux I__4023 (
            .O(N__35228),
            .I(N__35222));
    InMux I__4022 (
            .O(N__35225),
            .I(N__35219));
    Odrv4 I__4021 (
            .O(N__35222),
            .I(\pid_alt.error_d_reg_prev_esr_RNI4AJN1Z0Z_17 ));
    LocalMux I__4020 (
            .O(N__35219),
            .I(\pid_alt.error_d_reg_prev_esr_RNI4AJN1Z0Z_17 ));
    InMux I__4019 (
            .O(N__35214),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__4018 (
            .O(N__35211),
            .I(N__35208));
    LocalMux I__4017 (
            .O(N__35208),
            .I(N__35205));
    Span4Mux_h I__4016 (
            .O(N__35205),
            .I(N__35202));
    Odrv4 I__4015 (
            .O(N__35202),
            .I(\pid_alt.error_d_reg_prev_esr_RNISEDF3Z0Z_19 ));
    InMux I__4014 (
            .O(N__35199),
            .I(N__35195));
    CascadeMux I__4013 (
            .O(N__35198),
            .I(N__35192));
    LocalMux I__4012 (
            .O(N__35195),
            .I(N__35189));
    InMux I__4011 (
            .O(N__35192),
            .I(N__35186));
    Span4Mux_v I__4010 (
            .O(N__35189),
            .I(N__35183));
    LocalMux I__4009 (
            .O(N__35186),
            .I(N__35180));
    Odrv4 I__4008 (
            .O(N__35183),
            .I(\pid_alt.error_d_reg_prev_esr_RNICJKN1Z0Z_18 ));
    Odrv4 I__4007 (
            .O(N__35180),
            .I(\pid_alt.error_d_reg_prev_esr_RNICJKN1Z0Z_18 ));
    InMux I__4006 (
            .O(N__35175),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__4005 (
            .O(N__35172),
            .I(N__35169));
    LocalMux I__4004 (
            .O(N__35169),
            .I(N__35166));
    Span4Mux_v I__4003 (
            .O(N__35166),
            .I(N__35163));
    Odrv4 I__4002 (
            .O(N__35163),
            .I(\pid_alt.error_d_reg_prev_esr_RNI06021_0Z0Z_20 ));
    CascadeMux I__4001 (
            .O(N__35160),
            .I(N__35157));
    InMux I__4000 (
            .O(N__35157),
            .I(N__35154));
    LocalMux I__3999 (
            .O(N__35154),
            .I(N__35151));
    Span4Mux_h I__3998 (
            .O(N__35151),
            .I(N__35148));
    Odrv4 I__3997 (
            .O(N__35148),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGRON1Z0Z_19 ));
    InMux I__3996 (
            .O(N__35145),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__3995 (
            .O(N__35142),
            .I(N__35139));
    LocalMux I__3994 (
            .O(N__35139),
            .I(N__35136));
    Span4Mux_h I__3993 (
            .O(N__35136),
            .I(N__35133));
    Odrv4 I__3992 (
            .O(N__35133),
            .I(\pid_alt.error_d_reg_prev_esr_RNI06021_1Z0Z_20 ));
    InMux I__3991 (
            .O(N__35130),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    InMux I__3990 (
            .O(N__35127),
            .I(N__35124));
    LocalMux I__3989 (
            .O(N__35124),
            .I(N__35121));
    Span4Mux_h I__3988 (
            .O(N__35121),
            .I(N__35118));
    Odrv4 I__3987 (
            .O(N__35118),
            .I(\pid_alt.error_d_reg_prev_esr_RNIRUDT5Z0Z_6 ));
    CascadeMux I__3986 (
            .O(N__35115),
            .I(N__35112));
    InMux I__3985 (
            .O(N__35112),
            .I(N__35108));
    InMux I__3984 (
            .O(N__35111),
            .I(N__35105));
    LocalMux I__3983 (
            .O(N__35108),
            .I(N__35102));
    LocalMux I__3982 (
            .O(N__35105),
            .I(N__35097));
    Span4Mux_v I__3981 (
            .O(N__35102),
            .I(N__35097));
    Odrv4 I__3980 (
            .O(N__35097),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9AMU2Z0Z_5 ));
    InMux I__3979 (
            .O(N__35094),
            .I(bfn_4_12_0_));
    InMux I__3978 (
            .O(N__35091),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__3977 (
            .O(N__35088),
            .I(N__35085));
    LocalMux I__3976 (
            .O(N__35085),
            .I(N__35082));
    Span4Mux_h I__3975 (
            .O(N__35082),
            .I(N__35079));
    Odrv4 I__3974 (
            .O(N__35079),
            .I(\pid_alt.error_d_reg_prev_esr_RNIV7JT5Z0Z_8 ));
    InMux I__3973 (
            .O(N__35076),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    InMux I__3972 (
            .O(N__35073),
            .I(N__35070));
    LocalMux I__3971 (
            .O(N__35070),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKLA75Z0Z_9 ));
    CascadeMux I__3970 (
            .O(N__35067),
            .I(N__35063));
    InMux I__3969 (
            .O(N__35066),
            .I(N__35060));
    InMux I__3968 (
            .O(N__35063),
            .I(N__35057));
    LocalMux I__3967 (
            .O(N__35060),
            .I(N__35052));
    LocalMux I__3966 (
            .O(N__35057),
            .I(N__35052));
    Span4Mux_v I__3965 (
            .O(N__35052),
            .I(N__35049));
    Odrv4 I__3964 (
            .O(N__35049),
            .I(\pid_alt.error_d_reg_prev_esr_RNI49QU2Z0Z_8 ));
    InMux I__3963 (
            .O(N__35046),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__3962 (
            .O(N__35043),
            .I(N__35040));
    LocalMux I__3961 (
            .O(N__35040),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5H064Z0Z_10 ));
    CascadeMux I__3960 (
            .O(N__35037),
            .I(N__35033));
    CascadeMux I__3959 (
            .O(N__35036),
            .I(N__35030));
    InMux I__3958 (
            .O(N__35033),
            .I(N__35027));
    InMux I__3957 (
            .O(N__35030),
            .I(N__35024));
    LocalMux I__3956 (
            .O(N__35027),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGCG82Z0Z_9 ));
    LocalMux I__3955 (
            .O(N__35024),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGCG82Z0Z_9 ));
    InMux I__3954 (
            .O(N__35019),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__3953 (
            .O(N__35016),
            .I(N__35012));
    InMux I__3952 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__3951 (
            .O(N__35012),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL4GT1Z0Z_10 ));
    LocalMux I__3950 (
            .O(N__35009),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL4GT1Z0Z_10 ));
    CascadeMux I__3949 (
            .O(N__35004),
            .I(N__35001));
    InMux I__3948 (
            .O(N__35001),
            .I(N__34998));
    LocalMux I__3947 (
            .O(N__34998),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJJ1R3Z0Z_11 ));
    InMux I__3946 (
            .O(N__34995),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__3945 (
            .O(N__34992),
            .I(N__34989));
    LocalMux I__3944 (
            .O(N__34989),
            .I(\pid_alt.error_d_reg_prev_esr_RNIEF0O3Z0Z_12 ));
    CascadeMux I__3943 (
            .O(N__34986),
            .I(N__34982));
    CascadeMux I__3942 (
            .O(N__34985),
            .I(N__34979));
    InMux I__3941 (
            .O(N__34982),
            .I(N__34976));
    InMux I__3940 (
            .O(N__34979),
            .I(N__34973));
    LocalMux I__3939 (
            .O(N__34976),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUEHT1Z0Z_11 ));
    LocalMux I__3938 (
            .O(N__34973),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUEHT1Z0Z_11 ));
    InMux I__3937 (
            .O(N__34968),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__3936 (
            .O(N__34965),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    CascadeMux I__3935 (
            .O(N__34962),
            .I(\pid_alt.un1_reset_1_cascade_ ));
    InMux I__3934 (
            .O(N__34959),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__3933 (
            .O(N__34956),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__3932 (
            .O(N__34953),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    InMux I__3931 (
            .O(N__34950),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    CascadeMux I__3930 (
            .O(N__34947),
            .I(N__34944));
    InMux I__3929 (
            .O(N__34944),
            .I(N__34941));
    LocalMux I__3928 (
            .O(N__34941),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL2IS8Z0Z_3 ));
    InMux I__3927 (
            .O(N__34938),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__3926 (
            .O(N__34935),
            .I(N__34932));
    LocalMux I__3925 (
            .O(N__34932),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0K6S5Z0Z_4 ));
    CascadeMux I__3924 (
            .O(N__34929),
            .I(N__34925));
    CascadeMux I__3923 (
            .O(N__34928),
            .I(N__34922));
    InMux I__3922 (
            .O(N__34925),
            .I(N__34919));
    InMux I__3921 (
            .O(N__34922),
            .I(N__34916));
    LocalMux I__3920 (
            .O(N__34919),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0KHT2Z0Z_3 ));
    LocalMux I__3919 (
            .O(N__34916),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0KHT2Z0Z_3 ));
    InMux I__3918 (
            .O(N__34911),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__3917 (
            .O(N__34908),
            .I(N__34905));
    LocalMux I__3916 (
            .O(N__34905),
            .I(N__34902));
    Span4Mux_h I__3915 (
            .O(N__34902),
            .I(N__34899));
    Odrv4 I__3914 (
            .O(N__34899),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9ABT5Z0Z_5 ));
    InMux I__3913 (
            .O(N__34896),
            .I(N__34893));
    LocalMux I__3912 (
            .O(N__34893),
            .I(N__34889));
    CascadeMux I__3911 (
            .O(N__34892),
            .I(N__34886));
    Span4Mux_v I__3910 (
            .O(N__34889),
            .I(N__34883));
    InMux I__3909 (
            .O(N__34886),
            .I(N__34880));
    Odrv4 I__3908 (
            .O(N__34883),
            .I(\pid_alt.error_d_reg_prev_esr_RNI00LU2Z0Z_4 ));
    LocalMux I__3907 (
            .O(N__34880),
            .I(\pid_alt.error_d_reg_prev_esr_RNI00LU2Z0Z_4 ));
    InMux I__3906 (
            .O(N__34875),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__3905 (
            .O(N__34872),
            .I(N__34869));
    LocalMux I__3904 (
            .O(N__34869),
            .I(N__34865));
    InMux I__3903 (
            .O(N__34868),
            .I(N__34862));
    Odrv4 I__3902 (
            .O(N__34865),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    LocalMux I__3901 (
            .O(N__34862),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    InMux I__3900 (
            .O(N__34857),
            .I(N__34854));
    LocalMux I__3899 (
            .O(N__34854),
            .I(N__34850));
    InMux I__3898 (
            .O(N__34853),
            .I(N__34847));
    Odrv4 I__3897 (
            .O(N__34850),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__3896 (
            .O(N__34847),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    InMux I__3895 (
            .O(N__34842),
            .I(N__34837));
    InMux I__3894 (
            .O(N__34841),
            .I(N__34834));
    InMux I__3893 (
            .O(N__34840),
            .I(N__34831));
    LocalMux I__3892 (
            .O(N__34837),
            .I(N__34828));
    LocalMux I__3891 (
            .O(N__34834),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__3890 (
            .O(N__34831),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__3889 (
            .O(N__34828),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    CascadeMux I__3888 (
            .O(N__34821),
            .I(\pid_alt.m21_e_0_cascade_ ));
    InMux I__3887 (
            .O(N__34818),
            .I(N__34814));
    InMux I__3886 (
            .O(N__34817),
            .I(N__34811));
    LocalMux I__3885 (
            .O(N__34814),
            .I(N__34806));
    LocalMux I__3884 (
            .O(N__34811),
            .I(N__34806));
    Span4Mux_v I__3883 (
            .O(N__34806),
            .I(N__34802));
    InMux I__3882 (
            .O(N__34805),
            .I(N__34799));
    Odrv4 I__3881 (
            .O(N__34802),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__3880 (
            .O(N__34799),
            .I(\pid_alt.N_9_0 ));
    CascadeMux I__3879 (
            .O(N__34794),
            .I(N__34791));
    InMux I__3878 (
            .O(N__34791),
            .I(N__34788));
    LocalMux I__3877 (
            .O(N__34788),
            .I(\pid_alt.m21_e_9 ));
    InMux I__3876 (
            .O(N__34785),
            .I(N__34782));
    LocalMux I__3875 (
            .O(N__34782),
            .I(\pid_alt.m21_e_10 ));
    CascadeMux I__3874 (
            .O(N__34779),
            .I(\pid_alt.N_117_cascade_ ));
    CascadeMux I__3873 (
            .O(N__34776),
            .I(\pid_alt.un1_reset_1_0_i_cascade_ ));
    InMux I__3872 (
            .O(N__34773),
            .I(N__34769));
    InMux I__3871 (
            .O(N__34772),
            .I(N__34766));
    LocalMux I__3870 (
            .O(N__34769),
            .I(N__34760));
    LocalMux I__3869 (
            .O(N__34766),
            .I(N__34760));
    InMux I__3868 (
            .O(N__34765),
            .I(N__34756));
    Span4Mux_h I__3867 (
            .O(N__34760),
            .I(N__34753));
    InMux I__3866 (
            .O(N__34759),
            .I(N__34750));
    LocalMux I__3865 (
            .O(N__34756),
            .I(N__34747));
    Odrv4 I__3864 (
            .O(N__34753),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__3863 (
            .O(N__34750),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__3862 (
            .O(N__34747),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__3861 (
            .O(N__34740),
            .I(N__34736));
    InMux I__3860 (
            .O(N__34739),
            .I(N__34732));
    LocalMux I__3859 (
            .O(N__34736),
            .I(N__34729));
    InMux I__3858 (
            .O(N__34735),
            .I(N__34726));
    LocalMux I__3857 (
            .O(N__34732),
            .I(\pid_alt.error_i_acumm7lto13 ));
    Odrv4 I__3856 (
            .O(N__34729),
            .I(\pid_alt.error_i_acumm7lto13 ));
    LocalMux I__3855 (
            .O(N__34726),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__3854 (
            .O(N__34719),
            .I(N__34716));
    LocalMux I__3853 (
            .O(N__34716),
            .I(N__34712));
    InMux I__3852 (
            .O(N__34715),
            .I(N__34709));
    Odrv4 I__3851 (
            .O(N__34712),
            .I(\pid_alt.N_222 ));
    LocalMux I__3850 (
            .O(N__34709),
            .I(\pid_alt.N_222 ));
    InMux I__3849 (
            .O(N__34704),
            .I(N__34701));
    LocalMux I__3848 (
            .O(N__34701),
            .I(N__34698));
    Span4Mux_h I__3847 (
            .O(N__34698),
            .I(N__34695));
    Odrv4 I__3846 (
            .O(N__34695),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    InMux I__3845 (
            .O(N__34692),
            .I(N__34689));
    LocalMux I__3844 (
            .O(N__34689),
            .I(\pid_alt.drone_altitude_i_15 ));
    InMux I__3843 (
            .O(N__34686),
            .I(N__34683));
    LocalMux I__3842 (
            .O(N__34683),
            .I(N__34680));
    Odrv4 I__3841 (
            .O(N__34680),
            .I(\pid_alt.error_i_acumm_prereg15lt7 ));
    InMux I__3840 (
            .O(N__34677),
            .I(N__34674));
    LocalMux I__3839 (
            .O(N__34674),
            .I(\pid_alt.error_i_acumm_prereg15lto7Z0Z_2 ));
    InMux I__3838 (
            .O(N__34671),
            .I(bfn_3_19_0_));
    InMux I__3837 (
            .O(N__34668),
            .I(N__34665));
    LocalMux I__3836 (
            .O(N__34665),
            .I(\pid_alt.error_i_acumm_prereg_1_sqmuxa ));
    CEMux I__3835 (
            .O(N__34662),
            .I(N__34659));
    LocalMux I__3834 (
            .O(N__34659),
            .I(N__34654));
    CEMux I__3833 (
            .O(N__34658),
            .I(N__34651));
    CEMux I__3832 (
            .O(N__34657),
            .I(N__34648));
    Span4Mux_v I__3831 (
            .O(N__34654),
            .I(N__34644));
    LocalMux I__3830 (
            .O(N__34651),
            .I(N__34641));
    LocalMux I__3829 (
            .O(N__34648),
            .I(N__34638));
    CEMux I__3828 (
            .O(N__34647),
            .I(N__34635));
    Span4Mux_v I__3827 (
            .O(N__34644),
            .I(N__34632));
    Span4Mux_s3_h I__3826 (
            .O(N__34641),
            .I(N__34625));
    Span4Mux_v I__3825 (
            .O(N__34638),
            .I(N__34625));
    LocalMux I__3824 (
            .O(N__34635),
            .I(N__34625));
    Span4Mux_s3_h I__3823 (
            .O(N__34632),
            .I(N__34620));
    Span4Mux_v I__3822 (
            .O(N__34625),
            .I(N__34620));
    Span4Mux_v I__3821 (
            .O(N__34620),
            .I(N__34617));
    Odrv4 I__3820 (
            .O(N__34617),
            .I(\pid_alt.error_i_acumm_prereg_1_sqmuxa_0 ));
    CEMux I__3819 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__3818 (
            .O(N__34611),
            .I(\pid_alt.state_1_0_0 ));
    InMux I__3817 (
            .O(N__34608),
            .I(N__34605));
    LocalMux I__3816 (
            .O(N__34605),
            .I(N__34602));
    Span4Mux_h I__3815 (
            .O(N__34602),
            .I(N__34599));
    Odrv4 I__3814 (
            .O(N__34599),
            .I(\pid_alt.O_5_12 ));
    InMux I__3813 (
            .O(N__34596),
            .I(N__34592));
    InMux I__3812 (
            .O(N__34595),
            .I(N__34589));
    LocalMux I__3811 (
            .O(N__34592),
            .I(N__34586));
    LocalMux I__3810 (
            .O(N__34589),
            .I(N__34583));
    Span4Mux_h I__3809 (
            .O(N__34586),
            .I(N__34580));
    Span4Mux_v I__3808 (
            .O(N__34583),
            .I(N__34575));
    Span4Mux_v I__3807 (
            .O(N__34580),
            .I(N__34575));
    Odrv4 I__3806 (
            .O(N__34575),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__3805 (
            .O(N__34572),
            .I(N__34569));
    LocalMux I__3804 (
            .O(N__34569),
            .I(N__34566));
    Span4Mux_h I__3803 (
            .O(N__34566),
            .I(N__34563));
    Odrv4 I__3802 (
            .O(N__34563),
            .I(\pid_alt.O_5_11 ));
    InMux I__3801 (
            .O(N__34560),
            .I(N__34557));
    LocalMux I__3800 (
            .O(N__34557),
            .I(N__34554));
    Span4Mux_h I__3799 (
            .O(N__34554),
            .I(N__34551));
    Odrv4 I__3798 (
            .O(N__34551),
            .I(\pid_alt.O_3_5 ));
    CascadeMux I__3797 (
            .O(N__34548),
            .I(N__34544));
    CascadeMux I__3796 (
            .O(N__34547),
            .I(N__34541));
    InMux I__3795 (
            .O(N__34544),
            .I(N__34538));
    InMux I__3794 (
            .O(N__34541),
            .I(N__34534));
    LocalMux I__3793 (
            .O(N__34538),
            .I(N__34531));
    InMux I__3792 (
            .O(N__34537),
            .I(N__34528));
    LocalMux I__3791 (
            .O(N__34534),
            .I(alt_command_3));
    Odrv4 I__3790 (
            .O(N__34531),
            .I(alt_command_3));
    LocalMux I__3789 (
            .O(N__34528),
            .I(alt_command_3));
    CascadeMux I__3788 (
            .O(N__34521),
            .I(N__34518));
    InMux I__3787 (
            .O(N__34518),
            .I(N__34515));
    LocalMux I__3786 (
            .O(N__34515),
            .I(\pid_alt.alt_command_i_3 ));
    InMux I__3785 (
            .O(N__34512),
            .I(N__34509));
    LocalMux I__3784 (
            .O(N__34509),
            .I(N__34504));
    InMux I__3783 (
            .O(N__34508),
            .I(N__34499));
    InMux I__3782 (
            .O(N__34507),
            .I(N__34499));
    Odrv4 I__3781 (
            .O(N__34504),
            .I(drone_altitude_8));
    LocalMux I__3780 (
            .O(N__34499),
            .I(drone_altitude_8));
    InMux I__3779 (
            .O(N__34494),
            .I(N__34490));
    InMux I__3778 (
            .O(N__34493),
            .I(N__34486));
    LocalMux I__3777 (
            .O(N__34490),
            .I(N__34483));
    InMux I__3776 (
            .O(N__34489),
            .I(N__34480));
    LocalMux I__3775 (
            .O(N__34486),
            .I(alt_command_4));
    Odrv4 I__3774 (
            .O(N__34483),
            .I(alt_command_4));
    LocalMux I__3773 (
            .O(N__34480),
            .I(alt_command_4));
    CascadeMux I__3772 (
            .O(N__34473),
            .I(N__34470));
    InMux I__3771 (
            .O(N__34470),
            .I(N__34467));
    LocalMux I__3770 (
            .O(N__34467),
            .I(\pid_alt.alt_command_i_4 ));
    CascadeMux I__3769 (
            .O(N__34464),
            .I(N__34460));
    InMux I__3768 (
            .O(N__34463),
            .I(N__34456));
    InMux I__3767 (
            .O(N__34460),
            .I(N__34453));
    InMux I__3766 (
            .O(N__34459),
            .I(N__34450));
    LocalMux I__3765 (
            .O(N__34456),
            .I(alt_command_5));
    LocalMux I__3764 (
            .O(N__34453),
            .I(alt_command_5));
    LocalMux I__3763 (
            .O(N__34450),
            .I(alt_command_5));
    CascadeMux I__3762 (
            .O(N__34443),
            .I(N__34440));
    InMux I__3761 (
            .O(N__34440),
            .I(N__34437));
    LocalMux I__3760 (
            .O(N__34437),
            .I(\pid_alt.alt_command_i_5 ));
    InMux I__3759 (
            .O(N__34434),
            .I(N__34431));
    LocalMux I__3758 (
            .O(N__34431),
            .I(N__34426));
    InMux I__3757 (
            .O(N__34430),
            .I(N__34421));
    InMux I__3756 (
            .O(N__34429),
            .I(N__34421));
    Odrv4 I__3755 (
            .O(N__34426),
            .I(drone_altitude_10));
    LocalMux I__3754 (
            .O(N__34421),
            .I(drone_altitude_10));
    CascadeMux I__3753 (
            .O(N__34416),
            .I(N__34412));
    InMux I__3752 (
            .O(N__34415),
            .I(N__34408));
    InMux I__3751 (
            .O(N__34412),
            .I(N__34405));
    InMux I__3750 (
            .O(N__34411),
            .I(N__34402));
    LocalMux I__3749 (
            .O(N__34408),
            .I(alt_command_6));
    LocalMux I__3748 (
            .O(N__34405),
            .I(alt_command_6));
    LocalMux I__3747 (
            .O(N__34402),
            .I(alt_command_6));
    CascadeMux I__3746 (
            .O(N__34395),
            .I(N__34392));
    InMux I__3745 (
            .O(N__34392),
            .I(N__34389));
    LocalMux I__3744 (
            .O(N__34389),
            .I(\pid_alt.alt_command_i_6 ));
    InMux I__3743 (
            .O(N__34386),
            .I(N__34381));
    InMux I__3742 (
            .O(N__34385),
            .I(N__34376));
    InMux I__3741 (
            .O(N__34384),
            .I(N__34376));
    LocalMux I__3740 (
            .O(N__34381),
            .I(drone_altitude_11));
    LocalMux I__3739 (
            .O(N__34376),
            .I(drone_altitude_11));
    CascadeMux I__3738 (
            .O(N__34371),
            .I(N__34367));
    CascadeMux I__3737 (
            .O(N__34370),
            .I(N__34364));
    InMux I__3736 (
            .O(N__34367),
            .I(N__34360));
    InMux I__3735 (
            .O(N__34364),
            .I(N__34357));
    InMux I__3734 (
            .O(N__34363),
            .I(N__34354));
    LocalMux I__3733 (
            .O(N__34360),
            .I(alt_command_7));
    LocalMux I__3732 (
            .O(N__34357),
            .I(alt_command_7));
    LocalMux I__3731 (
            .O(N__34354),
            .I(alt_command_7));
    CascadeMux I__3730 (
            .O(N__34347),
            .I(N__34344));
    InMux I__3729 (
            .O(N__34344),
            .I(N__34341));
    LocalMux I__3728 (
            .O(N__34341),
            .I(\pid_alt.alt_command_i_7 ));
    InMux I__3727 (
            .O(N__34338),
            .I(N__34333));
    InMux I__3726 (
            .O(N__34337),
            .I(N__34328));
    InMux I__3725 (
            .O(N__34336),
            .I(N__34328));
    LocalMux I__3724 (
            .O(N__34333),
            .I(drone_altitude_12));
    LocalMux I__3723 (
            .O(N__34328),
            .I(drone_altitude_12));
    InMux I__3722 (
            .O(N__34323),
            .I(N__34320));
    LocalMux I__3721 (
            .O(N__34320),
            .I(N__34317));
    Span4Mux_v I__3720 (
            .O(N__34317),
            .I(N__34312));
    InMux I__3719 (
            .O(N__34316),
            .I(N__34307));
    InMux I__3718 (
            .O(N__34315),
            .I(N__34307));
    Odrv4 I__3717 (
            .O(N__34312),
            .I(drone_altitude_13));
    LocalMux I__3716 (
            .O(N__34307),
            .I(drone_altitude_13));
    InMux I__3715 (
            .O(N__34302),
            .I(N__34299));
    LocalMux I__3714 (
            .O(N__34299),
            .I(N__34296));
    Span4Mux_h I__3713 (
            .O(N__34296),
            .I(N__34291));
    InMux I__3712 (
            .O(N__34295),
            .I(N__34286));
    InMux I__3711 (
            .O(N__34294),
            .I(N__34286));
    Odrv4 I__3710 (
            .O(N__34291),
            .I(drone_altitude_14));
    LocalMux I__3709 (
            .O(N__34286),
            .I(drone_altitude_14));
    InMux I__3708 (
            .O(N__34281),
            .I(N__34276));
    InMux I__3707 (
            .O(N__34280),
            .I(N__34271));
    InMux I__3706 (
            .O(N__34279),
            .I(N__34271));
    LocalMux I__3705 (
            .O(N__34276),
            .I(N__34268));
    LocalMux I__3704 (
            .O(N__34271),
            .I(N__34265));
    Span4Mux_h I__3703 (
            .O(N__34268),
            .I(N__34262));
    Span12Mux_s5_h I__3702 (
            .O(N__34265),
            .I(N__34259));
    Span4Mux_v I__3701 (
            .O(N__34262),
            .I(N__34256));
    Span12Mux_v I__3700 (
            .O(N__34259),
            .I(N__34253));
    Span4Mux_v I__3699 (
            .O(N__34256),
            .I(N__34250));
    Odrv12 I__3698 (
            .O(N__34253),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    Odrv4 I__3697 (
            .O(N__34250),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__3696 (
            .O(N__34245),
            .I(N__34241));
    InMux I__3695 (
            .O(N__34244),
            .I(N__34238));
    LocalMux I__3694 (
            .O(N__34241),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    LocalMux I__3693 (
            .O(N__34238),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    InMux I__3692 (
            .O(N__34233),
            .I(N__34229));
    InMux I__3691 (
            .O(N__34232),
            .I(N__34226));
    LocalMux I__3690 (
            .O(N__34229),
            .I(N__34223));
    LocalMux I__3689 (
            .O(N__34226),
            .I(N__34220));
    Span4Mux_v I__3688 (
            .O(N__34223),
            .I(N__34216));
    Span4Mux_s2_h I__3687 (
            .O(N__34220),
            .I(N__34213));
    InMux I__3686 (
            .O(N__34219),
            .I(N__34210));
    Span4Mux_v I__3685 (
            .O(N__34216),
            .I(N__34207));
    Span4Mux_v I__3684 (
            .O(N__34213),
            .I(N__34204));
    LocalMux I__3683 (
            .O(N__34210),
            .I(N__34201));
    Span4Mux_v I__3682 (
            .O(N__34207),
            .I(N__34195));
    Span4Mux_v I__3681 (
            .O(N__34204),
            .I(N__34192));
    Span4Mux_s2_h I__3680 (
            .O(N__34201),
            .I(N__34189));
    InMux I__3679 (
            .O(N__34200),
            .I(N__34186));
    InMux I__3678 (
            .O(N__34199),
            .I(N__34181));
    InMux I__3677 (
            .O(N__34198),
            .I(N__34181));
    Odrv4 I__3676 (
            .O(N__34195),
            .I(drone_altitude_0));
    Odrv4 I__3675 (
            .O(N__34192),
            .I(drone_altitude_0));
    Odrv4 I__3674 (
            .O(N__34189),
            .I(drone_altitude_0));
    LocalMux I__3673 (
            .O(N__34186),
            .I(drone_altitude_0));
    LocalMux I__3672 (
            .O(N__34181),
            .I(drone_altitude_0));
    InMux I__3671 (
            .O(N__34170),
            .I(N__34165));
    InMux I__3670 (
            .O(N__34169),
            .I(N__34162));
    InMux I__3669 (
            .O(N__34168),
            .I(N__34159));
    LocalMux I__3668 (
            .O(N__34165),
            .I(drone_altitude_2));
    LocalMux I__3667 (
            .O(N__34162),
            .I(drone_altitude_2));
    LocalMux I__3666 (
            .O(N__34159),
            .I(drone_altitude_2));
    CascadeMux I__3665 (
            .O(N__34152),
            .I(N__34149));
    InMux I__3664 (
            .O(N__34149),
            .I(N__34144));
    InMux I__3663 (
            .O(N__34148),
            .I(N__34139));
    InMux I__3662 (
            .O(N__34147),
            .I(N__34139));
    LocalMux I__3661 (
            .O(N__34144),
            .I(drone_altitude_3));
    LocalMux I__3660 (
            .O(N__34139),
            .I(drone_altitude_3));
    InMux I__3659 (
            .O(N__34134),
            .I(N__34129));
    InMux I__3658 (
            .O(N__34133),
            .I(N__34124));
    InMux I__3657 (
            .O(N__34132),
            .I(N__34124));
    LocalMux I__3656 (
            .O(N__34129),
            .I(drone_altitude_4));
    LocalMux I__3655 (
            .O(N__34124),
            .I(drone_altitude_4));
    CascadeMux I__3654 (
            .O(N__34119),
            .I(N__34115));
    InMux I__3653 (
            .O(N__34118),
            .I(N__34111));
    InMux I__3652 (
            .O(N__34115),
            .I(N__34108));
    InMux I__3651 (
            .O(N__34114),
            .I(N__34105));
    LocalMux I__3650 (
            .O(N__34111),
            .I(alt_command_0));
    LocalMux I__3649 (
            .O(N__34108),
            .I(alt_command_0));
    LocalMux I__3648 (
            .O(N__34105),
            .I(alt_command_0));
    CascadeMux I__3647 (
            .O(N__34098),
            .I(N__34095));
    InMux I__3646 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__3645 (
            .O(N__34092),
            .I(\pid_alt.alt_command_i_0 ));
    CascadeMux I__3644 (
            .O(N__34089),
            .I(N__34084));
    InMux I__3643 (
            .O(N__34088),
            .I(N__34081));
    InMux I__3642 (
            .O(N__34087),
            .I(N__34078));
    InMux I__3641 (
            .O(N__34084),
            .I(N__34075));
    LocalMux I__3640 (
            .O(N__34081),
            .I(N__34072));
    LocalMux I__3639 (
            .O(N__34078),
            .I(alt_command_1));
    LocalMux I__3638 (
            .O(N__34075),
            .I(alt_command_1));
    Odrv4 I__3637 (
            .O(N__34072),
            .I(alt_command_1));
    CascadeMux I__3636 (
            .O(N__34065),
            .I(N__34062));
    InMux I__3635 (
            .O(N__34062),
            .I(N__34059));
    LocalMux I__3634 (
            .O(N__34059),
            .I(N__34056));
    Span4Mux_v I__3633 (
            .O(N__34056),
            .I(N__34051));
    InMux I__3632 (
            .O(N__34055),
            .I(N__34046));
    InMux I__3631 (
            .O(N__34054),
            .I(N__34046));
    Odrv4 I__3630 (
            .O(N__34051),
            .I(drone_altitude_5));
    LocalMux I__3629 (
            .O(N__34046),
            .I(drone_altitude_5));
    InMux I__3628 (
            .O(N__34041),
            .I(N__34038));
    LocalMux I__3627 (
            .O(N__34038),
            .I(\pid_alt.alt_command_i_1 ));
    InMux I__3626 (
            .O(N__34035),
            .I(N__34032));
    LocalMux I__3625 (
            .O(N__34032),
            .I(N__34028));
    InMux I__3624 (
            .O(N__34031),
            .I(N__34024));
    Span4Mux_h I__3623 (
            .O(N__34028),
            .I(N__34021));
    InMux I__3622 (
            .O(N__34027),
            .I(N__34018));
    LocalMux I__3621 (
            .O(N__34024),
            .I(drone_altitude_6));
    Odrv4 I__3620 (
            .O(N__34021),
            .I(drone_altitude_6));
    LocalMux I__3619 (
            .O(N__34018),
            .I(drone_altitude_6));
    CascadeMux I__3618 (
            .O(N__34011),
            .I(N__34008));
    InMux I__3617 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__3616 (
            .O(N__34005),
            .I(N__34001));
    InMux I__3615 (
            .O(N__34004),
            .I(N__33997));
    Span4Mux_s2_h I__3614 (
            .O(N__34001),
            .I(N__33994));
    InMux I__3613 (
            .O(N__34000),
            .I(N__33991));
    LocalMux I__3612 (
            .O(N__33997),
            .I(alt_command_2));
    Odrv4 I__3611 (
            .O(N__33994),
            .I(alt_command_2));
    LocalMux I__3610 (
            .O(N__33991),
            .I(alt_command_2));
    CascadeMux I__3609 (
            .O(N__33984),
            .I(N__33981));
    InMux I__3608 (
            .O(N__33981),
            .I(N__33978));
    LocalMux I__3607 (
            .O(N__33978),
            .I(\pid_alt.alt_command_i_2 ));
    InMux I__3606 (
            .O(N__33975),
            .I(N__33972));
    LocalMux I__3605 (
            .O(N__33972),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    CascadeMux I__3604 (
            .O(N__33969),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    InMux I__3603 (
            .O(N__33966),
            .I(N__33963));
    LocalMux I__3602 (
            .O(N__33963),
            .I(N__33960));
    Span4Mux_v I__3601 (
            .O(N__33960),
            .I(N__33955));
    InMux I__3600 (
            .O(N__33959),
            .I(N__33952));
    InMux I__3599 (
            .O(N__33958),
            .I(N__33949));
    Odrv4 I__3598 (
            .O(N__33955),
            .I(\pid_alt.un2_pid_prereg_cry_15_c_RNIP0DA ));
    LocalMux I__3597 (
            .O(N__33952),
            .I(\pid_alt.un2_pid_prereg_cry_15_c_RNIP0DA ));
    LocalMux I__3596 (
            .O(N__33949),
            .I(\pid_alt.un2_pid_prereg_cry_15_c_RNIP0DA ));
    InMux I__3595 (
            .O(N__33942),
            .I(N__33939));
    LocalMux I__3594 (
            .O(N__33939),
            .I(N__33936));
    Span4Mux_h I__3593 (
            .O(N__33936),
            .I(N__33933));
    Odrv4 I__3592 (
            .O(N__33933),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    InMux I__3591 (
            .O(N__33930),
            .I(N__33926));
    InMux I__3590 (
            .O(N__33929),
            .I(N__33923));
    LocalMux I__3589 (
            .O(N__33926),
            .I(N__33920));
    LocalMux I__3588 (
            .O(N__33923),
            .I(N__33917));
    Span4Mux_v I__3587 (
            .O(N__33920),
            .I(N__33911));
    Span4Mux_h I__3586 (
            .O(N__33917),
            .I(N__33911));
    InMux I__3585 (
            .O(N__33916),
            .I(N__33908));
    Odrv4 I__3584 (
            .O(N__33911),
            .I(\pid_alt.un2_pid_prereg_cry_6_c_RNINIBS ));
    LocalMux I__3583 (
            .O(N__33908),
            .I(\pid_alt.un2_pid_prereg_cry_6_c_RNINIBS ));
    InMux I__3582 (
            .O(N__33903),
            .I(N__33899));
    InMux I__3581 (
            .O(N__33902),
            .I(N__33896));
    LocalMux I__3580 (
            .O(N__33899),
            .I(N__33893));
    LocalMux I__3579 (
            .O(N__33896),
            .I(N__33888));
    Span4Mux_v I__3578 (
            .O(N__33893),
            .I(N__33888));
    Span4Mux_v I__3577 (
            .O(N__33888),
            .I(N__33885));
    Span4Mux_v I__3576 (
            .O(N__33885),
            .I(N__33882));
    Odrv4 I__3575 (
            .O(N__33882),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__3574 (
            .O(N__33879),
            .I(N__33876));
    LocalMux I__3573 (
            .O(N__33876),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    InMux I__3572 (
            .O(N__33873),
            .I(N__33867));
    InMux I__3571 (
            .O(N__33872),
            .I(N__33867));
    LocalMux I__3570 (
            .O(N__33867),
            .I(N__33864));
    Span4Mux_h I__3569 (
            .O(N__33864),
            .I(N__33861));
    Odrv4 I__3568 (
            .O(N__33861),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    CascadeMux I__3567 (
            .O(N__33858),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    InMux I__3566 (
            .O(N__33855),
            .I(N__33852));
    LocalMux I__3565 (
            .O(N__33852),
            .I(N__33847));
    InMux I__3564 (
            .O(N__33851),
            .I(N__33842));
    InMux I__3563 (
            .O(N__33850),
            .I(N__33842));
    Span4Mux_v I__3562 (
            .O(N__33847),
            .I(N__33839));
    LocalMux I__3561 (
            .O(N__33842),
            .I(N__33836));
    Odrv4 I__3560 (
            .O(N__33839),
            .I(\pid_alt.un2_pid_prereg_cry_18_c_RNIV9GA ));
    Odrv4 I__3559 (
            .O(N__33836),
            .I(\pid_alt.un2_pid_prereg_cry_18_c_RNIV9GA ));
    CascadeMux I__3558 (
            .O(N__33831),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ));
    InMux I__3557 (
            .O(N__33828),
            .I(N__33822));
    InMux I__3556 (
            .O(N__33827),
            .I(N__33822));
    LocalMux I__3555 (
            .O(N__33822),
            .I(N__33818));
    InMux I__3554 (
            .O(N__33821),
            .I(N__33815));
    Span4Mux_v I__3553 (
            .O(N__33818),
            .I(N__33810));
    LocalMux I__3552 (
            .O(N__33815),
            .I(N__33810));
    Span4Mux_v I__3551 (
            .O(N__33810),
            .I(N__33807));
    Span4Mux_v I__3550 (
            .O(N__33807),
            .I(N__33804));
    Odrv4 I__3549 (
            .O(N__33804),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    InMux I__3548 (
            .O(N__33801),
            .I(N__33797));
    InMux I__3547 (
            .O(N__33800),
            .I(N__33794));
    LocalMux I__3546 (
            .O(N__33797),
            .I(N__33791));
    LocalMux I__3545 (
            .O(N__33794),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    Odrv4 I__3544 (
            .O(N__33791),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    InMux I__3543 (
            .O(N__33786),
            .I(N__33783));
    LocalMux I__3542 (
            .O(N__33783),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    InMux I__3541 (
            .O(N__33780),
            .I(N__33773));
    InMux I__3540 (
            .O(N__33779),
            .I(N__33773));
    InMux I__3539 (
            .O(N__33778),
            .I(N__33770));
    LocalMux I__3538 (
            .O(N__33773),
            .I(N__33767));
    LocalMux I__3537 (
            .O(N__33770),
            .I(N__33764));
    Span4Mux_v I__3536 (
            .O(N__33767),
            .I(N__33761));
    Odrv4 I__3535 (
            .O(N__33764),
            .I(\pid_alt.un2_pid_prereg_cry_8_c_RNITQDS ));
    Odrv4 I__3534 (
            .O(N__33761),
            .I(\pid_alt.un2_pid_prereg_cry_8_c_RNITQDS ));
    InMux I__3533 (
            .O(N__33756),
            .I(N__33750));
    InMux I__3532 (
            .O(N__33755),
            .I(N__33750));
    LocalMux I__3531 (
            .O(N__33750),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__3530 (
            .O(N__33747),
            .I(N__33741));
    InMux I__3529 (
            .O(N__33746),
            .I(N__33741));
    LocalMux I__3528 (
            .O(N__33741),
            .I(N__33738));
    Span4Mux_v I__3527 (
            .O(N__33738),
            .I(N__33735));
    Span4Mux_v I__3526 (
            .O(N__33735),
            .I(N__33732));
    Span4Mux_v I__3525 (
            .O(N__33732),
            .I(N__33729));
    Odrv4 I__3524 (
            .O(N__33729),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    InMux I__3523 (
            .O(N__33726),
            .I(N__33719));
    InMux I__3522 (
            .O(N__33725),
            .I(N__33719));
    InMux I__3521 (
            .O(N__33724),
            .I(N__33716));
    LocalMux I__3520 (
            .O(N__33719),
            .I(N__33711));
    LocalMux I__3519 (
            .O(N__33716),
            .I(N__33711));
    Span12Mux_v I__3518 (
            .O(N__33711),
            .I(N__33708));
    Odrv12 I__3517 (
            .O(N__33708),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__3516 (
            .O(N__33705),
            .I(N__33702));
    LocalMux I__3515 (
            .O(N__33702),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    CascadeMux I__3514 (
            .O(N__33699),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ));
    InMux I__3513 (
            .O(N__33696),
            .I(N__33693));
    LocalMux I__3512 (
            .O(N__33693),
            .I(N__33690));
    Span4Mux_v I__3511 (
            .O(N__33690),
            .I(N__33685));
    InMux I__3510 (
            .O(N__33689),
            .I(N__33680));
    InMux I__3509 (
            .O(N__33688),
            .I(N__33680));
    Odrv4 I__3508 (
            .O(N__33685),
            .I(\pid_alt.un2_pid_prereg_cry_16_c_RNIR3EA ));
    LocalMux I__3507 (
            .O(N__33680),
            .I(\pid_alt.un2_pid_prereg_cry_16_c_RNIR3EA ));
    CascadeMux I__3506 (
            .O(N__33675),
            .I(N__33672));
    InMux I__3505 (
            .O(N__33672),
            .I(N__33668));
    InMux I__3504 (
            .O(N__33671),
            .I(N__33665));
    LocalMux I__3503 (
            .O(N__33668),
            .I(N__33660));
    LocalMux I__3502 (
            .O(N__33665),
            .I(N__33660));
    Span12Mux_v I__3501 (
            .O(N__33660),
            .I(N__33657));
    Odrv12 I__3500 (
            .O(N__33657),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    InMux I__3499 (
            .O(N__33654),
            .I(N__33648));
    InMux I__3498 (
            .O(N__33653),
            .I(N__33648));
    LocalMux I__3497 (
            .O(N__33648),
            .I(N__33645));
    Odrv4 I__3496 (
            .O(N__33645),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    InMux I__3495 (
            .O(N__33642),
            .I(N__33636));
    InMux I__3494 (
            .O(N__33641),
            .I(N__33636));
    LocalMux I__3493 (
            .O(N__33636),
            .I(N__33632));
    InMux I__3492 (
            .O(N__33635),
            .I(N__33629));
    Span4Mux_v I__3491 (
            .O(N__33632),
            .I(N__33624));
    LocalMux I__3490 (
            .O(N__33629),
            .I(N__33624));
    Span4Mux_v I__3489 (
            .O(N__33624),
            .I(N__33621));
    Span4Mux_v I__3488 (
            .O(N__33621),
            .I(N__33618));
    Odrv4 I__3487 (
            .O(N__33618),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    InMux I__3486 (
            .O(N__33615),
            .I(N__33611));
    InMux I__3485 (
            .O(N__33614),
            .I(N__33608));
    LocalMux I__3484 (
            .O(N__33611),
            .I(N__33605));
    LocalMux I__3483 (
            .O(N__33608),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    Odrv4 I__3482 (
            .O(N__33605),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__3481 (
            .O(N__33600),
            .I(N__33597));
    LocalMux I__3480 (
            .O(N__33597),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    InMux I__3479 (
            .O(N__33594),
            .I(N__33585));
    InMux I__3478 (
            .O(N__33593),
            .I(N__33585));
    InMux I__3477 (
            .O(N__33592),
            .I(N__33585));
    LocalMux I__3476 (
            .O(N__33585),
            .I(N__33582));
    Span4Mux_v I__3475 (
            .O(N__33582),
            .I(N__33579));
    Span4Mux_v I__3474 (
            .O(N__33579),
            .I(N__33576));
    Odrv4 I__3473 (
            .O(N__33576),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    InMux I__3472 (
            .O(N__33573),
            .I(N__33567));
    InMux I__3471 (
            .O(N__33572),
            .I(N__33567));
    LocalMux I__3470 (
            .O(N__33567),
            .I(N__33564));
    Span4Mux_v I__3469 (
            .O(N__33564),
            .I(N__33561));
    Span4Mux_v I__3468 (
            .O(N__33561),
            .I(N__33558));
    Span4Mux_v I__3467 (
            .O(N__33558),
            .I(N__33555));
    Odrv4 I__3466 (
            .O(N__33555),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    CascadeMux I__3465 (
            .O(N__33552),
            .I(N__33549));
    InMux I__3464 (
            .O(N__33549),
            .I(N__33543));
    InMux I__3463 (
            .O(N__33548),
            .I(N__33543));
    LocalMux I__3462 (
            .O(N__33543),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__3461 (
            .O(N__33540),
            .I(N__33537));
    LocalMux I__3460 (
            .O(N__33537),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    CascadeMux I__3459 (
            .O(N__33534),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ));
    InMux I__3458 (
            .O(N__33531),
            .I(N__33528));
    LocalMux I__3457 (
            .O(N__33528),
            .I(N__33525));
    Span4Mux_h I__3456 (
            .O(N__33525),
            .I(N__33520));
    InMux I__3455 (
            .O(N__33524),
            .I(N__33515));
    InMux I__3454 (
            .O(N__33523),
            .I(N__33515));
    Odrv4 I__3453 (
            .O(N__33520),
            .I(\pid_alt.un2_pid_prereg_cry_9_c_RNIEPOG ));
    LocalMux I__3452 (
            .O(N__33515),
            .I(\pid_alt.un2_pid_prereg_cry_9_c_RNIEPOG ));
    InMux I__3451 (
            .O(N__33510),
            .I(N__33507));
    LocalMux I__3450 (
            .O(N__33507),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    CascadeMux I__3449 (
            .O(N__33504),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17_cascade_ ));
    InMux I__3448 (
            .O(N__33501),
            .I(N__33498));
    LocalMux I__3447 (
            .O(N__33498),
            .I(N__33495));
    Span4Mux_v I__3446 (
            .O(N__33495),
            .I(N__33490));
    InMux I__3445 (
            .O(N__33494),
            .I(N__33485));
    InMux I__3444 (
            .O(N__33493),
            .I(N__33485));
    Odrv4 I__3443 (
            .O(N__33490),
            .I(\pid_alt.un2_pid_prereg_cry_17_c_RNIT6FA ));
    LocalMux I__3442 (
            .O(N__33485),
            .I(\pid_alt.un2_pid_prereg_cry_17_c_RNIT6FA ));
    InMux I__3441 (
            .O(N__33480),
            .I(N__33474));
    InMux I__3440 (
            .O(N__33479),
            .I(N__33474));
    LocalMux I__3439 (
            .O(N__33474),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    InMux I__3438 (
            .O(N__33471),
            .I(N__33465));
    InMux I__3437 (
            .O(N__33470),
            .I(N__33465));
    LocalMux I__3436 (
            .O(N__33465),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    InMux I__3435 (
            .O(N__33462),
            .I(N__33453));
    InMux I__3434 (
            .O(N__33461),
            .I(N__33453));
    InMux I__3433 (
            .O(N__33460),
            .I(N__33453));
    LocalMux I__3432 (
            .O(N__33453),
            .I(N__33450));
    Span12Mux_h I__3431 (
            .O(N__33450),
            .I(N__33447));
    Odrv12 I__3430 (
            .O(N__33447),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    CascadeMux I__3429 (
            .O(N__33444),
            .I(N__33441));
    InMux I__3428 (
            .O(N__33441),
            .I(N__33435));
    InMux I__3427 (
            .O(N__33440),
            .I(N__33435));
    LocalMux I__3426 (
            .O(N__33435),
            .I(N__33432));
    Span4Mux_h I__3425 (
            .O(N__33432),
            .I(N__33429));
    Span4Mux_v I__3424 (
            .O(N__33429),
            .I(N__33426));
    Span4Mux_v I__3423 (
            .O(N__33426),
            .I(N__33423));
    Odrv4 I__3422 (
            .O(N__33423),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__3421 (
            .O(N__33420),
            .I(N__33414));
    InMux I__3420 (
            .O(N__33419),
            .I(N__33414));
    LocalMux I__3419 (
            .O(N__33414),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    InMux I__3418 (
            .O(N__33411),
            .I(N__33408));
    LocalMux I__3417 (
            .O(N__33408),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    CascadeMux I__3416 (
            .O(N__33405),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__3415 (
            .O(N__33402),
            .I(N__33399));
    LocalMux I__3414 (
            .O(N__33399),
            .I(N__33396));
    Span4Mux_h I__3413 (
            .O(N__33396),
            .I(N__33391));
    InMux I__3412 (
            .O(N__33395),
            .I(N__33386));
    InMux I__3411 (
            .O(N__33394),
            .I(N__33386));
    Odrv4 I__3410 (
            .O(N__33391),
            .I(\pid_alt.un2_pid_prereg_cry_11_c_RNIRGEG ));
    LocalMux I__3409 (
            .O(N__33386),
            .I(\pid_alt.un2_pid_prereg_cry_11_c_RNIRGEG ));
    InMux I__3408 (
            .O(N__33381),
            .I(N__33378));
    LocalMux I__3407 (
            .O(N__33378),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    CascadeMux I__3406 (
            .O(N__33375),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ));
    InMux I__3405 (
            .O(N__33372),
            .I(N__33369));
    LocalMux I__3404 (
            .O(N__33369),
            .I(N__33366));
    Span4Mux_h I__3403 (
            .O(N__33366),
            .I(N__33361));
    InMux I__3402 (
            .O(N__33365),
            .I(N__33356));
    InMux I__3401 (
            .O(N__33364),
            .I(N__33356));
    Odrv4 I__3400 (
            .O(N__33361),
            .I(\pid_alt.un2_pid_prereg_cry_10_c_RNIOCDG ));
    LocalMux I__3399 (
            .O(N__33356),
            .I(\pid_alt.un2_pid_prereg_cry_10_c_RNIOCDG ));
    InMux I__3398 (
            .O(N__33351),
            .I(N__33345));
    InMux I__3397 (
            .O(N__33350),
            .I(N__33345));
    LocalMux I__3396 (
            .O(N__33345),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ));
    CascadeMux I__3395 (
            .O(N__33342),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ));
    InMux I__3394 (
            .O(N__33339),
            .I(N__33336));
    LocalMux I__3393 (
            .O(N__33336),
            .I(N__33331));
    InMux I__3392 (
            .O(N__33335),
            .I(N__33326));
    InMux I__3391 (
            .O(N__33334),
            .I(N__33326));
    Odrv4 I__3390 (
            .O(N__33331),
            .I(\pid_alt.un2_pid_prereg_cry_4_c_RNIHA9S ));
    LocalMux I__3389 (
            .O(N__33326),
            .I(\pid_alt.un2_pid_prereg_cry_4_c_RNIHA9S ));
    InMux I__3388 (
            .O(N__33321),
            .I(N__33315));
    InMux I__3387 (
            .O(N__33320),
            .I(N__33315));
    LocalMux I__3386 (
            .O(N__33315),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    InMux I__3385 (
            .O(N__33312),
            .I(N__33306));
    InMux I__3384 (
            .O(N__33311),
            .I(N__33306));
    LocalMux I__3383 (
            .O(N__33306),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__3382 (
            .O(N__33303),
            .I(N__33299));
    InMux I__3381 (
            .O(N__33302),
            .I(N__33296));
    LocalMux I__3380 (
            .O(N__33299),
            .I(N__33291));
    LocalMux I__3379 (
            .O(N__33296),
            .I(N__33291));
    Span12Mux_s4_h I__3378 (
            .O(N__33291),
            .I(N__33288));
    Span12Mux_v I__3377 (
            .O(N__33288),
            .I(N__33285));
    Odrv12 I__3376 (
            .O(N__33285),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    InMux I__3375 (
            .O(N__33282),
            .I(N__33273));
    InMux I__3374 (
            .O(N__33281),
            .I(N__33273));
    InMux I__3373 (
            .O(N__33280),
            .I(N__33273));
    LocalMux I__3372 (
            .O(N__33273),
            .I(N__33270));
    Span12Mux_h I__3371 (
            .O(N__33270),
            .I(N__33267));
    Odrv12 I__3370 (
            .O(N__33267),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    InMux I__3369 (
            .O(N__33264),
            .I(N__33261));
    LocalMux I__3368 (
            .O(N__33261),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    InMux I__3367 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__3366 (
            .O(N__33255),
            .I(N__33250));
    InMux I__3365 (
            .O(N__33254),
            .I(N__33245));
    InMux I__3364 (
            .O(N__33253),
            .I(N__33245));
    Odrv4 I__3363 (
            .O(N__33250),
            .I(\pid_alt.un2_pid_prereg_cry_3_c_RNIN46R ));
    LocalMux I__3362 (
            .O(N__33245),
            .I(\pid_alt.un2_pid_prereg_cry_3_c_RNIN46R ));
    CascadeMux I__3361 (
            .O(N__33240),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ));
    InMux I__3360 (
            .O(N__33237),
            .I(N__33234));
    LocalMux I__3359 (
            .O(N__33234),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    CascadeMux I__3358 (
            .O(N__33231),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ));
    InMux I__3357 (
            .O(N__33228),
            .I(N__33225));
    LocalMux I__3356 (
            .O(N__33225),
            .I(N__33222));
    Span4Mux_h I__3355 (
            .O(N__33222),
            .I(N__33217));
    InMux I__3354 (
            .O(N__33221),
            .I(N__33212));
    InMux I__3353 (
            .O(N__33220),
            .I(N__33212));
    Odrv4 I__3352 (
            .O(N__33217),
            .I(\pid_alt.un2_pid_prereg_cry_12_c_RNI7SBD ));
    LocalMux I__3351 (
            .O(N__33212),
            .I(\pid_alt.un2_pid_prereg_cry_12_c_RNI7SBD ));
    InMux I__3350 (
            .O(N__33207),
            .I(N__33202));
    InMux I__3349 (
            .O(N__33206),
            .I(N__33199));
    InMux I__3348 (
            .O(N__33205),
            .I(N__33196));
    LocalMux I__3347 (
            .O(N__33202),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3346 (
            .O(N__33199),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3345 (
            .O(N__33196),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__3344 (
            .O(N__33189),
            .I(N__33184));
    InMux I__3343 (
            .O(N__33188),
            .I(N__33179));
    InMux I__3342 (
            .O(N__33187),
            .I(N__33179));
    LocalMux I__3341 (
            .O(N__33184),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__3340 (
            .O(N__33179),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    CascadeMux I__3339 (
            .O(N__33174),
            .I(N__33170));
    InMux I__3338 (
            .O(N__33173),
            .I(N__33166));
    InMux I__3337 (
            .O(N__33170),
            .I(N__33163));
    InMux I__3336 (
            .O(N__33169),
            .I(N__33160));
    LocalMux I__3335 (
            .O(N__33166),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__3334 (
            .O(N__33163),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__3333 (
            .O(N__33160),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    InMux I__3332 (
            .O(N__33153),
            .I(N__33148));
    InMux I__3331 (
            .O(N__33152),
            .I(N__33143));
    InMux I__3330 (
            .O(N__33151),
            .I(N__33143));
    LocalMux I__3329 (
            .O(N__33148),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__3328 (
            .O(N__33143),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    CascadeMux I__3327 (
            .O(N__33138),
            .I(N__33135));
    InMux I__3326 (
            .O(N__33135),
            .I(N__33132));
    LocalMux I__3325 (
            .O(N__33132),
            .I(N__33129));
    Span4Mux_h I__3324 (
            .O(N__33129),
            .I(N__33125));
    InMux I__3323 (
            .O(N__33128),
            .I(N__33122));
    Odrv4 I__3322 (
            .O(N__33125),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__3321 (
            .O(N__33122),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    InMux I__3320 (
            .O(N__33117),
            .I(N__33114));
    LocalMux I__3319 (
            .O(N__33114),
            .I(N__33110));
    InMux I__3318 (
            .O(N__33113),
            .I(N__33107));
    Odrv4 I__3317 (
            .O(N__33110),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    LocalMux I__3316 (
            .O(N__33107),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    CascadeMux I__3315 (
            .O(N__33102),
            .I(\pid_alt.m21_e_8_cascade_ ));
    InMux I__3314 (
            .O(N__33099),
            .I(N__33096));
    LocalMux I__3313 (
            .O(N__33096),
            .I(\pid_alt.m21_e_2 ));
    InMux I__3312 (
            .O(N__33093),
            .I(N__33090));
    LocalMux I__3311 (
            .O(N__33090),
            .I(N__33085));
    InMux I__3310 (
            .O(N__33089),
            .I(N__33080));
    InMux I__3309 (
            .O(N__33088),
            .I(N__33080));
    Odrv4 I__3308 (
            .O(N__33085),
            .I(\pid_alt.un2_pid_prereg_cry_5_c_RNIKEAS ));
    LocalMux I__3307 (
            .O(N__33080),
            .I(\pid_alt.un2_pid_prereg_cry_5_c_RNIKEAS ));
    CascadeMux I__3306 (
            .O(N__33075),
            .I(N__33071));
    CascadeMux I__3305 (
            .O(N__33074),
            .I(N__33067));
    InMux I__3304 (
            .O(N__33071),
            .I(N__33062));
    InMux I__3303 (
            .O(N__33070),
            .I(N__33062));
    InMux I__3302 (
            .O(N__33067),
            .I(N__33059));
    LocalMux I__3301 (
            .O(N__33062),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__3300 (
            .O(N__33059),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__3299 (
            .O(N__33054),
            .I(N__33049));
    InMux I__3298 (
            .O(N__33053),
            .I(N__33044));
    InMux I__3297 (
            .O(N__33052),
            .I(N__33044));
    LocalMux I__3296 (
            .O(N__33049),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__3295 (
            .O(N__33044),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    InMux I__3294 (
            .O(N__33039),
            .I(N__33035));
    InMux I__3293 (
            .O(N__33038),
            .I(N__33031));
    LocalMux I__3292 (
            .O(N__33035),
            .I(N__33028));
    InMux I__3291 (
            .O(N__33034),
            .I(N__33025));
    LocalMux I__3290 (
            .O(N__33031),
            .I(N__33022));
    Span4Mux_v I__3289 (
            .O(N__33028),
            .I(N__33019));
    LocalMux I__3288 (
            .O(N__33025),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    Odrv12 I__3287 (
            .O(N__33022),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    Odrv4 I__3286 (
            .O(N__33019),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    InMux I__3285 (
            .O(N__33012),
            .I(N__33008));
    InMux I__3284 (
            .O(N__33011),
            .I(N__33005));
    LocalMux I__3283 (
            .O(N__33008),
            .I(N__33002));
    LocalMux I__3282 (
            .O(N__33005),
            .I(N__32997));
    Span4Mux_h I__3281 (
            .O(N__33002),
            .I(N__32997));
    Span4Mux_v I__3280 (
            .O(N__32997),
            .I(N__32994));
    Span4Mux_v I__3279 (
            .O(N__32994),
            .I(N__32991));
    Odrv4 I__3278 (
            .O(N__32991),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__3277 (
            .O(N__32988),
            .I(N__32984));
    InMux I__3276 (
            .O(N__32987),
            .I(N__32981));
    LocalMux I__3275 (
            .O(N__32984),
            .I(N__32978));
    LocalMux I__3274 (
            .O(N__32981),
            .I(N__32975));
    Span4Mux_v I__3273 (
            .O(N__32978),
            .I(N__32972));
    Span4Mux_v I__3272 (
            .O(N__32975),
            .I(N__32969));
    Odrv4 I__3271 (
            .O(N__32972),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    Odrv4 I__3270 (
            .O(N__32969),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    InMux I__3269 (
            .O(N__32964),
            .I(N__32961));
    LocalMux I__3268 (
            .O(N__32961),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    InMux I__3267 (
            .O(N__32958),
            .I(N__32955));
    LocalMux I__3266 (
            .O(N__32955),
            .I(N__32951));
    CascadeMux I__3265 (
            .O(N__32954),
            .I(N__32948));
    Span4Mux_h I__3264 (
            .O(N__32951),
            .I(N__32945));
    InMux I__3263 (
            .O(N__32948),
            .I(N__32942));
    Odrv4 I__3262 (
            .O(N__32945),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    LocalMux I__3261 (
            .O(N__32942),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__3260 (
            .O(N__32937),
            .I(N__32934));
    LocalMux I__3259 (
            .O(N__32934),
            .I(N__32930));
    InMux I__3258 (
            .O(N__32933),
            .I(N__32927));
    Odrv4 I__3257 (
            .O(N__32930),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    LocalMux I__3256 (
            .O(N__32927),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__3255 (
            .O(N__32922),
            .I(N__32919));
    LocalMux I__3254 (
            .O(N__32919),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    CascadeMux I__3253 (
            .O(N__32916),
            .I(N__32913));
    InMux I__3252 (
            .O(N__32913),
            .I(N__32910));
    LocalMux I__3251 (
            .O(N__32910),
            .I(\pid_alt.m35_e_3 ));
    InMux I__3250 (
            .O(N__32907),
            .I(N__32904));
    LocalMux I__3249 (
            .O(N__32904),
            .I(N__32901));
    Odrv4 I__3248 (
            .O(N__32901),
            .I(alt_kp_3));
    InMux I__3247 (
            .O(N__32898),
            .I(N__32895));
    LocalMux I__3246 (
            .O(N__32895),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    CascadeMux I__3245 (
            .O(N__32892),
            .I(\pid_alt.m7_e_4_cascade_ ));
    CascadeMux I__3244 (
            .O(N__32889),
            .I(\pid_alt.N_222_cascade_ ));
    InMux I__3243 (
            .O(N__32886),
            .I(N__32883));
    LocalMux I__3242 (
            .O(N__32883),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__3241 (
            .O(N__32880),
            .I(N__32877));
    LocalMux I__3240 (
            .O(N__32877),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    InMux I__3239 (
            .O(N__32874),
            .I(N__32871));
    LocalMux I__3238 (
            .O(N__32871),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__3237 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__3236 (
            .O(N__32865),
            .I(N__32862));
    Span4Mux_v I__3235 (
            .O(N__32862),
            .I(N__32857));
    InMux I__3234 (
            .O(N__32861),
            .I(N__32852));
    InMux I__3233 (
            .O(N__32860),
            .I(N__32852));
    Odrv4 I__3232 (
            .O(N__32857),
            .I(\pid_alt.un2_pid_prereg_cry_19_c_RNIO4IA ));
    LocalMux I__3231 (
            .O(N__32852),
            .I(\pid_alt.un2_pid_prereg_cry_19_c_RNIO4IA ));
    CascadeMux I__3230 (
            .O(N__32847),
            .I(N__32844));
    InMux I__3229 (
            .O(N__32844),
            .I(N__32841));
    LocalMux I__3228 (
            .O(N__32841),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__3227 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__3226 (
            .O(N__32835),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__3225 (
            .O(N__32832),
            .I(N__32829));
    LocalMux I__3224 (
            .O(N__32829),
            .I(N__32826));
    Span4Mux_s2_h I__3223 (
            .O(N__32826),
            .I(N__32823));
    Odrv4 I__3222 (
            .O(N__32823),
            .I(alt_kp_6));
    InMux I__3221 (
            .O(N__32820),
            .I(N__32817));
    LocalMux I__3220 (
            .O(N__32817),
            .I(N__32814));
    Span4Mux_s2_h I__3219 (
            .O(N__32814),
            .I(N__32811));
    Odrv4 I__3218 (
            .O(N__32811),
            .I(alt_kp_2));
    InMux I__3217 (
            .O(N__32808),
            .I(N__32805));
    LocalMux I__3216 (
            .O(N__32805),
            .I(N__32802));
    Span4Mux_v I__3215 (
            .O(N__32802),
            .I(N__32799));
    Odrv4 I__3214 (
            .O(N__32799),
            .I(alt_kp_7));
    InMux I__3213 (
            .O(N__32796),
            .I(N__32793));
    LocalMux I__3212 (
            .O(N__32793),
            .I(N__32790));
    Span4Mux_v I__3211 (
            .O(N__32790),
            .I(N__32787));
    Odrv4 I__3210 (
            .O(N__32787),
            .I(alt_kp_1));
    CascadeMux I__3209 (
            .O(N__32784),
            .I(N__32781));
    InMux I__3208 (
            .O(N__32781),
            .I(N__32778));
    LocalMux I__3207 (
            .O(N__32778),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__3206 (
            .O(N__32775),
            .I(N__32772));
    LocalMux I__3205 (
            .O(N__32772),
            .I(drone_altitude_i_4));
    InMux I__3204 (
            .O(N__32769),
            .I(N__32766));
    LocalMux I__3203 (
            .O(N__32766),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__3202 (
            .O(N__32763),
            .I(N__32759));
    InMux I__3201 (
            .O(N__32762),
            .I(N__32756));
    LocalMux I__3200 (
            .O(N__32759),
            .I(\pid_alt.drone_altitude_i_0 ));
    LocalMux I__3199 (
            .O(N__32756),
            .I(\pid_alt.drone_altitude_i_0 ));
    CascadeMux I__3198 (
            .O(N__32751),
            .I(N__32748));
    InMux I__3197 (
            .O(N__32748),
            .I(N__32745));
    LocalMux I__3196 (
            .O(N__32745),
            .I(N__32742));
    Odrv4 I__3195 (
            .O(N__32742),
            .I(drone_altitude_i_8));
    InMux I__3194 (
            .O(N__32739),
            .I(N__32736));
    LocalMux I__3193 (
            .O(N__32736),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__3192 (
            .O(N__32733),
            .I(N__32730));
    LocalMux I__3191 (
            .O(N__32730),
            .I(N__32727));
    Odrv4 I__3190 (
            .O(N__32727),
            .I(drone_altitude_i_10));
    InMux I__3189 (
            .O(N__32724),
            .I(N__32721));
    LocalMux I__3188 (
            .O(N__32721),
            .I(drone_altitude_i_11));
    InMux I__3187 (
            .O(N__32718),
            .I(N__32712));
    InMux I__3186 (
            .O(N__32717),
            .I(N__32712));
    LocalMux I__3185 (
            .O(N__32712),
            .I(N__32709));
    Span4Mux_v I__3184 (
            .O(N__32709),
            .I(N__32706));
    Odrv4 I__3183 (
            .O(N__32706),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__3182 (
            .O(N__32703),
            .I(\pid_alt.un2_pid_prereg_cry_20 ));
    CascadeMux I__3181 (
            .O(N__32700),
            .I(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB_cascade_ ));
    CascadeMux I__3180 (
            .O(N__32697),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15_cascade_ ));
    InMux I__3179 (
            .O(N__32694),
            .I(N__32691));
    LocalMux I__3178 (
            .O(N__32691),
            .I(N__32684));
    InMux I__3177 (
            .O(N__32690),
            .I(N__32681));
    InMux I__3176 (
            .O(N__32689),
            .I(N__32674));
    InMux I__3175 (
            .O(N__32688),
            .I(N__32674));
    InMux I__3174 (
            .O(N__32687),
            .I(N__32674));
    Odrv12 I__3173 (
            .O(N__32684),
            .I(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB ));
    LocalMux I__3172 (
            .O(N__32681),
            .I(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB ));
    LocalMux I__3171 (
            .O(N__32674),
            .I(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB ));
    CascadeMux I__3170 (
            .O(N__32667),
            .I(N__32664));
    InMux I__3169 (
            .O(N__32664),
            .I(N__32656));
    InMux I__3168 (
            .O(N__32663),
            .I(N__32656));
    CascadeMux I__3167 (
            .O(N__32662),
            .I(N__32652));
    CascadeMux I__3166 (
            .O(N__32661),
            .I(N__32649));
    LocalMux I__3165 (
            .O(N__32656),
            .I(N__32645));
    InMux I__3164 (
            .O(N__32655),
            .I(N__32638));
    InMux I__3163 (
            .O(N__32652),
            .I(N__32638));
    InMux I__3162 (
            .O(N__32649),
            .I(N__32638));
    InMux I__3161 (
            .O(N__32648),
            .I(N__32635));
    Span4Mux_h I__3160 (
            .O(N__32645),
            .I(N__32630));
    LocalMux I__3159 (
            .O(N__32638),
            .I(N__32630));
    LocalMux I__3158 (
            .O(N__32635),
            .I(N__32627));
    Span4Mux_v I__3157 (
            .O(N__32630),
            .I(N__32624));
    Sp12to4 I__3156 (
            .O(N__32627),
            .I(N__32621));
    Odrv4 I__3155 (
            .O(N__32624),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    Odrv12 I__3154 (
            .O(N__32621),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    CascadeMux I__3153 (
            .O(N__32616),
            .I(N__32613));
    InMux I__3152 (
            .O(N__32613),
            .I(N__32604));
    InMux I__3151 (
            .O(N__32612),
            .I(N__32604));
    InMux I__3150 (
            .O(N__32611),
            .I(N__32604));
    LocalMux I__3149 (
            .O(N__32604),
            .I(N__32599));
    InMux I__3148 (
            .O(N__32603),
            .I(N__32594));
    InMux I__3147 (
            .O(N__32602),
            .I(N__32594));
    Span4Mux_v I__3146 (
            .O(N__32599),
            .I(N__32591));
    LocalMux I__3145 (
            .O(N__32594),
            .I(N__32584));
    Sp12to4 I__3144 (
            .O(N__32591),
            .I(N__32584));
    InMux I__3143 (
            .O(N__32590),
            .I(N__32579));
    InMux I__3142 (
            .O(N__32589),
            .I(N__32579));
    Span12Mux_h I__3141 (
            .O(N__32584),
            .I(N__32574));
    LocalMux I__3140 (
            .O(N__32579),
            .I(N__32574));
    Odrv12 I__3139 (
            .O(N__32574),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    InMux I__3138 (
            .O(N__32571),
            .I(N__32560));
    InMux I__3137 (
            .O(N__32570),
            .I(N__32560));
    InMux I__3136 (
            .O(N__32569),
            .I(N__32560));
    InMux I__3135 (
            .O(N__32568),
            .I(N__32554));
    InMux I__3134 (
            .O(N__32567),
            .I(N__32554));
    LocalMux I__3133 (
            .O(N__32560),
            .I(N__32551));
    InMux I__3132 (
            .O(N__32559),
            .I(N__32548));
    LocalMux I__3131 (
            .O(N__32554),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    Odrv4 I__3130 (
            .O(N__32551),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__3129 (
            .O(N__32548),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__3128 (
            .O(N__32541),
            .I(N__32538));
    LocalMux I__3127 (
            .O(N__32538),
            .I(N__32535));
    Span4Mux_v I__3126 (
            .O(N__32535),
            .I(N__32532));
    Odrv4 I__3125 (
            .O(N__32532),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    CascadeMux I__3124 (
            .O(N__32529),
            .I(N__32526));
    InMux I__3123 (
            .O(N__32526),
            .I(N__32522));
    InMux I__3122 (
            .O(N__32525),
            .I(N__32519));
    LocalMux I__3121 (
            .O(N__32522),
            .I(N__32516));
    LocalMux I__3120 (
            .O(N__32519),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    Odrv4 I__3119 (
            .O(N__32516),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__3118 (
            .O(N__32511),
            .I(\pid_alt.un2_pid_prereg_cry_11 ));
    CascadeMux I__3117 (
            .O(N__32508),
            .I(N__32505));
    InMux I__3116 (
            .O(N__32505),
            .I(N__32502));
    LocalMux I__3115 (
            .O(N__32502),
            .I(N__32499));
    Odrv4 I__3114 (
            .O(N__32499),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__3113 (
            .O(N__32496),
            .I(\pid_alt.un2_pid_prereg_cry_12 ));
    InMux I__3112 (
            .O(N__32493),
            .I(N__32490));
    LocalMux I__3111 (
            .O(N__32490),
            .I(N__32487));
    Span4Mux_v I__3110 (
            .O(N__32487),
            .I(N__32484));
    Odrv4 I__3109 (
            .O(N__32484),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__3108 (
            .O(N__32481),
            .I(\pid_alt.un2_pid_prereg_cry_13 ));
    InMux I__3107 (
            .O(N__32478),
            .I(N__32475));
    LocalMux I__3106 (
            .O(N__32475),
            .I(N__32472));
    Span4Mux_h I__3105 (
            .O(N__32472),
            .I(N__32469));
    Odrv4 I__3104 (
            .O(N__32469),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__3103 (
            .O(N__32466),
            .I(\pid_alt.un2_pid_prereg_cry_14 ));
    InMux I__3102 (
            .O(N__32463),
            .I(N__32460));
    LocalMux I__3101 (
            .O(N__32460),
            .I(N__32457));
    Span4Mux_v I__3100 (
            .O(N__32457),
            .I(N__32454));
    Odrv4 I__3099 (
            .O(N__32454),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__3098 (
            .O(N__32451),
            .I(bfn_2_14_0_));
    InMux I__3097 (
            .O(N__32448),
            .I(N__32445));
    LocalMux I__3096 (
            .O(N__32445),
            .I(N__32442));
    Odrv4 I__3095 (
            .O(N__32442),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__3094 (
            .O(N__32439),
            .I(\pid_alt.un2_pid_prereg_cry_16 ));
    InMux I__3093 (
            .O(N__32436),
            .I(N__32433));
    LocalMux I__3092 (
            .O(N__32433),
            .I(N__32430));
    Span4Mux_v I__3091 (
            .O(N__32430),
            .I(N__32427));
    Odrv4 I__3090 (
            .O(N__32427),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__3089 (
            .O(N__32424),
            .I(\pid_alt.un2_pid_prereg_cry_17 ));
    InMux I__3088 (
            .O(N__32421),
            .I(N__32418));
    LocalMux I__3087 (
            .O(N__32418),
            .I(N__32415));
    Span4Mux_v I__3086 (
            .O(N__32415),
            .I(N__32412));
    Odrv4 I__3085 (
            .O(N__32412),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__3084 (
            .O(N__32409),
            .I(\pid_alt.un2_pid_prereg_cry_18 ));
    InMux I__3083 (
            .O(N__32406),
            .I(\pid_alt.un2_pid_prereg_cry_19 ));
    CascadeMux I__3082 (
            .O(N__32403),
            .I(N__32400));
    InMux I__3081 (
            .O(N__32400),
            .I(N__32397));
    LocalMux I__3080 (
            .O(N__32397),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__3079 (
            .O(N__32394),
            .I(\pid_alt.un2_pid_prereg_cry_3 ));
    CascadeMux I__3078 (
            .O(N__32391),
            .I(N__32388));
    InMux I__3077 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__3076 (
            .O(N__32385),
            .I(N__32382));
    Odrv4 I__3075 (
            .O(N__32382),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__3074 (
            .O(N__32379),
            .I(\pid_alt.un2_pid_prereg_cry_4 ));
    InMux I__3073 (
            .O(N__32376),
            .I(N__32372));
    InMux I__3072 (
            .O(N__32375),
            .I(N__32369));
    LocalMux I__3071 (
            .O(N__32372),
            .I(N__32366));
    LocalMux I__3070 (
            .O(N__32369),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__3069 (
            .O(N__32366),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    CascadeMux I__3068 (
            .O(N__32361),
            .I(N__32358));
    InMux I__3067 (
            .O(N__32358),
            .I(N__32355));
    LocalMux I__3066 (
            .O(N__32355),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__3065 (
            .O(N__32352),
            .I(\pid_alt.un2_pid_prereg_cry_5 ));
    CascadeMux I__3064 (
            .O(N__32349),
            .I(N__32345));
    InMux I__3063 (
            .O(N__32348),
            .I(N__32342));
    InMux I__3062 (
            .O(N__32345),
            .I(N__32339));
    LocalMux I__3061 (
            .O(N__32342),
            .I(N__32336));
    LocalMux I__3060 (
            .O(N__32339),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv12 I__3059 (
            .O(N__32336),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    CascadeMux I__3058 (
            .O(N__32331),
            .I(N__32328));
    InMux I__3057 (
            .O(N__32328),
            .I(N__32325));
    LocalMux I__3056 (
            .O(N__32325),
            .I(N__32322));
    Span4Mux_h I__3055 (
            .O(N__32322),
            .I(N__32319));
    Odrv4 I__3054 (
            .O(N__32319),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__3053 (
            .O(N__32316),
            .I(\pid_alt.un2_pid_prereg_cry_6 ));
    CascadeMux I__3052 (
            .O(N__32313),
            .I(N__32310));
    InMux I__3051 (
            .O(N__32310),
            .I(N__32306));
    InMux I__3050 (
            .O(N__32309),
            .I(N__32303));
    LocalMux I__3049 (
            .O(N__32306),
            .I(N__32298));
    LocalMux I__3048 (
            .O(N__32303),
            .I(N__32298));
    Odrv4 I__3047 (
            .O(N__32298),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    CascadeMux I__3046 (
            .O(N__32295),
            .I(N__32292));
    InMux I__3045 (
            .O(N__32292),
            .I(N__32289));
    LocalMux I__3044 (
            .O(N__32289),
            .I(N__32286));
    Odrv4 I__3043 (
            .O(N__32286),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__3042 (
            .O(N__32283),
            .I(bfn_2_13_0_));
    CascadeMux I__3041 (
            .O(N__32280),
            .I(N__32276));
    InMux I__3040 (
            .O(N__32279),
            .I(N__32273));
    InMux I__3039 (
            .O(N__32276),
            .I(N__32270));
    LocalMux I__3038 (
            .O(N__32273),
            .I(N__32267));
    LocalMux I__3037 (
            .O(N__32270),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    Odrv4 I__3036 (
            .O(N__32267),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    CascadeMux I__3035 (
            .O(N__32262),
            .I(N__32259));
    InMux I__3034 (
            .O(N__32259),
            .I(N__32256));
    LocalMux I__3033 (
            .O(N__32256),
            .I(N__32253));
    Span4Mux_v I__3032 (
            .O(N__32253),
            .I(N__32250));
    Odrv4 I__3031 (
            .O(N__32250),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__3030 (
            .O(N__32247),
            .I(\pid_alt.un2_pid_prereg_cry_8 ));
    CascadeMux I__3029 (
            .O(N__32244),
            .I(N__32240));
    InMux I__3028 (
            .O(N__32243),
            .I(N__32237));
    InMux I__3027 (
            .O(N__32240),
            .I(N__32234));
    LocalMux I__3026 (
            .O(N__32237),
            .I(N__32231));
    LocalMux I__3025 (
            .O(N__32234),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv12 I__3024 (
            .O(N__32231),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    CascadeMux I__3023 (
            .O(N__32226),
            .I(N__32223));
    InMux I__3022 (
            .O(N__32223),
            .I(N__32220));
    LocalMux I__3021 (
            .O(N__32220),
            .I(N__32217));
    Odrv4 I__3020 (
            .O(N__32217),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__3019 (
            .O(N__32214),
            .I(\pid_alt.un2_pid_prereg_cry_9 ));
    InMux I__3018 (
            .O(N__32211),
            .I(N__32207));
    CascadeMux I__3017 (
            .O(N__32210),
            .I(N__32204));
    LocalMux I__3016 (
            .O(N__32207),
            .I(N__32201));
    InMux I__3015 (
            .O(N__32204),
            .I(N__32198));
    Span4Mux_v I__3014 (
            .O(N__32201),
            .I(N__32195));
    LocalMux I__3013 (
            .O(N__32198),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv4 I__3012 (
            .O(N__32195),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    CascadeMux I__3011 (
            .O(N__32190),
            .I(N__32187));
    InMux I__3010 (
            .O(N__32187),
            .I(N__32184));
    LocalMux I__3009 (
            .O(N__32184),
            .I(N__32181));
    Span4Mux_v I__3008 (
            .O(N__32181),
            .I(N__32178));
    Odrv4 I__3007 (
            .O(N__32178),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__3006 (
            .O(N__32175),
            .I(\pid_alt.un2_pid_prereg_cry_10 ));
    InMux I__3005 (
            .O(N__32172),
            .I(N__32169));
    LocalMux I__3004 (
            .O(N__32169),
            .I(\pid_alt.m35_e_2 ));
    CascadeMux I__3003 (
            .O(N__32166),
            .I(\pid_alt.N_62_mux_cascade_ ));
    CascadeMux I__3002 (
            .O(N__32163),
            .I(\pid_alt.N_94_cascade_ ));
    InMux I__3001 (
            .O(N__32160),
            .I(N__32151));
    InMux I__3000 (
            .O(N__32159),
            .I(N__32151));
    InMux I__2999 (
            .O(N__32158),
            .I(N__32151));
    LocalMux I__2998 (
            .O(N__32151),
            .I(\pid_alt.N_94 ));
    InMux I__2997 (
            .O(N__32148),
            .I(N__32145));
    LocalMux I__2996 (
            .O(N__32145),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    CascadeMux I__2995 (
            .O(N__32142),
            .I(N__32139));
    InMux I__2994 (
            .O(N__32139),
            .I(N__32136));
    LocalMux I__2993 (
            .O(N__32136),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__2992 (
            .O(N__32133),
            .I(\pid_alt.un2_pid_prereg_cry_0 ));
    InMux I__2991 (
            .O(N__32130),
            .I(N__32127));
    LocalMux I__2990 (
            .O(N__32127),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    CascadeMux I__2989 (
            .O(N__32124),
            .I(N__32121));
    InMux I__2988 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__2987 (
            .O(N__32118),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    InMux I__2986 (
            .O(N__32115),
            .I(\pid_alt.un2_pid_prereg_cry_1 ));
    InMux I__2985 (
            .O(N__32112),
            .I(N__32109));
    LocalMux I__2984 (
            .O(N__32109),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    CascadeMux I__2983 (
            .O(N__32106),
            .I(N__32103));
    InMux I__2982 (
            .O(N__32103),
            .I(N__32100));
    LocalMux I__2981 (
            .O(N__32100),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__2980 (
            .O(N__32097),
            .I(\pid_alt.un2_pid_prereg_cry_2 ));
    InMux I__2979 (
            .O(N__32094),
            .I(N__32091));
    LocalMux I__2978 (
            .O(N__32091),
            .I(N__32088));
    Odrv12 I__2977 (
            .O(N__32088),
            .I(alt_kd_4));
    InMux I__2976 (
            .O(N__32085),
            .I(N__32082));
    LocalMux I__2975 (
            .O(N__32082),
            .I(N__32079));
    Odrv12 I__2974 (
            .O(N__32079),
            .I(alt_kd_6));
    InMux I__2973 (
            .O(N__32076),
            .I(N__32073));
    LocalMux I__2972 (
            .O(N__32073),
            .I(N__32070));
    Span4Mux_s3_h I__2971 (
            .O(N__32070),
            .I(N__32067));
    Odrv4 I__2970 (
            .O(N__32067),
            .I(alt_kd_3));
    InMux I__2969 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__2968 (
            .O(N__32061),
            .I(N__32058));
    Odrv4 I__2967 (
            .O(N__32058),
            .I(\pid_alt.O_5_16 ));
    InMux I__2966 (
            .O(N__32055),
            .I(N__32052));
    LocalMux I__2965 (
            .O(N__32052),
            .I(\pid_alt.O_5_8 ));
    InMux I__2964 (
            .O(N__32049),
            .I(N__32046));
    LocalMux I__2963 (
            .O(N__32046),
            .I(\pid_alt.O_5_15 ));
    InMux I__2962 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__2961 (
            .O(N__32040),
            .I(\pid_alt.O_5_10 ));
    InMux I__2960 (
            .O(N__32037),
            .I(N__32031));
    InMux I__2959 (
            .O(N__32036),
            .I(N__32031));
    LocalMux I__2958 (
            .O(N__32031),
            .I(N__32028));
    Span12Mux_v I__2957 (
            .O(N__32028),
            .I(N__32025));
    Odrv12 I__2956 (
            .O(N__32025),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__2955 (
            .O(N__32022),
            .I(N__32019));
    LocalMux I__2954 (
            .O(N__32019),
            .I(N__32016));
    Span4Mux_s2_h I__2953 (
            .O(N__32016),
            .I(N__32013));
    Odrv4 I__2952 (
            .O(N__32013),
            .I(alt_kd_1));
    InMux I__2951 (
            .O(N__32010),
            .I(N__32007));
    LocalMux I__2950 (
            .O(N__32007),
            .I(N__32004));
    Span4Mux_s2_h I__2949 (
            .O(N__32004),
            .I(N__32001));
    Odrv4 I__2948 (
            .O(N__32001),
            .I(alt_kd_2));
    InMux I__2947 (
            .O(N__31998),
            .I(N__31995));
    LocalMux I__2946 (
            .O(N__31995),
            .I(N__31992));
    Span4Mux_v I__2945 (
            .O(N__31992),
            .I(N__31989));
    Odrv4 I__2944 (
            .O(N__31989),
            .I(alt_kd_0));
    InMux I__2943 (
            .O(N__31986),
            .I(N__31983));
    LocalMux I__2942 (
            .O(N__31983),
            .I(N__31980));
    Span4Mux_v I__2941 (
            .O(N__31980),
            .I(N__31977));
    Odrv4 I__2940 (
            .O(N__31977),
            .I(alt_kd_5));
    InMux I__2939 (
            .O(N__31974),
            .I(N__31971));
    LocalMux I__2938 (
            .O(N__31971),
            .I(N__31968));
    Span4Mux_s2_h I__2937 (
            .O(N__31968),
            .I(N__31965));
    Odrv4 I__2936 (
            .O(N__31965),
            .I(alt_kd_7));
    InMux I__2935 (
            .O(N__31962),
            .I(N__31959));
    LocalMux I__2934 (
            .O(N__31959),
            .I(N__31956));
    Span4Mux_h I__2933 (
            .O(N__31956),
            .I(N__31953));
    Odrv4 I__2932 (
            .O(N__31953),
            .I(\pid_alt.O_5_14 ));
    InMux I__2931 (
            .O(N__31950),
            .I(N__31947));
    LocalMux I__2930 (
            .O(N__31947),
            .I(N__31944));
    Span4Mux_h I__2929 (
            .O(N__31944),
            .I(N__31941));
    Odrv4 I__2928 (
            .O(N__31941),
            .I(\pid_alt.O_5_24 ));
    InMux I__2927 (
            .O(N__31938),
            .I(N__31935));
    LocalMux I__2926 (
            .O(N__31935),
            .I(N__31932));
    Span4Mux_h I__2925 (
            .O(N__31932),
            .I(N__31929));
    Odrv4 I__2924 (
            .O(N__31929),
            .I(\pid_alt.O_5_17 ));
    InMux I__2923 (
            .O(N__31926),
            .I(N__31923));
    LocalMux I__2922 (
            .O(N__31923),
            .I(N__31920));
    Odrv4 I__2921 (
            .O(N__31920),
            .I(\pid_alt.O_5_18 ));
    InMux I__2920 (
            .O(N__31917),
            .I(N__31914));
    LocalMux I__2919 (
            .O(N__31914),
            .I(N__31911));
    Span4Mux_h I__2918 (
            .O(N__31911),
            .I(N__31908));
    Odrv4 I__2917 (
            .O(N__31908),
            .I(\pid_alt.O_5_19 ));
    InMux I__2916 (
            .O(N__31905),
            .I(N__31902));
    LocalMux I__2915 (
            .O(N__31902),
            .I(N__31899));
    Odrv4 I__2914 (
            .O(N__31899),
            .I(\pid_alt.O_5_20 ));
    InMux I__2913 (
            .O(N__31896),
            .I(N__31893));
    LocalMux I__2912 (
            .O(N__31893),
            .I(N__31890));
    Odrv4 I__2911 (
            .O(N__31890),
            .I(\pid_alt.O_5_21 ));
    InMux I__2910 (
            .O(N__31887),
            .I(N__31884));
    LocalMux I__2909 (
            .O(N__31884),
            .I(N__31881));
    Odrv4 I__2908 (
            .O(N__31881),
            .I(\pid_alt.O_5_22 ));
    InMux I__2907 (
            .O(N__31878),
            .I(N__31875));
    LocalMux I__2906 (
            .O(N__31875),
            .I(N__31872));
    Odrv4 I__2905 (
            .O(N__31872),
            .I(\pid_alt.O_5_23 ));
    InMux I__2904 (
            .O(N__31869),
            .I(N__31863));
    InMux I__2903 (
            .O(N__31868),
            .I(N__31863));
    LocalMux I__2902 (
            .O(N__31863),
            .I(N__31860));
    Odrv12 I__2901 (
            .O(N__31860),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    InMux I__2900 (
            .O(N__31857),
            .I(\pid_alt.error_cry_14 ));
    InMux I__2899 (
            .O(N__31854),
            .I(N__31851));
    LocalMux I__2898 (
            .O(N__31851),
            .I(N__31848));
    Span4Mux_s1_h I__2897 (
            .O(N__31848),
            .I(N__31843));
    InMux I__2896 (
            .O(N__31847),
            .I(N__31840));
    InMux I__2895 (
            .O(N__31846),
            .I(N__31837));
    Span4Mux_v I__2894 (
            .O(N__31843),
            .I(N__31832));
    LocalMux I__2893 (
            .O(N__31840),
            .I(N__31832));
    LocalMux I__2892 (
            .O(N__31837),
            .I(N__31829));
    Span4Mux_v I__2891 (
            .O(N__31832),
            .I(N__31826));
    Span4Mux_v I__2890 (
            .O(N__31829),
            .I(N__31823));
    Odrv4 I__2889 (
            .O(N__31826),
            .I(\pid_alt.error_15 ));
    Odrv4 I__2888 (
            .O(N__31823),
            .I(\pid_alt.error_15 ));
    CascadeMux I__2887 (
            .O(N__31818),
            .I(N__31815));
    InMux I__2886 (
            .O(N__31815),
            .I(N__31812));
    LocalMux I__2885 (
            .O(N__31812),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__2884 (
            .O(N__31809),
            .I(N__31806));
    LocalMux I__2883 (
            .O(N__31806),
            .I(N__31803));
    Odrv4 I__2882 (
            .O(N__31803),
            .I(drone_altitude_i_5));
    InMux I__2881 (
            .O(N__31800),
            .I(N__31797));
    LocalMux I__2880 (
            .O(N__31797),
            .I(N__31794));
    Odrv4 I__2879 (
            .O(N__31794),
            .I(drone_altitude_i_6));
    CascadeMux I__2878 (
            .O(N__31791),
            .I(N__31788));
    InMux I__2877 (
            .O(N__31788),
            .I(N__31785));
    LocalMux I__2876 (
            .O(N__31785),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__2875 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__2874 (
            .O(N__31779),
            .I(N__31776));
    Odrv4 I__2873 (
            .O(N__31776),
            .I(\pid_alt.O_5_9 ));
    InMux I__2872 (
            .O(N__31773),
            .I(N__31770));
    LocalMux I__2871 (
            .O(N__31770),
            .I(N__31766));
    InMux I__2870 (
            .O(N__31769),
            .I(N__31762));
    Span4Mux_s1_h I__2869 (
            .O(N__31766),
            .I(N__31759));
    InMux I__2868 (
            .O(N__31765),
            .I(N__31756));
    LocalMux I__2867 (
            .O(N__31762),
            .I(N__31753));
    Span4Mux_v I__2866 (
            .O(N__31759),
            .I(N__31748));
    LocalMux I__2865 (
            .O(N__31756),
            .I(N__31748));
    Span4Mux_v I__2864 (
            .O(N__31753),
            .I(N__31745));
    Span4Mux_v I__2863 (
            .O(N__31748),
            .I(N__31740));
    Span4Mux_v I__2862 (
            .O(N__31745),
            .I(N__31740));
    Odrv4 I__2861 (
            .O(N__31740),
            .I(\pid_alt.error_7 ));
    InMux I__2860 (
            .O(N__31737),
            .I(\pid_alt.error_cry_6 ));
    InMux I__2859 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__2858 (
            .O(N__31731),
            .I(N__31726));
    InMux I__2857 (
            .O(N__31730),
            .I(N__31723));
    InMux I__2856 (
            .O(N__31729),
            .I(N__31720));
    Span4Mux_v I__2855 (
            .O(N__31726),
            .I(N__31717));
    LocalMux I__2854 (
            .O(N__31723),
            .I(N__31714));
    LocalMux I__2853 (
            .O(N__31720),
            .I(N__31711));
    Span4Mux_v I__2852 (
            .O(N__31717),
            .I(N__31706));
    Span4Mux_v I__2851 (
            .O(N__31714),
            .I(N__31706));
    Span4Mux_v I__2850 (
            .O(N__31711),
            .I(N__31703));
    Span4Mux_v I__2849 (
            .O(N__31706),
            .I(N__31698));
    Span4Mux_v I__2848 (
            .O(N__31703),
            .I(N__31698));
    Odrv4 I__2847 (
            .O(N__31698),
            .I(\pid_alt.error_8 ));
    InMux I__2846 (
            .O(N__31695),
            .I(bfn_1_18_0_));
    InMux I__2845 (
            .O(N__31692),
            .I(N__31688));
    InMux I__2844 (
            .O(N__31691),
            .I(N__31684));
    LocalMux I__2843 (
            .O(N__31688),
            .I(N__31681));
    InMux I__2842 (
            .O(N__31687),
            .I(N__31678));
    LocalMux I__2841 (
            .O(N__31684),
            .I(N__31675));
    Span4Mux_v I__2840 (
            .O(N__31681),
            .I(N__31672));
    LocalMux I__2839 (
            .O(N__31678),
            .I(N__31669));
    Span12Mux_s1_h I__2838 (
            .O(N__31675),
            .I(N__31666));
    Sp12to4 I__2837 (
            .O(N__31672),
            .I(N__31661));
    Sp12to4 I__2836 (
            .O(N__31669),
            .I(N__31661));
    Odrv12 I__2835 (
            .O(N__31666),
            .I(\pid_alt.error_9 ));
    Odrv12 I__2834 (
            .O(N__31661),
            .I(\pid_alt.error_9 ));
    InMux I__2833 (
            .O(N__31656),
            .I(\pid_alt.error_cry_8 ));
    InMux I__2832 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__2831 (
            .O(N__31650),
            .I(N__31647));
    Span4Mux_s1_h I__2830 (
            .O(N__31647),
            .I(N__31642));
    InMux I__2829 (
            .O(N__31646),
            .I(N__31639));
    InMux I__2828 (
            .O(N__31645),
            .I(N__31636));
    Span4Mux_v I__2827 (
            .O(N__31642),
            .I(N__31631));
    LocalMux I__2826 (
            .O(N__31639),
            .I(N__31631));
    LocalMux I__2825 (
            .O(N__31636),
            .I(N__31628));
    Span4Mux_v I__2824 (
            .O(N__31631),
            .I(N__31625));
    Span4Mux_v I__2823 (
            .O(N__31628),
            .I(N__31622));
    Odrv4 I__2822 (
            .O(N__31625),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2821 (
            .O(N__31622),
            .I(\pid_alt.error_10 ));
    InMux I__2820 (
            .O(N__31617),
            .I(\pid_alt.error_cry_9 ));
    InMux I__2819 (
            .O(N__31614),
            .I(N__31611));
    LocalMux I__2818 (
            .O(N__31611),
            .I(N__31608));
    Span4Mux_v I__2817 (
            .O(N__31608),
            .I(N__31603));
    InMux I__2816 (
            .O(N__31607),
            .I(N__31600));
    InMux I__2815 (
            .O(N__31606),
            .I(N__31597));
    Span4Mux_s1_h I__2814 (
            .O(N__31603),
            .I(N__31592));
    LocalMux I__2813 (
            .O(N__31600),
            .I(N__31592));
    LocalMux I__2812 (
            .O(N__31597),
            .I(N__31589));
    Sp12to4 I__2811 (
            .O(N__31592),
            .I(N__31586));
    Sp12to4 I__2810 (
            .O(N__31589),
            .I(N__31583));
    Odrv12 I__2809 (
            .O(N__31586),
            .I(\pid_alt.error_11 ));
    Odrv12 I__2808 (
            .O(N__31583),
            .I(\pid_alt.error_11 ));
    InMux I__2807 (
            .O(N__31578),
            .I(\pid_alt.error_cry_10 ));
    InMux I__2806 (
            .O(N__31575),
            .I(N__31571));
    InMux I__2805 (
            .O(N__31574),
            .I(N__31567));
    LocalMux I__2804 (
            .O(N__31571),
            .I(N__31564));
    InMux I__2803 (
            .O(N__31570),
            .I(N__31561));
    LocalMux I__2802 (
            .O(N__31567),
            .I(N__31558));
    Span4Mux_v I__2801 (
            .O(N__31564),
            .I(N__31553));
    LocalMux I__2800 (
            .O(N__31561),
            .I(N__31553));
    Span4Mux_s1_h I__2799 (
            .O(N__31558),
            .I(N__31550));
    Span4Mux_v I__2798 (
            .O(N__31553),
            .I(N__31547));
    Span4Mux_v I__2797 (
            .O(N__31550),
            .I(N__31544));
    Odrv4 I__2796 (
            .O(N__31547),
            .I(\pid_alt.error_12 ));
    Odrv4 I__2795 (
            .O(N__31544),
            .I(\pid_alt.error_12 ));
    InMux I__2794 (
            .O(N__31539),
            .I(\pid_alt.error_cry_11 ));
    InMux I__2793 (
            .O(N__31536),
            .I(N__31533));
    LocalMux I__2792 (
            .O(N__31533),
            .I(N__31528));
    InMux I__2791 (
            .O(N__31532),
            .I(N__31525));
    InMux I__2790 (
            .O(N__31531),
            .I(N__31522));
    Span4Mux_v I__2789 (
            .O(N__31528),
            .I(N__31517));
    LocalMux I__2788 (
            .O(N__31525),
            .I(N__31517));
    LocalMux I__2787 (
            .O(N__31522),
            .I(N__31514));
    Span4Mux_v I__2786 (
            .O(N__31517),
            .I(N__31511));
    Span4Mux_v I__2785 (
            .O(N__31514),
            .I(N__31508));
    Odrv4 I__2784 (
            .O(N__31511),
            .I(\pid_alt.error_13 ));
    Odrv4 I__2783 (
            .O(N__31508),
            .I(\pid_alt.error_13 ));
    InMux I__2782 (
            .O(N__31503),
            .I(\pid_alt.error_cry_12 ));
    InMux I__2781 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__2780 (
            .O(N__31497),
            .I(N__31494));
    Span4Mux_s1_h I__2779 (
            .O(N__31494),
            .I(N__31489));
    InMux I__2778 (
            .O(N__31493),
            .I(N__31486));
    InMux I__2777 (
            .O(N__31492),
            .I(N__31483));
    Span4Mux_v I__2776 (
            .O(N__31489),
            .I(N__31478));
    LocalMux I__2775 (
            .O(N__31486),
            .I(N__31478));
    LocalMux I__2774 (
            .O(N__31483),
            .I(N__31475));
    Span4Mux_v I__2773 (
            .O(N__31478),
            .I(N__31472));
    Span4Mux_v I__2772 (
            .O(N__31475),
            .I(N__31469));
    Odrv4 I__2771 (
            .O(N__31472),
            .I(\pid_alt.error_14 ));
    Odrv4 I__2770 (
            .O(N__31469),
            .I(\pid_alt.error_14 ));
    InMux I__2769 (
            .O(N__31464),
            .I(\pid_alt.error_cry_13 ));
    InMux I__2768 (
            .O(N__31461),
            .I(N__31458));
    LocalMux I__2767 (
            .O(N__31458),
            .I(\pid_front.O_0_22 ));
    InMux I__2766 (
            .O(N__31455),
            .I(N__31452));
    LocalMux I__2765 (
            .O(N__31452),
            .I(\pid_front.O_0_9 ));
    InMux I__2764 (
            .O(N__31449),
            .I(N__31446));
    LocalMux I__2763 (
            .O(N__31446),
            .I(N__31443));
    Span4Mux_s1_h I__2762 (
            .O(N__31443),
            .I(N__31438));
    InMux I__2761 (
            .O(N__31442),
            .I(N__31435));
    InMux I__2760 (
            .O(N__31441),
            .I(N__31432));
    Span4Mux_v I__2759 (
            .O(N__31438),
            .I(N__31427));
    LocalMux I__2758 (
            .O(N__31435),
            .I(N__31427));
    LocalMux I__2757 (
            .O(N__31432),
            .I(N__31424));
    Span4Mux_v I__2756 (
            .O(N__31427),
            .I(N__31421));
    Sp12to4 I__2755 (
            .O(N__31424),
            .I(N__31418));
    Odrv4 I__2754 (
            .O(N__31421),
            .I(\pid_alt.error_1 ));
    Odrv12 I__2753 (
            .O(N__31418),
            .I(\pid_alt.error_1 ));
    InMux I__2752 (
            .O(N__31413),
            .I(\pid_alt.error_cry_0 ));
    InMux I__2751 (
            .O(N__31410),
            .I(N__31405));
    InMux I__2750 (
            .O(N__31409),
            .I(N__31402));
    InMux I__2749 (
            .O(N__31408),
            .I(N__31399));
    LocalMux I__2748 (
            .O(N__31405),
            .I(N__31396));
    LocalMux I__2747 (
            .O(N__31402),
            .I(N__31393));
    LocalMux I__2746 (
            .O(N__31399),
            .I(N__31390));
    Span4Mux_v I__2745 (
            .O(N__31396),
            .I(N__31387));
    Span4Mux_v I__2744 (
            .O(N__31393),
            .I(N__31384));
    Span12Mux_s1_h I__2743 (
            .O(N__31390),
            .I(N__31381));
    Span4Mux_v I__2742 (
            .O(N__31387),
            .I(N__31376));
    Span4Mux_v I__2741 (
            .O(N__31384),
            .I(N__31376));
    Odrv12 I__2740 (
            .O(N__31381),
            .I(\pid_alt.error_2 ));
    Odrv4 I__2739 (
            .O(N__31376),
            .I(\pid_alt.error_2 ));
    InMux I__2738 (
            .O(N__31371),
            .I(\pid_alt.error_cry_1 ));
    InMux I__2737 (
            .O(N__31368),
            .I(N__31365));
    LocalMux I__2736 (
            .O(N__31365),
            .I(N__31360));
    InMux I__2735 (
            .O(N__31364),
            .I(N__31357));
    InMux I__2734 (
            .O(N__31363),
            .I(N__31354));
    Span4Mux_v I__2733 (
            .O(N__31360),
            .I(N__31349));
    LocalMux I__2732 (
            .O(N__31357),
            .I(N__31349));
    LocalMux I__2731 (
            .O(N__31354),
            .I(N__31346));
    Span4Mux_v I__2730 (
            .O(N__31349),
            .I(N__31343));
    Span4Mux_v I__2729 (
            .O(N__31346),
            .I(N__31340));
    Span4Mux_v I__2728 (
            .O(N__31343),
            .I(N__31335));
    Span4Mux_v I__2727 (
            .O(N__31340),
            .I(N__31335));
    Odrv4 I__2726 (
            .O(N__31335),
            .I(\pid_alt.error_3 ));
    InMux I__2725 (
            .O(N__31332),
            .I(\pid_alt.error_cry_2 ));
    InMux I__2724 (
            .O(N__31329),
            .I(N__31324));
    InMux I__2723 (
            .O(N__31328),
            .I(N__31321));
    InMux I__2722 (
            .O(N__31327),
            .I(N__31318));
    LocalMux I__2721 (
            .O(N__31324),
            .I(N__31315));
    LocalMux I__2720 (
            .O(N__31321),
            .I(N__31312));
    LocalMux I__2719 (
            .O(N__31318),
            .I(N__31309));
    Span4Mux_v I__2718 (
            .O(N__31315),
            .I(N__31306));
    Span4Mux_s1_h I__2717 (
            .O(N__31312),
            .I(N__31303));
    Span4Mux_v I__2716 (
            .O(N__31309),
            .I(N__31300));
    Span4Mux_v I__2715 (
            .O(N__31306),
            .I(N__31297));
    Span4Mux_v I__2714 (
            .O(N__31303),
            .I(N__31292));
    Span4Mux_v I__2713 (
            .O(N__31300),
            .I(N__31292));
    Odrv4 I__2712 (
            .O(N__31297),
            .I(\pid_alt.error_4 ));
    Odrv4 I__2711 (
            .O(N__31292),
            .I(\pid_alt.error_4 ));
    InMux I__2710 (
            .O(N__31287),
            .I(\pid_alt.error_cry_3 ));
    InMux I__2709 (
            .O(N__31284),
            .I(N__31281));
    LocalMux I__2708 (
            .O(N__31281),
            .I(N__31278));
    Span4Mux_v I__2707 (
            .O(N__31278),
            .I(N__31273));
    InMux I__2706 (
            .O(N__31277),
            .I(N__31270));
    InMux I__2705 (
            .O(N__31276),
            .I(N__31267));
    Span4Mux_v I__2704 (
            .O(N__31273),
            .I(N__31262));
    LocalMux I__2703 (
            .O(N__31270),
            .I(N__31262));
    LocalMux I__2702 (
            .O(N__31267),
            .I(N__31259));
    Span4Mux_s1_h I__2701 (
            .O(N__31262),
            .I(N__31256));
    Span4Mux_v I__2700 (
            .O(N__31259),
            .I(N__31253));
    Span4Mux_v I__2699 (
            .O(N__31256),
            .I(N__31248));
    Span4Mux_v I__2698 (
            .O(N__31253),
            .I(N__31248));
    Odrv4 I__2697 (
            .O(N__31248),
            .I(\pid_alt.error_5 ));
    InMux I__2696 (
            .O(N__31245),
            .I(\pid_alt.error_cry_4 ));
    InMux I__2695 (
            .O(N__31242),
            .I(N__31239));
    LocalMux I__2694 (
            .O(N__31239),
            .I(N__31234));
    InMux I__2693 (
            .O(N__31238),
            .I(N__31231));
    InMux I__2692 (
            .O(N__31237),
            .I(N__31228));
    Span4Mux_v I__2691 (
            .O(N__31234),
            .I(N__31223));
    LocalMux I__2690 (
            .O(N__31231),
            .I(N__31223));
    LocalMux I__2689 (
            .O(N__31228),
            .I(N__31220));
    Span4Mux_v I__2688 (
            .O(N__31223),
            .I(N__31217));
    Span4Mux_v I__2687 (
            .O(N__31220),
            .I(N__31214));
    Span4Mux_v I__2686 (
            .O(N__31217),
            .I(N__31209));
    Span4Mux_v I__2685 (
            .O(N__31214),
            .I(N__31209));
    Odrv4 I__2684 (
            .O(N__31209),
            .I(\pid_alt.error_6 ));
    InMux I__2683 (
            .O(N__31206),
            .I(\pid_alt.error_cry_5 ));
    InMux I__2682 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__2681 (
            .O(N__31200),
            .I(\pid_front.O_0_5 ));
    InMux I__2680 (
            .O(N__31197),
            .I(N__31194));
    LocalMux I__2679 (
            .O(N__31194),
            .I(\pid_front.O_0_10 ));
    InMux I__2678 (
            .O(N__31191),
            .I(N__31188));
    LocalMux I__2677 (
            .O(N__31188),
            .I(\pid_front.O_0_11 ));
    InMux I__2676 (
            .O(N__31185),
            .I(N__31182));
    LocalMux I__2675 (
            .O(N__31182),
            .I(\pid_front.O_0_16 ));
    InMux I__2674 (
            .O(N__31179),
            .I(N__31176));
    LocalMux I__2673 (
            .O(N__31176),
            .I(\pid_front.O_0_17 ));
    InMux I__2672 (
            .O(N__31173),
            .I(N__31170));
    LocalMux I__2671 (
            .O(N__31170),
            .I(\pid_front.O_0_18 ));
    InMux I__2670 (
            .O(N__31167),
            .I(N__31164));
    LocalMux I__2669 (
            .O(N__31164),
            .I(\pid_front.O_0_19 ));
    InMux I__2668 (
            .O(N__31161),
            .I(N__31158));
    LocalMux I__2667 (
            .O(N__31158),
            .I(\pid_front.O_0_20 ));
    InMux I__2666 (
            .O(N__31155),
            .I(N__31152));
    LocalMux I__2665 (
            .O(N__31152),
            .I(\pid_front.O_0_21 ));
    InMux I__2664 (
            .O(N__31149),
            .I(N__31146));
    LocalMux I__2663 (
            .O(N__31146),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    InMux I__2662 (
            .O(N__31143),
            .I(N__31137));
    InMux I__2661 (
            .O(N__31142),
            .I(N__31137));
    LocalMux I__2660 (
            .O(N__31137),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    InMux I__2659 (
            .O(N__31134),
            .I(N__31128));
    InMux I__2658 (
            .O(N__31133),
            .I(N__31128));
    LocalMux I__2657 (
            .O(N__31128),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    InMux I__2656 (
            .O(N__31125),
            .I(N__31116));
    InMux I__2655 (
            .O(N__31124),
            .I(N__31116));
    InMux I__2654 (
            .O(N__31123),
            .I(N__31116));
    LocalMux I__2653 (
            .O(N__31116),
            .I(N__31113));
    Odrv12 I__2652 (
            .O(N__31113),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    InMux I__2651 (
            .O(N__31110),
            .I(N__31107));
    LocalMux I__2650 (
            .O(N__31107),
            .I(N__31104));
    Odrv4 I__2649 (
            .O(N__31104),
            .I(\pid_front.O_0_23 ));
    InMux I__2648 (
            .O(N__31101),
            .I(N__31098));
    LocalMux I__2647 (
            .O(N__31098),
            .I(N__31095));
    Odrv4 I__2646 (
            .O(N__31095),
            .I(\pid_front.O_0_24 ));
    InMux I__2645 (
            .O(N__31092),
            .I(N__31089));
    LocalMux I__2644 (
            .O(N__31089),
            .I(\pid_front.O_0_12 ));
    InMux I__2643 (
            .O(N__31086),
            .I(N__31083));
    LocalMux I__2642 (
            .O(N__31083),
            .I(\pid_front.O_0_7 ));
    InMux I__2641 (
            .O(N__31080),
            .I(N__31077));
    LocalMux I__2640 (
            .O(N__31077),
            .I(\pid_front.O_0_8 ));
    InMux I__2639 (
            .O(N__31074),
            .I(N__31071));
    LocalMux I__2638 (
            .O(N__31071),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__2637 (
            .O(N__31068),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ));
    CascadeMux I__2636 (
            .O(N__31065),
            .I(N__31061));
    InMux I__2635 (
            .O(N__31064),
            .I(N__31056));
    InMux I__2634 (
            .O(N__31061),
            .I(N__31056));
    LocalMux I__2633 (
            .O(N__31056),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    InMux I__2632 (
            .O(N__31053),
            .I(N__31044));
    InMux I__2631 (
            .O(N__31052),
            .I(N__31044));
    InMux I__2630 (
            .O(N__31051),
            .I(N__31044));
    LocalMux I__2629 (
            .O(N__31044),
            .I(N__31041));
    Span12Mux_v I__2628 (
            .O(N__31041),
            .I(N__31038));
    Odrv12 I__2627 (
            .O(N__31038),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    CascadeMux I__2626 (
            .O(N__31035),
            .I(N__31032));
    InMux I__2625 (
            .O(N__31032),
            .I(N__31026));
    InMux I__2624 (
            .O(N__31031),
            .I(N__31026));
    LocalMux I__2623 (
            .O(N__31026),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    CascadeMux I__2622 (
            .O(N__31023),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6_cascade_ ));
    CascadeMux I__2621 (
            .O(N__31020),
            .I(\pid_alt.un1_pid_prereg_236_1_cascade_ ));
    InMux I__2620 (
            .O(N__31017),
            .I(N__31014));
    LocalMux I__2619 (
            .O(N__31014),
            .I(\pid_alt.O_4_20 ));
    InMux I__2618 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__2617 (
            .O(N__31008),
            .I(\pid_alt.O_4_15 ));
    InMux I__2616 (
            .O(N__31005),
            .I(N__31002));
    LocalMux I__2615 (
            .O(N__31002),
            .I(\pid_alt.O_4_6 ));
    InMux I__2614 (
            .O(N__30999),
            .I(N__30996));
    LocalMux I__2613 (
            .O(N__30996),
            .I(\pid_alt.O_4_5 ));
    InMux I__2612 (
            .O(N__30993),
            .I(N__30990));
    LocalMux I__2611 (
            .O(N__30990),
            .I(\pid_alt.O_4_8 ));
    InMux I__2610 (
            .O(N__30987),
            .I(N__30984));
    LocalMux I__2609 (
            .O(N__30984),
            .I(\pid_alt.O_4_7 ));
    InMux I__2608 (
            .O(N__30981),
            .I(N__30978));
    LocalMux I__2607 (
            .O(N__30978),
            .I(\pid_alt.O_4_10 ));
    InMux I__2606 (
            .O(N__30975),
            .I(N__30972));
    LocalMux I__2605 (
            .O(N__30972),
            .I(N__30969));
    Span4Mux_h I__2604 (
            .O(N__30969),
            .I(N__30966));
    Odrv4 I__2603 (
            .O(N__30966),
            .I(\pid_alt.O_4_4 ));
    InMux I__2602 (
            .O(N__30963),
            .I(N__30960));
    LocalMux I__2601 (
            .O(N__30960),
            .I(\pid_alt.O_4_21 ));
    InMux I__2600 (
            .O(N__30957),
            .I(N__30954));
    LocalMux I__2599 (
            .O(N__30954),
            .I(N__30951));
    Odrv4 I__2598 (
            .O(N__30951),
            .I(\pid_alt.O_4_13 ));
    InMux I__2597 (
            .O(N__30948),
            .I(N__30945));
    LocalMux I__2596 (
            .O(N__30945),
            .I(N__30942));
    Odrv4 I__2595 (
            .O(N__30942),
            .I(\pid_alt.O_4_16 ));
    InMux I__2594 (
            .O(N__30939),
            .I(N__30936));
    LocalMux I__2593 (
            .O(N__30936),
            .I(N__30933));
    Odrv4 I__2592 (
            .O(N__30933),
            .I(\pid_alt.O_4_22 ));
    InMux I__2591 (
            .O(N__30930),
            .I(N__30927));
    LocalMux I__2590 (
            .O(N__30927),
            .I(N__30924));
    Odrv4 I__2589 (
            .O(N__30924),
            .I(\pid_alt.O_4_17 ));
    InMux I__2588 (
            .O(N__30921),
            .I(N__30918));
    LocalMux I__2587 (
            .O(N__30918),
            .I(\pid_alt.O_4_14 ));
    InMux I__2586 (
            .O(N__30915),
            .I(N__30912));
    LocalMux I__2585 (
            .O(N__30912),
            .I(\pid_alt.O_4_9 ));
    InMux I__2584 (
            .O(N__30909),
            .I(N__30906));
    LocalMux I__2583 (
            .O(N__30906),
            .I(N__30903));
    Odrv4 I__2582 (
            .O(N__30903),
            .I(\pid_alt.O_4_23 ));
    InMux I__2581 (
            .O(N__30900),
            .I(N__30897));
    LocalMux I__2580 (
            .O(N__30897),
            .I(N__30894));
    Odrv4 I__2579 (
            .O(N__30894),
            .I(\pid_alt.O_4_19 ));
    InMux I__2578 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__2577 (
            .O(N__30888),
            .I(\pid_alt.O_4_12 ));
    InMux I__2576 (
            .O(N__30885),
            .I(N__30882));
    LocalMux I__2575 (
            .O(N__30882),
            .I(N__30879));
    Span4Mux_v I__2574 (
            .O(N__30879),
            .I(N__30876));
    Odrv4 I__2573 (
            .O(N__30876),
            .I(alt_ki_2));
    InMux I__2572 (
            .O(N__30873),
            .I(N__30870));
    LocalMux I__2571 (
            .O(N__30870),
            .I(N__30867));
    Odrv4 I__2570 (
            .O(N__30867),
            .I(alt_ki_3));
    InMux I__2569 (
            .O(N__30864),
            .I(N__30861));
    LocalMux I__2568 (
            .O(N__30861),
            .I(N__30858));
    Span4Mux_s2_h I__2567 (
            .O(N__30858),
            .I(N__30855));
    Odrv4 I__2566 (
            .O(N__30855),
            .I(alt_ki_4));
    InMux I__2565 (
            .O(N__30852),
            .I(N__30849));
    LocalMux I__2564 (
            .O(N__30849),
            .I(N__30846));
    Odrv4 I__2563 (
            .O(N__30846),
            .I(alt_ki_5));
    InMux I__2562 (
            .O(N__30843),
            .I(N__30840));
    LocalMux I__2561 (
            .O(N__30840),
            .I(N__30837));
    Span4Mux_s2_h I__2560 (
            .O(N__30837),
            .I(N__30834));
    Odrv4 I__2559 (
            .O(N__30834),
            .I(alt_ki_6));
    InMux I__2558 (
            .O(N__30831),
            .I(N__30828));
    LocalMux I__2557 (
            .O(N__30828),
            .I(N__30825));
    Span4Mux_v I__2556 (
            .O(N__30825),
            .I(N__30822));
    Odrv4 I__2555 (
            .O(N__30822),
            .I(alt_ki_7));
    InMux I__2554 (
            .O(N__30819),
            .I(N__30816));
    LocalMux I__2553 (
            .O(N__30816),
            .I(N__30813));
    Span4Mux_h I__2552 (
            .O(N__30813),
            .I(N__30810));
    Odrv4 I__2551 (
            .O(N__30810),
            .I(\pid_alt.O_4_24 ));
    InMux I__2550 (
            .O(N__30807),
            .I(N__30804));
    LocalMux I__2549 (
            .O(N__30804),
            .I(N__30801));
    Odrv4 I__2548 (
            .O(N__30801),
            .I(\pid_alt.O_4_11 ));
    InMux I__2547 (
            .O(N__30798),
            .I(N__30795));
    LocalMux I__2546 (
            .O(N__30795),
            .I(N__30792));
    Odrv4 I__2545 (
            .O(N__30792),
            .I(\pid_alt.O_4_18 ));
    InMux I__2544 (
            .O(N__30789),
            .I(N__30786));
    LocalMux I__2543 (
            .O(N__30786),
            .I(\pid_alt.O_3_6 ));
    InMux I__2542 (
            .O(N__30783),
            .I(N__30780));
    LocalMux I__2541 (
            .O(N__30780),
            .I(\pid_alt.O_3_7 ));
    InMux I__2540 (
            .O(N__30777),
            .I(N__30774));
    LocalMux I__2539 (
            .O(N__30774),
            .I(\pid_alt.O_3_8 ));
    InMux I__2538 (
            .O(N__30771),
            .I(N__30768));
    LocalMux I__2537 (
            .O(N__30768),
            .I(\pid_alt.O_3_16 ));
    InMux I__2536 (
            .O(N__30765),
            .I(N__30762));
    LocalMux I__2535 (
            .O(N__30762),
            .I(\pid_alt.O_3_20 ));
    InMux I__2534 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__2533 (
            .O(N__30756),
            .I(\pid_alt.O_3_9 ));
    InMux I__2532 (
            .O(N__30753),
            .I(N__30750));
    LocalMux I__2531 (
            .O(N__30750),
            .I(\pid_alt.O_3_13 ));
    InMux I__2530 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__2529 (
            .O(N__30744),
            .I(N__30741));
    Span4Mux_v I__2528 (
            .O(N__30741),
            .I(N__30738));
    Odrv4 I__2527 (
            .O(N__30738),
            .I(alt_ki_0));
    InMux I__2526 (
            .O(N__30735),
            .I(N__30732));
    LocalMux I__2525 (
            .O(N__30732),
            .I(N__30729));
    Span4Mux_v I__2524 (
            .O(N__30729),
            .I(N__30726));
    Odrv4 I__2523 (
            .O(N__30726),
            .I(alt_ki_1));
    InMux I__2522 (
            .O(N__30723),
            .I(N__30720));
    LocalMux I__2521 (
            .O(N__30720),
            .I(\pid_alt.O_3_15 ));
    InMux I__2520 (
            .O(N__30717),
            .I(N__30714));
    LocalMux I__2519 (
            .O(N__30714),
            .I(N__30711));
    Odrv4 I__2518 (
            .O(N__30711),
            .I(\pid_alt.O_3_19 ));
    InMux I__2517 (
            .O(N__30708),
            .I(N__30705));
    LocalMux I__2516 (
            .O(N__30705),
            .I(N__30702));
    Odrv4 I__2515 (
            .O(N__30702),
            .I(\pid_alt.O_3_17 ));
    InMux I__2514 (
            .O(N__30699),
            .I(N__30696));
    LocalMux I__2513 (
            .O(N__30696),
            .I(N__30693));
    Odrv4 I__2512 (
            .O(N__30693),
            .I(\pid_alt.O_3_18 ));
    InMux I__2511 (
            .O(N__30690),
            .I(N__30687));
    LocalMux I__2510 (
            .O(N__30687),
            .I(\pid_alt.O_3_10 ));
    InMux I__2509 (
            .O(N__30684),
            .I(N__30681));
    LocalMux I__2508 (
            .O(N__30681),
            .I(\pid_alt.O_3_14 ));
    InMux I__2507 (
            .O(N__30678),
            .I(N__30675));
    LocalMux I__2506 (
            .O(N__30675),
            .I(N__30672));
    Odrv4 I__2505 (
            .O(N__30672),
            .I(\pid_alt.O_3_24 ));
    InMux I__2504 (
            .O(N__30669),
            .I(N__30666));
    LocalMux I__2503 (
            .O(N__30666),
            .I(\pid_alt.O_3_22 ));
    InMux I__2502 (
            .O(N__30663),
            .I(N__30660));
    LocalMux I__2501 (
            .O(N__30660),
            .I(\pid_alt.O_3_23 ));
    InMux I__2500 (
            .O(N__30657),
            .I(N__30654));
    LocalMux I__2499 (
            .O(N__30654),
            .I(N__30651));
    Odrv4 I__2498 (
            .O(N__30651),
            .I(\pid_alt.O_3_12 ));
    InMux I__2497 (
            .O(N__30648),
            .I(N__30645));
    LocalMux I__2496 (
            .O(N__30645),
            .I(N__30642));
    Odrv4 I__2495 (
            .O(N__30642),
            .I(\pid_alt.O_3_21 ));
    InMux I__2494 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__2493 (
            .O(N__30636),
            .I(\pid_alt.O_3_11 ));
    IoInMux I__2492 (
            .O(N__30633),
            .I(N__30630));
    LocalMux I__2491 (
            .O(N__30630),
            .I(N__30627));
    Span4Mux_s0_v I__2490 (
            .O(N__30627),
            .I(N__30624));
    Sp12to4 I__2489 (
            .O(N__30624),
            .I(N__30621));
    Span12Mux_h I__2488 (
            .O(N__30621),
            .I(N__30618));
    Span12Mux_v I__2487 (
            .O(N__30618),
            .I(N__30615));
    Span12Mux_v I__2486 (
            .O(N__30615),
            .I(N__30612));
    Odrv12 I__2485 (
            .O(N__30612),
            .I(\Pc2drone_pll_inst.clk_system_pll ));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_21_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_8_0_));
    defparam IN_MUX_bfv_21_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_9_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_21_9_0_));
    defparam IN_MUX_bfv_21_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_21_10_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\pid_side.un11lto30_i_a2_6 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\pid_front.un11lto30_i_a2_6 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\pid_alt.error_i_acumm_prereg6_cry_7 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\pid_alt.error_i_acumm_prereg6 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_14_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_2_0_));
    defparam IN_MUX_bfv_14_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_3_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_14_3_0_));
    defparam IN_MUX_bfv_14_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_4_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_14_4_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\pid_side.error_cry_3_0 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(\pid_front.error_cry_3_0 ),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\pid_alt.un2_pid_prereg_cry_7 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pid_alt.un2_pid_prereg_cry_15 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_9_6_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__54900),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_side.state_RNIL5IF_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__62334),
            .GLOBALBUFFEROUTPUT(\pid_side.N_478_g ));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__36528),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_579_0_g ));
    ICE_GB \Pc2drone_pll_inst.PLLOUTCORE_derived_clock_RNI5FOA  (
            .USERSIGNALTOGLOBALBUFFER(N__30633),
            .GLOBALBUFFEROUTPUT(clk_system_pll_g));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__76710),
            .GLOBALBUFFEROUTPUT(N_580_g));
    ICE_GB \pid_side.state_RNIIIOO_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__63816),
            .GLOBALBUFFEROUTPUT(\pid_side.N_1352_g ));
    ICE_GB \pid_front.state_RNIPKTD_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__42198),
            .GLOBALBUFFEROUTPUT(\pid_front.N_404_g ));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__50007),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_8_LC_1_4_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_4_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_1_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30657),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83907),
            .ce(N__36268),
            .sr(N__82894));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30648),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83907),
            .ce(N__36268),
            .sr(N__82894));
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30639),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_11_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30723),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30717),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30708),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30699),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_5_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30690),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30684),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83918),
            .ce(N__36270),
            .sr(N__82893));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30678),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30669),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30663),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_6_3  (
            .in0(N__30789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_6_4  (
            .in0(N__30783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__30777),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30771),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30765),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83931),
            .ce(N__36271),
            .sr(N__82892));
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30759),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83943),
            .ce(N__36272),
            .sr(N__82891));
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30753),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83943),
            .ce(N__36272),
            .sr(N__82891));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_8_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_1_8_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__80515),
            .in2(_gnd_net_),
            .in3(N__83029),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_1_8_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_1_8_1  (
            .in0(N__83030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73740),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_1_8_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_1_8_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__80248),
            .in2(_gnd_net_),
            .in3(N__83031),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_8_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_1_8_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_1_8_3  (
            .in0(N__83032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79720),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_1_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__79276),
            .in2(_gnd_net_),
            .in3(N__83033),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_8_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_1_8_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_1_8_5  (
            .in0(N__83034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80108),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_1_8_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__81076),
            .in2(_gnd_net_),
            .in3(N__83035),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_1_8_7  (
            .in0(N__83036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79890),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83958),
            .ce(N__38325),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30819),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83972),
            .ce(N__36273),
            .sr(N__82890));
    defparam \pid_alt.error_i_reg_esr_7_LC_1_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30807),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83972),
            .ce(N__36273),
            .sr(N__82890));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30798),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83972),
            .ce(N__36273),
            .sr(N__82890));
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30957),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83972),
            .ce(N__36273),
            .sr(N__82890));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30948),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30939),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30930),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30921),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_10_4  (
            .in0(N__30915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30909),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30900),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83988),
            .ce(N__36274),
            .sr(N__82888));
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30891),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31017),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31011),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31005),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_1_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30999),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__30993),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30987),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30981),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84006),
            .ce(N__36275),
            .sr(N__82887));
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30975),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84023),
            .ce(N__36276),
            .sr(N__82886));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30963),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84023),
            .ce(N__36276),
            .sr(N__82886));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9ABT5_5_LC_1_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9ABT5_5_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9ABT5_5_LC_1_13_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9ABT5_5_LC_1_13_0  (
            .in0(N__31074),
            .in1(N__34896),
            .in2(N__31065),
            .in3(N__33088),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9ABT5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_1_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_1_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_1_13_1  (
            .in0(N__33011),
            .in1(N__32987),
            .in2(_gnd_net_),
            .in3(N__33038),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9AMU2_5_LC_1_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9AMU2_5_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9AMU2_5_LC_1_13_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9AMU2_5_LC_1_13_2  (
            .in0(N__31064),
            .in1(_gnd_net_),
            .in2(N__31068),
            .in3(N__33089),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9AMU2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31053),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84038),
            .ce(N__37530),
            .sr(N__77300));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_1_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_1_13_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_1_13_5  (
            .in0(N__32036),
            .in1(N__31031),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_13_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_1_13_6  (
            .in0(N__31052),
            .in1(_gnd_net_),
            .in2(N__31035),
            .in3(N__32037),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUDT5_6_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUDT5_6_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUDT5_6_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIRUDT5_6_LC_1_13_7  (
            .in0(N__35111),
            .in1(N__35331),
            .in2(N__31023),
            .in3(N__33916),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIRUDT5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_1_14_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_1_14_1  (
            .in0(N__32648),
            .in1(N__32559),
            .in2(_gnd_net_),
            .in3(N__32589),
            .lcout(\pid_alt.un1_pid_prereg_236_1 ),
            .ltout(\pid_alt.un1_pid_prereg_236_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISEDF3_19_LC_1_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISEDF3_19_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISEDF3_19_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISEDF3_19_LC_1_14_2  (
            .in0(N__35199),
            .in1(N__31142),
            .in2(N__31020),
            .in3(N__32860),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISEDF3Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_1_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_1_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32590),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84053),
            .ce(N__37527),
            .sr(N__77310));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGRON1_19_LC_1_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGRON1_19_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGRON1_19_LC_1_14_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGRON1_19_LC_1_14_4  (
            .in0(N__31149),
            .in1(N__31143),
            .in2(_gnd_net_),
            .in3(N__32861),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGRON1Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_1_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_1_14_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_1_14_5  (
            .in0(N__31869),
            .in1(N__31134),
            .in2(_gnd_net_),
            .in3(N__31124),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_1_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_1_14_6  (
            .in0(N__31125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84053),
            .ce(N__37527),
            .sr(N__77310));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_14_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_14_7  (
            .in0(N__31868),
            .in1(N__31133),
            .in2(_gnd_net_),
            .in3(N__31123),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_20_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31110),
            .lcout(\pid_front.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_21_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31101),
            .lcout(\pid_front.error_p_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_9_LC_1_15_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_9_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_9_LC_1_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_9_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31092),
            .lcout(\pid_front.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_4_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31086),
            .lcout(\pid_front.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_5_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31080),
            .lcout(\pid_front.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_2_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31203),
            .lcout(\pid_front.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_7_LC_1_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_7_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_7_LC_1_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_7_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31197),
            .lcout(\pid_front.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_8_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31191),
            .lcout(\pid_front.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84072),
            .ce(N__83133),
            .sr(N__82885));
    defparam \pid_front.error_p_reg_esr_13_LC_1_16_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_13_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_13_LC_1_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_13_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31185),
            .lcout(\pid_front.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_14_LC_1_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_14_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_14_LC_1_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_14_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31179),
            .lcout(\pid_front.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_15_LC_1_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_15_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_15_LC_1_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_15_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31173),
            .lcout(\pid_front.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_16_LC_1_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_16_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31167),
            .lcout(\pid_front.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_17_LC_1_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_17_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31161),
            .lcout(\pid_front.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_18_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_18_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_18_LC_1_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_18_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31155),
            .lcout(\pid_front.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_19_LC_1_16_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_19_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_19_LC_1_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_19_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31461),
            .lcout(\pid_front.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_6_LC_1_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_6_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31455),
            .lcout(\pid_front.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84084),
            .ce(N__83131),
            .sr(N__82884));
    defparam \pid_alt.error_cry_0_c_LC_1_17_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_1_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__32762),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNIO4P5_LC_1_17_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNIO4P5_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNIO4P5_LC_1_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNIO4P5_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__36441),
            .in2(_gnd_net_),
            .in3(N__31413),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNIQ7Q5_LC_1_17_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNIQ7Q5_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNIQ7Q5_LC_1_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNIQ7Q5_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__32739),
            .in2(_gnd_net_),
            .in3(N__31371),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNISAR5_LC_1_17_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNISAR5_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNISAR5_LC_1_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_2_c_RNISAR5_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32784),
            .in3(N__31332),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKI0D_LC_1_17_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKI0D_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKI0D_LC_1_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKI0D_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__32775),
            .in2(N__34119),
            .in3(N__31287),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINM1D_LC_1_17_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINM1D_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINM1D_LC_1_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINM1D_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__31809),
            .in2(N__34089),
            .in3(N__31245),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQQ2D_LC_1_17_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQQ2D_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQQ2D_LC_1_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQQ2D_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__31800),
            .in2(N__34011),
            .in3(N__31206),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITU3D_LC_1_17_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITU3D_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITU3D_LC_1_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITU3D_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__52743),
            .in2(N__34548),
            .in3(N__31737),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI035D_LC_1_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI035D_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI035D_LC_1_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI035D_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__34494),
            .in2(N__32751),
            .in3(N__31695),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNI376D_LC_1_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNI376D_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNI376D_LC_1_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNI376D_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__36402),
            .in2(N__34464),
            .in3(N__31656),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIDR2H_LC_1_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIDR2H_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIDR2H_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIDR2H_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__32733),
            .in2(N__34416),
            .in3(N__31617),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNIN0IL_LC_1_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNIN0IL_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNIN0IL_LC_1_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNIN0IL_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__32724),
            .in2(N__34370),
            .in3(N__31578),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNISNEE_LC_1_18_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNISNEE_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNISNEE_LC_1_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_11_c_RNISNEE_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__32769),
            .in2(_gnd_net_),
            .in3(N__31539),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNIUQFE_LC_1_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNIUQFE_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNIUQFE_LC_1_18_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_12_c_RNIUQFE_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31818),
            .in3(N__31503),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI0UGE_LC_1_18_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI0UGE_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI0UGE_LC_1_18_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_13_c_RNI0UGE_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31791),
            .in3(N__31464),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNI21IE_LC_1_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNI21IE_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNI21IE_LC_1_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNI21IE_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__52881),
            .in2(_gnd_net_),
            .in3(N__31857),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_13_LC_1_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_13_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_13_LC_1_19_0 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_13_LC_1_19_0  (
            .in0(N__34316),
            .in1(N__52850),
            .in2(N__58510),
            .in3(N__68636),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84102),
            .ce(),
            .sr(N__77343));
    defparam \pid_alt.error_axb_13_LC_1_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_1_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34315),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_5_LC_1_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_5_LC_1_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_5_LC_1_19_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_5_LC_1_19_2  (
            .in0(N__34055),
            .in1(N__52852),
            .in2(N__58512),
            .in3(N__68637),
            .lcout(drone_altitude_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84102),
            .ce(),
            .sr(N__77343));
    defparam \dron_frame_decoder_1.source_Altitude_RNI9143_5_LC_1_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNI9143_5_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNI9143_5_LC_1_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNI9143_5_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34054),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_14_LC_1_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_14_LC_1_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_14_LC_1_19_4 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_14_LC_1_19_4  (
            .in0(N__34295),
            .in1(N__52851),
            .in2(N__58511),
            .in3(N__68573),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84102),
            .ce(),
            .sr(N__77343));
    defparam \dron_frame_decoder_1.source_Altitude_6_LC_1_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_6_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_6_LC_1_19_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_6_LC_1_19_5  (
            .in0(N__52853),
            .in1(N__34031),
            .in2(N__68574),
            .in3(N__58495),
            .lcout(drone_altitude_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84102),
            .ce(),
            .sr(N__77343));
    defparam \dron_frame_decoder_1.source_Altitude_RNIA243_6_LC_1_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNIA243_6_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNIA243_6_LC_1_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNIA243_6_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34027),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_14_LC_1_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_1_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34294),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31782),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31962),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31950),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31938),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31926),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31917),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31905),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84109),
            .ce(N__36281),
            .sr(N__82881));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31896),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31887),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31878),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32064),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32055),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_23_6  (
            .in0(N__32049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32043),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84112),
            .ce(N__36282),
            .sr(N__82878));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_5_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_5_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_2_5_1  (
            .in0(N__83040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73728),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83909),
            .ce(N__38310),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_5_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_5_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__80275),
            .in2(_gnd_net_),
            .in3(N__83041),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83909),
            .ce(N__38310),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_5_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_5_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__80500),
            .in2(_gnd_net_),
            .in3(N__83039),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83909),
            .ce(N__38310),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_5_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_5_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_2_5_5  (
            .in0(N__83042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80100),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83909),
            .ce(N__38310),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_5_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_5_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_2_5_7  (
            .in0(N__83043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79909),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83909),
            .ce(N__38310),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_6_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__79258),
            .in2(_gnd_net_),
            .in3(N__83037),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83920),
            .ce(N__38308),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__81080),
            .in2(_gnd_net_),
            .in3(N__83038),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83920),
            .ce(N__38308),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__79697),
            .in2(_gnd_net_),
            .in3(N__83028),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83933),
            .ce(N__38309),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_2_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_2_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37660),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83945),
            .ce(N__37533),
            .sr(N__77256));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_8_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33034),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83945),
            .ce(N__37533),
            .sr(N__77256));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32694),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83960),
            .ce(N__34658),
            .sr(N__77263));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_2_9_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36034),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83960),
            .ce(N__34658),
            .sr(N__77263));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_2_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37759),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83960),
            .ce(N__34658),
            .sr(N__77263));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_2_9_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33339),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83960),
            .ce(N__34658),
            .sr(N__77263));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_2_9_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_2_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33930),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83960),
            .ce(N__34658),
            .sr(N__77263));
    defparam \pid_alt.error_i_acumm_10_LC_2_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_2_10_0 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_2_10_0  (
            .in0(N__36984),
            .in1(N__47726),
            .in2(N__32244),
            .in3(N__33054),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_11_LC_2_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_2_10_1 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_2_10_1  (
            .in0(N__47723),
            .in1(N__33153),
            .in2(N__32210),
            .in3(N__36985),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_6_LC_2_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_2_10_2 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_2_10_2  (
            .in0(N__36986),
            .in1(N__32375),
            .in2(N__33075),
            .in3(N__47730),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_7_LC_2_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_2_10_3 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_2_10_3  (
            .in0(N__47724),
            .in1(N__34841),
            .in2(N__32349),
            .in3(N__36987),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_8_LC_2_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_2_10_4 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_2_10_4  (
            .in0(N__36988),
            .in1(N__33173),
            .in2(N__32313),
            .in3(N__47731),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_9_LC_2_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_2_10_5 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_2_10_5  (
            .in0(N__47725),
            .in1(N__33189),
            .in2(N__32280),
            .in3(N__36989),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_10_6  (
            .in0(N__33070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34840),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_12_LC_2_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_2_10_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_2_10_7  (
            .in0(N__34818),
            .in1(N__32525),
            .in2(N__47733),
            .in3(N__33207),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83976),
            .ce(),
            .sr(N__46503));
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_2_11_0 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_2_11_0  (
            .in0(N__32159),
            .in1(N__37029),
            .in2(N__33138),
            .in3(N__46626),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83992),
            .ce(N__36935),
            .sr(N__46507));
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_2_11_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_2_11_1  (
            .in0(N__46627),
            .in1(N__33117),
            .in2(N__37037),
            .in3(N__32160),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83992),
            .ce(N__36935),
            .sr(N__46507));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_2_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_2_11_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_2_11_2  (
            .in0(N__36982),
            .in1(N__32172),
            .in2(N__32916),
            .in3(N__34817),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(\pid_alt.N_62_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_2_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_2_11_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__46576),
            .in2(N__32166),
            .in3(N__36983),
            .lcout(\pid_alt.N_94 ),
            .ltout(\pid_alt.N_94_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_2_11_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_2_11_4  (
            .in0(N__34857),
            .in1(N__37028),
            .in2(N__32163),
            .in3(N__46625),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83992),
            .ce(N__36935),
            .sr(N__46507));
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_2_11_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_2_11_5  (
            .in0(N__46624),
            .in1(N__34872),
            .in2(N__37036),
            .in3(N__32158),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83992),
            .ce(N__36935),
            .sr(N__46507));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_12_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_12_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__32933),
            .in2(N__32954),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pid_alt.un2_pid_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_0_c_RNIEO2R_LC_2_12_1 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_0_c_RNIEO2R_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_0_c_RNIEO2R_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_0_c_RNIEO2R_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__32148),
            .in2(N__32142),
            .in3(N__32133),
            .lcout(\pid_alt.un2_pid_prereg_cry_0_c_RNIEO2R ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_0 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_1_c_RNIHS3R_LC_2_12_2 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_1_c_RNIHS3R_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_1_c_RNIHS3R_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_1_c_RNIHS3R_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__32130),
            .in2(N__32124),
            .in3(N__32115),
            .lcout(\pid_alt.un2_pid_prereg_cry_1_c_RNIHS3R ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_1 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_2_c_RNIK05R_LC_2_12_3 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_2_c_RNIK05R_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_2_c_RNIK05R_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_2_c_RNIK05R_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__32112),
            .in2(N__32106),
            .in3(N__32097),
            .lcout(\pid_alt.un2_pid_prereg_cry_2_c_RNIK05R ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_2 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_3_c_RNIN46R_LC_2_12_4 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_3_c_RNIN46R_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_3_c_RNIN46R_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_3_c_RNIN46R_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__36948),
            .in2(N__32403),
            .in3(N__32394),
            .lcout(\pid_alt.un2_pid_prereg_cry_3_c_RNIN46R ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_3 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_4_c_RNIHA9S_LC_2_12_5 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_4_c_RNIHA9S_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_4_c_RNIHA9S_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_4_c_RNIHA9S_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__46545),
            .in2(N__32391),
            .in3(N__32379),
            .lcout(\pid_alt.un2_pid_prereg_cry_4_c_RNIHA9S ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_4 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_5_c_RNIKEAS_LC_2_12_6 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_5_c_RNIKEAS_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_5_c_RNIKEAS_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_5_c_RNIKEAS_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__32376),
            .in2(N__32361),
            .in3(N__32352),
            .lcout(\pid_alt.un2_pid_prereg_cry_5_c_RNIKEAS ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_5 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_6_c_RNINIBS_LC_2_12_7 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_6_c_RNINIBS_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_6_c_RNINIBS_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_6_c_RNINIBS_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__32348),
            .in2(N__32331),
            .in3(N__32316),
            .lcout(\pid_alt.un2_pid_prereg_cry_6_c_RNINIBS ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_6 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_7_c_RNIQMCS_LC_2_13_0 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_7_c_RNIQMCS_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_7_c_RNIQMCS_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_7_c_RNIQMCS_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__32309),
            .in2(N__32295),
            .in3(N__32283),
            .lcout(\pid_alt.un2_pid_prereg_cry_7_c_RNIQMCS ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pid_alt.un2_pid_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_8_c_RNITQDS_LC_2_13_1 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_8_c_RNITQDS_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_8_c_RNITQDS_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_8_c_RNITQDS_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__32279),
            .in2(N__32262),
            .in3(N__32247),
            .lcout(\pid_alt.un2_pid_prereg_cry_8_c_RNITQDS ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_8 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_9_c_RNIEPOG_LC_2_13_2 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_9_c_RNIEPOG_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_9_c_RNIEPOG_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_9_c_RNIEPOG_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__32243),
            .in2(N__32226),
            .in3(N__32214),
            .lcout(\pid_alt.un2_pid_prereg_cry_9_c_RNIEPOG ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_9 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_10_c_RNIOCDG_LC_2_13_3 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_10_c_RNIOCDG_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_10_c_RNIOCDG_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_10_c_RNIOCDG_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__32211),
            .in2(N__32190),
            .in3(N__32175),
            .lcout(\pid_alt.un2_pid_prereg_cry_10_c_RNIOCDG ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_10 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_11_c_RNIRGEG_LC_2_13_4 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_11_c_RNIRGEG_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_11_c_RNIRGEG_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_11_c_RNIRGEG_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__32541),
            .in2(N__32529),
            .in3(N__32511),
            .lcout(\pid_alt.un2_pid_prereg_cry_11_c_RNIRGEG ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_11 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_12_c_RNI7SBD_LC_2_13_5 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_12_c_RNI7SBD_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_12_c_RNI7SBD_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_12_c_RNI7SBD_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__34704),
            .in2(N__32508),
            .in3(N__32496),
            .lcout(\pid_alt.un2_pid_prereg_cry_12_c_RNI7SBD ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_12 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_13_c_RNILQAA_LC_2_13_6 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_13_c_RNILQAA_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_13_c_RNILQAA_LC_2_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_13_c_RNILQAA_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__32493),
            .in2(_gnd_net_),
            .in3(N__32481),
            .lcout(\pid_alt.un2_pid_prereg_cry_13_c_RNILQAA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_13 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_14_c_RNINTBA_LC_2_13_7 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_14_c_RNINTBA_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_14_c_RNINTBA_LC_2_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_14_c_RNINTBA_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__32478),
            .in2(_gnd_net_),
            .in3(N__32466),
            .lcout(\pid_alt.un2_pid_prereg_cry_14_c_RNINTBA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_14 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_15_c_RNIP0DA_LC_2_14_0 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_15_c_RNIP0DA_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_15_c_RNIP0DA_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_15_c_RNIP0DA_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__32463),
            .in2(_gnd_net_),
            .in3(N__32451),
            .lcout(\pid_alt.un2_pid_prereg_cry_15_c_RNIP0DA ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pid_alt.un2_pid_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_16_c_RNIR3EA_LC_2_14_1 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_16_c_RNIR3EA_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_16_c_RNIR3EA_LC_2_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_16_c_RNIR3EA_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__32448),
            .in2(_gnd_net_),
            .in3(N__32439),
            .lcout(\pid_alt.un2_pid_prereg_cry_16_c_RNIR3EA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_16 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_17_c_RNIT6FA_LC_2_14_2 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_17_c_RNIT6FA_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_17_c_RNIT6FA_LC_2_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_17_c_RNIT6FA_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__32436),
            .in2(_gnd_net_),
            .in3(N__32424),
            .lcout(\pid_alt.un2_pid_prereg_cry_17_c_RNIT6FA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_17 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_18_c_RNIV9GA_LC_2_14_3 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_18_c_RNIV9GA_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_18_c_RNIV9GA_LC_2_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_18_c_RNIV9GA_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__32421),
            .in2(_gnd_net_),
            .in3(N__32409),
            .lcout(\pid_alt.un2_pid_prereg_cry_18_c_RNIV9GA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_18 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_19_c_RNIO4IA_LC_2_14_4 .C_ON=1'b1;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_19_c_RNIO4IA_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_19_c_RNIO4IA_LC_2_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_19_c_RNIO4IA_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__32717),
            .in2(_gnd_net_),
            .in3(N__32406),
            .lcout(\pid_alt.un2_pid_prereg_cry_19_c_RNIO4IA ),
            .ltout(),
            .carryin(\pid_alt.un2_pid_prereg_cry_19 ),
            .carryout(\pid_alt.un2_pid_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_20_c_RNIGLBB_LC_2_14_5 .C_ON=1'b0;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_20_c_RNIGLBB_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_20_c_RNIGLBB_LC_2_14_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un2_pid_prereg_un2_pid_prereg_cry_20_c_RNIGLBB_LC_2_14_5  (
            .in0(N__32718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32703),
            .lcout(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB ),
            .ltout(\pid_alt.un2_pid_prereg_cry_20_c_RNIGLBB_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_20_LC_2_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_20_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_20_LC_2_14_6 .LUT_INIT=16'b1111010011010000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI06021_20_LC_2_14_6  (
            .in0(N__32567),
            .in1(N__32663),
            .in2(N__32700),
            .in3(N__32602),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI06021Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_2_20_LC_2_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_2_20_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_2_20_LC_2_14_7 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI06021_2_20_LC_2_14_7  (
            .in0(N__32603),
            .in1(N__32568),
            .in2(N__32667),
            .in3(N__32690),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI06021_2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_1_20_LC_2_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_1_20_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_1_20_LC_2_15_0 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI06021_1_20_LC_2_15_0  (
            .in0(N__32570),
            .in1(N__32612),
            .in2(N__32662),
            .in3(N__32688),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI06021_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_0_20_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_0_20_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI06021_0_20_LC_2_15_2 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI06021_0_20_LC_2_15_2  (
            .in0(N__32569),
            .in1(N__32611),
            .in2(N__32661),
            .in3(N__32687),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI06021_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_2_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_2_15_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_2_15_5  (
            .in0(N__37716),
            .in1(N__37688),
            .in2(_gnd_net_),
            .in3(N__37668),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI060F3_15_LC_2_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI060F3_15_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI060F3_15_LC_2_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI060F3_15_LC_2_15_6  (
            .in0(N__33600),
            .in1(N__37736),
            .in2(N__32697),
            .in3(N__33958),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI060F3Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_15_7 .LUT_INIT=16'b1111111001111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_15_7  (
            .in0(N__32689),
            .in1(N__32655),
            .in2(N__32616),
            .in3(N__32571),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_0_LC_2_16_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_0_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_0_LC_2_16_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_0_LC_2_16_0  (
            .in0(N__34199),
            .in1(N__52854),
            .in2(N__58504),
            .in3(N__72042),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84076),
            .ce(),
            .sr(N__77317));
    defparam \pid_alt.error_cry_0_c_inv_LC_2_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_2_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_2_16_1  (
            .in0(N__32763),
            .in1(N__60630),
            .in2(_gnd_net_),
            .in3(N__34198),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_8_LC_2_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_8_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_8_LC_2_16_2 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_8_LC_2_16_2  (
            .in0(N__34508),
            .in1(N__52857),
            .in2(N__58506),
            .in3(N__72043),
            .lcout(drone_altitude_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84076),
            .ce(),
            .sr(N__77317));
    defparam \dron_frame_decoder_1.source_Altitude_RNIC443_8_LC_2_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNIC443_8_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNIC443_8_LC_2_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNIC443_8_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34507),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_10_LC_2_16_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_10_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_10_LC_2_16_4 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_10_LC_2_16_4  (
            .in0(N__34430),
            .in1(N__52855),
            .in2(N__58505),
            .in3(N__71833),
            .lcout(drone_altitude_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84076),
            .ce(),
            .sr(N__77317));
    defparam \dron_frame_decoder_1.source_Altitude_2_LC_2_16_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_2_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_2_LC_2_16_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_2_LC_2_16_5  (
            .in0(N__52856),
            .in1(N__34170),
            .in2(N__71842),
            .in3(N__58470),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84076),
            .ce(),
            .sr(N__77317));
    defparam \pid_alt.error_axb_2_LC_2_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_2_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34168),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_RNILMV6_10_LC_2_16_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNILMV6_10_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNILMV6_10_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNILMV6_10_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34429),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_11_LC_2_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_11_LC_2_17_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_11_LC_2_17_0 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_11_LC_2_17_0  (
            .in0(N__34385),
            .in1(N__52803),
            .in2(N__58507),
            .in3(N__64997),
            .lcout(drone_altitude_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84087),
            .ce(),
            .sr(N__77324));
    defparam \dron_frame_decoder_1.source_Altitude_RNIMNV6_11_LC_2_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNIMNV6_11_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNIMNV6_11_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNIMNV6_11_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34384),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_3_LC_2_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_3_LC_2_17_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_3_LC_2_17_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_3_LC_2_17_2  (
            .in0(N__34148),
            .in1(N__52805),
            .in2(N__58509),
            .in3(N__64998),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84087),
            .ce(),
            .sr(N__77324));
    defparam \pid_alt.error_axb_3_LC_2_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_2_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34147),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_12_LC_2_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_12_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_12_LC_2_17_4 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_12_LC_2_17_4  (
            .in0(N__34337),
            .in1(N__52804),
            .in2(N__58508),
            .in3(N__65209),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84087),
            .ce(),
            .sr(N__77324));
    defparam \dron_frame_decoder_1.source_Altitude_4_LC_2_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_4_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_4_LC_2_17_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_4_LC_2_17_5  (
            .in0(N__34133),
            .in1(N__58483),
            .in2(N__52824),
            .in3(N__65210),
            .lcout(drone_altitude_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84087),
            .ce(),
            .sr(N__77324));
    defparam \dron_frame_decoder_1.source_Altitude_RNI8043_4_LC_2_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNI8043_4_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNI8043_4_LC_2_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNI8043_4_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34132),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_2_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_2_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34336),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg15lto3_LC_2_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg15lto3_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg15lto3_LC_2_18_0 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \pid_alt.error_i_acumm_prereg15lto3_LC_2_18_0  (
            .in0(N__34004),
            .in1(N__34087),
            .in2(N__34547),
            .in3(N__34118),
            .lcout(\pid_alt.error_i_acumm_prereg15lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_0_LC_2_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_0_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_0_LC_2_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_0_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80517),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \Commands_frame_decoder.source_CH1data_esr_1_LC_2_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_1_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_1_LC_2_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_1_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73739),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \Commands_frame_decoder.source_CH1data_esr_2_LC_2_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_2_LC_2_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_2_LC_2_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_2_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80297),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \Commands_frame_decoder.source_CH1data_esr_3_LC_2_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_3_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_3_LC_2_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_3_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79715),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \pid_alt.error_i_acumm_prereg15lto7_2_LC_2_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg15lto7_2_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg15lto7_2_LC_2_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg15lto7_2_LC_2_18_5  (
            .in0(N__34415),
            .in1(N__34463),
            .in2(N__34371),
            .in3(N__34493),
            .lcout(\pid_alt.error_i_acumm_prereg15lto7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_18_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79288),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80088),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84094),
            .ce(N__37410),
            .sr(N__77331));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81101),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84101),
            .ce(N__37409),
            .sr(N__77340));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_19_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79930),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84101),
            .ce(N__37409),
            .sr(N__77340));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_21_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_21_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_21_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__81085),
            .in2(_gnd_net_),
            .in3(N__83026),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84104),
            .ce(N__38763),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(N__80296),
            .in2(_gnd_net_),
            .in3(N__83025),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84107),
            .ce(N__38773),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_23_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_23_4  (
            .in0(N__83024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79932),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84111),
            .ce(N__38774),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(N__73788),
            .in2(_gnd_net_),
            .in3(N__83023),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84111),
            .ce(N__38774),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__79730),
            .in2(_gnd_net_),
            .in3(N__83015),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84114),
            .ce(N__38775),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_3_8_0  (
            .in0(N__32874),
            .in1(N__32880),
            .in2(N__32847),
            .in3(N__32886),
            .lcout(),
            .ltout(\pid_alt.m7_e_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_8_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_8_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_3_8_1  (
            .in0(N__32922),
            .in1(N__32898),
            .in2(N__32892),
            .in3(N__32838),
            .lcout(\pid_alt.N_222 ),
            .ltout(\pid_alt.N_222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_8_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_8_2 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_3_8_2  (
            .in0(N__33206),
            .in1(N__34759),
            .in2(N__32889),
            .in3(N__34740),
            .lcout(\pid_alt.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_3_8_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_3_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_3_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33966),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83934),
            .ce(N__34662),
            .sr(N__77251));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_8_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_3_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33501),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83934),
            .ce(N__34662),
            .sr(N__77251));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_8_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_8_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_3_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33855),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83934),
            .ce(N__34662),
            .sr(N__77251));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_8_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_3_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_3_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32868),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83934),
            .ce(N__34662),
            .sr(N__77251));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_3_8_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_3_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_3_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37458),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83934),
            .ce(N__34662),
            .sr(N__77251));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_3_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_3_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_3_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__32958),
            .in2(_gnd_net_),
            .in3(N__32937),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_9_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_3_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35536),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_3_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33372),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_9_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_3_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33402),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_9_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33228),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_9_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33258),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_9_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_3_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33696),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_9_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36127),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83946),
            .ce(N__34657),
            .sr(N__77257));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_3_10_0  (
            .in0(N__33188),
            .in1(N__33152),
            .in2(N__33174),
            .in3(N__33053),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_3_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35866),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83961),
            .ce(N__34647),
            .sr(N__77264));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__33052),
            .in2(_gnd_net_),
            .in3(N__33205),
            .lcout(\pid_alt.m21_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_3_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33778),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83961),
            .ce(N__34647),
            .sr(N__77264));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_3_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_3_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_3_10_4  (
            .in0(N__33187),
            .in1(N__33169),
            .in2(N__33074),
            .in3(N__33151),
            .lcout(),
            .ltout(\pid_alt.m21_e_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_10_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_3_10_5  (
            .in0(N__33128),
            .in1(N__33113),
            .in2(N__33102),
            .in3(N__33099),
            .lcout(\pid_alt.m21_e_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33093),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83961),
            .ce(N__34647),
            .sr(N__77264));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33531),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83961),
            .ce(N__34647),
            .sr(N__77264));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0K6S5_4_LC_3_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0K6S5_4_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0K6S5_4_LC_3_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0K6S5_4_LC_3_11_0  (
            .in0(N__32964),
            .in1(N__33320),
            .in2(N__34929),
            .in3(N__33334),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0K6S5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_11_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_3_11_1  (
            .in0(N__33039),
            .in1(N__33012),
            .in2(_gnd_net_),
            .in3(N__32988),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI00LU2_4_LC_3_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI00LU2_4_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI00LU2_4_LC_3_11_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI00LU2_4_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__33321),
            .in2(N__33342),
            .in3(N__33335),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI00LU2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_11_3 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_3_11_3  (
            .in0(N__33280),
            .in1(N__33302),
            .in2(_gnd_net_),
            .in3(N__33311),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_3_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33282),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83977),
            .ce(N__37531),
            .sr(N__77271));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0KHT2_3_LC_3_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0KHT2_3_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0KHT2_3_LC_3_11_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0KHT2_3_LC_3_11_5  (
            .in0(N__35925),
            .in1(N__33264),
            .in2(_gnd_net_),
            .in3(N__33254),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0KHT2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_11_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_3_11_6  (
            .in0(N__33312),
            .in1(N__33303),
            .in2(_gnd_net_),
            .in3(N__33281),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2IS8_3_LC_3_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2IS8_3_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2IS8_3_LC_3_11_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL2IS8_3_LC_3_11_7  (
            .in0(N__35924),
            .in1(N__33253),
            .in2(N__33240),
            .in3(N__35982),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL2IS8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIEF0O3_12_LC_3_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIEF0O3_12_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIEF0O3_12_LC_3_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIEF0O3_12_LC_3_12_0  (
            .in0(N__33470),
            .in1(N__33237),
            .in2(N__34986),
            .in3(N__33220),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIEF0O3Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_12_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_3_12_1  (
            .in0(N__33419),
            .in1(N__33440),
            .in2(_gnd_net_),
            .in3(N__33460),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG0FQ1_12_LC_3_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG0FQ1_12_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG0FQ1_12_LC_3_12_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG0FQ1_12_LC_3_12_2  (
            .in0(N__33471),
            .in1(_gnd_net_),
            .in2(N__33231),
            .in3(N__33221),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG0FQ1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_12_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_3_12_3  (
            .in0(N__35742),
            .in1(N__35688),
            .in2(_gnd_net_),
            .in3(N__35708),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_3_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_3_12_4  (
            .in0(N__33462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83993),
            .ce(N__37528),
            .sr(N__77276));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUEHT1_11_LC_3_12_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUEHT1_11_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUEHT1_11_LC_3_12_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUEHT1_11_LC_3_12_5  (
            .in0(N__33654),
            .in1(N__33411),
            .in2(_gnd_net_),
            .in3(N__33395),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUEHT1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_12_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_3_12_6  (
            .in0(N__33461),
            .in1(_gnd_net_),
            .in2(N__33444),
            .in3(N__33420),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJJ1R3_11_LC_3_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJJ1R3_11_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJJ1R3_11_LC_3_12_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJJ1R3_11_LC_3_12_7  (
            .in0(N__33653),
            .in1(N__35016),
            .in2(N__33405),
            .in3(N__33394),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJJ1R3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5H064_10_LC_3_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5H064_10_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5H064_10_LC_3_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5H064_10_LC_3_13_0  (
            .in0(N__33350),
            .in1(N__33381),
            .in2(N__35037),
            .in3(N__33364),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5H064Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_3_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_3_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_3_13_1  (
            .in0(N__33572),
            .in1(N__33548),
            .in2(_gnd_net_),
            .in3(N__33592),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL4GT1_10_LC_3_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL4GT1_10_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL4GT1_10_LC_3_13_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL4GT1_10_LC_3_13_2  (
            .in0(N__33351),
            .in1(_gnd_net_),
            .in2(N__33375),
            .in3(N__33365),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL4GT1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_3_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_3_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_3_13_3  (
            .in0(N__33635),
            .in1(N__33671),
            .in2(_gnd_net_),
            .in3(N__33615),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_3_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_3_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_3_13_4  (
            .in0(N__33594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84012),
            .ce(N__37525),
            .sr(N__77281));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGCG82_9_LC_3_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGCG82_9_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGCG82_9_LC_3_13_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGCG82_9_LC_3_13_5  (
            .in0(N__33540),
            .in1(N__35754),
            .in2(_gnd_net_),
            .in3(N__33524),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGCG82Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_3_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_3_13_6 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_3_13_6  (
            .in0(N__33593),
            .in1(N__33573),
            .in2(N__33552),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKLA75_9_LC_3_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKLA75_9_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKLA75_9_LC_3_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKLA75_9_LC_3_13_7  (
            .in0(N__35066),
            .in1(N__35753),
            .in2(N__33534),
            .in3(N__33523),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKLA75Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0B5F3_17_LC_3_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0B5F3_17_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0B5F3_17_LC_3_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0B5F3_17_LC_3_14_0  (
            .in0(N__33479),
            .in1(N__33510),
            .in2(N__35262),
            .in3(N__33493),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0B5F3Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_3_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_3_14_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_3_14_1  (
            .in0(N__33746),
            .in1(N__33755),
            .in2(_gnd_net_),
            .in3(N__33724),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI4AJN1_17_LC_3_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI4AJN1_17_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI4AJN1_17_LC_3_14_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI4AJN1_17_LC_3_14_2  (
            .in0(N__33480),
            .in1(_gnd_net_),
            .in2(N__33504),
            .in3(N__33494),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI4AJN1Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_3_14_3  (
            .in0(N__33903),
            .in1(N__33801),
            .in2(_gnd_net_),
            .in3(N__33821),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_3_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_3_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33726),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84026),
            .ce(N__37523),
            .sr(N__77291));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0IN1_16_LC_3_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0IN1_16_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0IN1_16_LC_3_14_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0IN1_16_LC_3_14_5  (
            .in0(N__35646),
            .in1(N__33705),
            .in2(_gnd_net_),
            .in3(N__33689),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0IN1Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_14_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_14_6  (
            .in0(N__33756),
            .in1(N__33747),
            .in2(_gnd_net_),
            .in3(N__33725),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGO2F3_16_LC_3_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGO2F3_16_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGO2F3_16_LC_3_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGO2F3_16_LC_3_14_7  (
            .in0(N__35645),
            .in1(N__35285),
            .in2(N__33699),
            .in3(N__33688),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGO2F3Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_3_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_3_15_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_3_15_0  (
            .in0(N__35394),
            .in1(N__35370),
            .in2(_gnd_net_),
            .in3(N__35357),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_3_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_3_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_3_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_3_15_1  (
            .in0(N__35358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84043),
            .ce(N__37521),
            .sr(N__77301));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_3_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_3_15_2 .LUT_INIT=16'b1010000011111010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_3_15_2  (
            .in0(N__33641),
            .in1(_gnd_net_),
            .in2(N__33675),
            .in3(N__33614),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_3_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_3_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_3_15_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__33642),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84043),
            .ce(N__37521),
            .sr(N__77301));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_3_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_3_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_3_15_4  (
            .in0(N__34244),
            .in1(N__34596),
            .in2(_gnd_net_),
            .in3(N__34281),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_15_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_15_5  (
            .in0(N__35603),
            .in1(N__35669),
            .in2(_gnd_net_),
            .in3(N__35629),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKNGN1_15_LC_3_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKNGN1_15_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKNGN1_15_LC_3_15_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKNGN1_15_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__33975),
            .in2(N__33969),
            .in3(N__33959),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKNGN1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIIKNU2_6_LC_3_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIKNU2_6_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIKNU2_6_LC_3_15_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIIKNU2_6_LC_3_15_7  (
            .in0(N__33942),
            .in1(N__35327),
            .in2(_gnd_net_),
            .in3(N__33929),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIIKNU2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICJKN1_18_LC_3_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICJKN1_18_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICJKN1_18_LC_3_16_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICJKN1_18_LC_3_16_0  (
            .in0(N__33879),
            .in1(N__33873),
            .in2(_gnd_net_),
            .in3(N__33851),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICJKN1Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_16_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_3_16_1  (
            .in0(N__33902),
            .in1(N__33827),
            .in2(_gnd_net_),
            .in3(N__33800),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGT7F3_18_LC_3_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGT7F3_18_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGT7F3_18_LC_3_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGT7F3_18_LC_3_16_2  (
            .in0(N__35232),
            .in1(N__33872),
            .in2(N__33858),
            .in3(N__33850),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGT7F3Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_16_3 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_3_16_3  (
            .in0(N__34279),
            .in1(N__34595),
            .in2(_gnd_net_),
            .in3(N__34245),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIV7JT5_8_LC_3_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIV7JT5_8_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIV7JT5_8_LC_3_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIV7JT5_8_LC_3_16_4  (
            .in0(N__35810),
            .in1(N__35795),
            .in2(N__33831),
            .in3(N__33779),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIV7JT5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_3_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_3_16_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__33828),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84058),
            .ce(N__37520),
            .sr(N__77311));
    defparam \pid_alt.error_d_reg_prev_esr_RNI49QU2_8_LC_3_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI49QU2_8_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI49QU2_8_LC_3_16_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI49QU2_8_LC_3_16_6  (
            .in0(N__33786),
            .in1(N__35796),
            .in2(_gnd_net_),
            .in3(N__33780),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI49QU2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_3_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_3_16_7  (
            .in0(N__34280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84058),
            .ce(N__37520),
            .sr(N__77311));
    defparam \pid_alt.error_i_acumm_prereg6_cry_0_c_LC_3_17_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_0_c_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_0_c_LC_3_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_0_c_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__34200),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_1_c_LC_3_17_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_1_c_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_1_c_LC_3_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_1_c_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__60631),
            .in2(N__36462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_0 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_2_c_LC_3_17_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_2_c_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_2_c_LC_3_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_2_c_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__34169),
            .in2(N__60652),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_1 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_3_c_LC_3_17_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_3_c_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_3_c_LC_3_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_3_c_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__60635),
            .in2(N__34152),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_2 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_4_c_inv_LC_3_17_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_4_c_inv_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_4_c_inv_LC_3_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_4_c_inv_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__34134),
            .in2(N__34098),
            .in3(N__34114),
            .lcout(\pid_alt.alt_command_i_0 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_3 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_5_c_inv_LC_3_17_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_5_c_inv_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_5_c_inv_LC_3_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_5_c_inv_LC_3_17_5  (
            .in0(N__34088),
            .in1(N__34041),
            .in2(N__34065),
            .in3(_gnd_net_),
            .lcout(\pid_alt.alt_command_i_1 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_4 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_6_c_inv_LC_3_17_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_6_c_inv_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_6_c_inv_LC_3_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_6_c_inv_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__34035),
            .in2(N__33984),
            .in3(N__34000),
            .lcout(\pid_alt.alt_command_i_2 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_5 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_7_c_inv_LC_3_17_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_7_c_inv_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_7_c_inv_LC_3_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_7_c_inv_LC_3_17_7  (
            .in0(N__34537),
            .in1(N__52770),
            .in2(N__34521),
            .in3(_gnd_net_),
            .lcout(\pid_alt.alt_command_i_3 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_6 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_8_c_inv_LC_3_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_8_c_inv_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_8_c_inv_LC_3_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_8_c_inv_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__34512),
            .in2(N__34473),
            .in3(N__34489),
            .lcout(\pid_alt.alt_command_i_4 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_9_c_inv_LC_3_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_9_c_inv_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_9_c_inv_LC_3_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_9_c_inv_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__36417),
            .in2(N__34443),
            .in3(N__34459),
            .lcout(\pid_alt.alt_command_i_5 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_8 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_10_c_inv_LC_3_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_10_c_inv_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_10_c_inv_LC_3_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_10_c_inv_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__34434),
            .in2(N__34395),
            .in3(N__34411),
            .lcout(\pid_alt.alt_command_i_6 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_9 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_11_c_inv_LC_3_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_11_c_inv_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_11_c_inv_LC_3_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_11_c_inv_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__34386),
            .in2(N__34347),
            .in3(N__34363),
            .lcout(\pid_alt.alt_command_i_7 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_10 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_12_c_LC_3_18_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_12_c_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_12_c_LC_3_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_12_c_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__34338),
            .in2(N__60653),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_11 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_13_c_LC_3_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_13_c_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_13_c_LC_3_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_13_c_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__34323),
            .in2(N__60629),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_12 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_14_c_LC_3_18_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_14_c_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_14_c_LC_3_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_14_c_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__34302),
            .in2(N__60654),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_13 ),
            .carryout(\pid_alt.error_i_acumm_prereg6_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_inv_LC_3_18_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_inv_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_inv_LC_3_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_15_c_inv_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__34692),
            .in2(_gnd_net_),
            .in3(N__52880),
            .lcout(\pid_alt.drone_altitude_i_15 ),
            .ltout(),
            .carryin(\pid_alt.error_i_acumm_prereg6_cry_14 ),
            .carryout(\pid_alt.error_i_acumm_prereg6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIT0JE2_LC_3_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIT0JE2_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIT0JE2_LC_3_19_0 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIT0JE2_LC_3_19_0  (
            .in0(N__34686),
            .in1(N__34677),
            .in2(N__50068),
            .in3(N__34671),
            .lcout(\pid_alt.error_i_acumm_prereg_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIQDPN2_LC_3_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIQDPN2_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIQDPN2_LC_3_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg6_cry_15_c_RNIQDPN2_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__54983),
            .in2(_gnd_net_),
            .in3(N__34668),
            .lcout(\pid_alt.error_i_acumm_prereg_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_3_19_2 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_3_19_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_3_19_2  (
            .in0(N__50061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77632),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_3_19_3 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_3_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47685),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84095),
            .ce(N__34614),
            .sr(N__77332));
    defparam \pid_alt.error_p_reg_esr_8_LC_3_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_3_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_3_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_3_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34608),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84108),
            .ce(N__36280),
            .sr(N__82874));
    defparam \pid_alt.error_p_reg_esr_7_LC_3_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_3_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_3_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_3_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34572),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84108),
            .ce(N__36280),
            .sr(N__82874));
    defparam \pid_alt.error_d_reg_esr_1_LC_4_7_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_4_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34560),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83910),
            .ce(N__36269),
            .sr(N__82889));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35415),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83921),
            .ce(N__37532),
            .sr(N__77249));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_9_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__34868),
            .in2(_gnd_net_),
            .in3(N__34853),
            .lcout(),
            .ltout(\pid_alt.m21_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_9_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_4_9_2  (
            .in0(N__34842),
            .in1(N__46572),
            .in2(N__34821),
            .in3(N__37012),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_9_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_9_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_9_3  (
            .in0(N__34765),
            .in1(N__34735),
            .in2(_gnd_net_),
            .in3(N__34715),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_10_1 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_10_1  (
            .in0(N__34805),
            .in1(N__34772),
            .in2(N__34794),
            .in3(N__34785),
            .lcout(),
            .ltout(\pid_alt.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_10_2 .C_ON=1'b0;
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_10_2 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \pid_alt.state_RNIAAPN5_1_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__47721),
            .in2(N__34779),
            .in3(N__54968),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(\pid_alt.un1_reset_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIVV066_1_LC_4_10_3 .C_ON=1'b0;
    defparam \pid_alt.state_RNIVV066_1_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIVV066_1_LC_4_10_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_alt.state_RNIVV066_1_LC_4_10_3  (
            .in0(N__47722),
            .in1(_gnd_net_),
            .in2(N__34776),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_76_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_13_LC_4_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_4_10_5 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_4_10_5  (
            .in0(N__34773),
            .in1(N__34739),
            .in2(_gnd_net_),
            .in3(N__34719),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83947),
            .ce(N__36922),
            .sr(N__46490));
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6  (
            .in0(N__36765),
            .in1(N__47720),
            .in2(N__37150),
            .in3(N__54967),
            .lcout(),
            .ltout(\pid_alt.un1_reset_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_7 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_7  (
            .in0(N__37202),
            .in1(N__36621),
            .in2(N__34962),
            .in3(N__37259),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_11_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__39806),
            .in2(N__39810),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_4_11_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__35445),
            .in2(N__35480),
            .in3(N__34959),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_1_LC_4_11_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__35505),
            .in2(N__35538),
            .in3(N__34956),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_2_LC_4_11_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__36099),
            .in2(N__36137),
            .in3(N__34953),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_3_LC_4_11_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__36000),
            .in2(N__36038),
            .in3(N__34950),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_4_LC_4_11_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__35978),
            .in2(N__34947),
            .in3(N__34938),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_5_LC_4_11_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(N__34935),
            .in2(N__34928),
            .in3(N__34911),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_6_LC_4_11_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(N__34908),
            .in2(N__34892),
            .in3(N__34875),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__83962),
            .ce(N__37529),
            .sr(N__77265));
    defparam \pid_alt.pid_prereg_esr_7_LC_4_12_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__35127),
            .in2(N__35115),
            .in3(N__35094),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_8_LC_4_12_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__35880),
            .in2(N__35909),
            .in3(N__35091),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_9_LC_4_12_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__35088),
            .in2(N__35817),
            .in3(N__35076),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_10_LC_4_12_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__35073),
            .in2(N__35067),
            .in3(N__35046),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_11_LC_4_12_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__35043),
            .in2(N__35036),
            .in3(N__35019),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_12_LC_4_12_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__35015),
            .in2(N__35004),
            .in3(N__34995),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_13_LC_4_12_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__34992),
            .in2(N__34985),
            .in3(N__34968),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_14_LC_4_12_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__37581),
            .in2(N__37601),
            .in3(N__34965),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__83978),
            .ce(N__37526),
            .sr(N__77272));
    defparam \pid_alt.pid_prereg_esr_15_LC_4_13_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__36906),
            .in2(N__37431),
            .in3(N__35313),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_16_LC_4_13_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__35310),
            .in2(N__37737),
            .in3(N__35298),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_17_LC_4_13_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__35295),
            .in2(N__35289),
            .in3(N__35271),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_18_LC_4_13_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__35268),
            .in2(N__35261),
            .in3(N__35244),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_19_LC_4_13_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__35241),
            .in2(N__35231),
            .in3(N__35214),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_20_LC_4_13_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__35211),
            .in2(N__35198),
            .in3(N__35175),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_21_LC_4_13_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__35172),
            .in2(N__35160),
            .in3(N__35145),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_22_LC_4_13_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__35142),
            .in2(N__35592),
            .in3(N__35130),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__83994),
            .ce(N__37524),
            .sr(N__77277));
    defparam \pid_alt.pid_prereg_esr_23_LC_4_14_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__35588),
            .in2(N__35568),
            .in3(N__35556),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__84013),
            .ce(N__37522),
            .sr(N__77282));
    defparam \pid_alt.pid_prereg_esr_24_LC_4_14_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__35553),
            .in2(_gnd_net_),
            .in3(N__35541),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84013),
            .ce(N__37522),
            .sr(N__77282));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_4_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_4_15_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__35453),
            .in2(_gnd_net_),
            .in3(N__35407),
            .lcout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ),
            .ltout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3RCL2_1_LC_4_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3RCL2_1_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3RCL2_1_LC_4_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3RCL2_1_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__35537),
            .in2(N__35508),
            .in3(N__36162),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3RCL2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_4_15_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_4_15_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_4_15_2  (
            .in0(N__58410),
            .in1(N__39753),
            .in2(_gnd_net_),
            .in3(N__58305),
            .lcout(\dron_frame_decoder_1.state_ns_i_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_0_LC_4_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_4_15_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__35496),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84027),
            .ce(N__36277),
            .sr(N__82883));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_15_4  (
            .in0(N__35484),
            .in1(N__35454),
            .in2(_gnd_net_),
            .in3(N__35408),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_0_LC_4_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35433),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84027),
            .ce(N__36277),
            .sr(N__82883));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_15_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_4_15_6  (
            .in0(N__35393),
            .in1(N__35369),
            .in2(_gnd_net_),
            .in3(N__35356),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_4_16_0  (
            .in0(N__36293),
            .in1(N__35786),
            .in2(_gnd_net_),
            .in3(N__35776),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_4_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_4_16_1  (
            .in0(N__35778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84044),
            .ce(N__37518),
            .sr(N__77302));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_4_16_2  (
            .in0(N__36294),
            .in1(N__35787),
            .in2(_gnd_net_),
            .in3(N__35777),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_4_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_4_16_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_4_16_3  (
            .in0(N__35741),
            .in1(N__35684),
            .in2(_gnd_net_),
            .in3(N__35714),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_4_16_4  (
            .in0(N__35715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84044),
            .ce(N__37518),
            .sr(N__77302));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_16_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_4_16_5  (
            .in0(N__35670),
            .in1(N__35604),
            .in2(_gnd_net_),
            .in3(N__35630),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_4_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_4_16_6  (
            .in0(N__35631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84044),
            .ce(N__37518),
            .sr(N__77302));
    defparam \pid_front.error_axb_8_l_ofx_LC_4_16_7 .C_ON=1'b0;
    defparam \pid_front.error_axb_8_l_ofx_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_8_l_ofx_LC_4_16_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_front.error_axb_8_l_ofx_LC_4_16_7  (
            .in0(N__49727),
            .in1(N__48153),
            .in2(_gnd_net_),
            .in3(N__48122),
            .lcout(\pid_front.error_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9F5Q6_2_LC_4_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9F5Q6_2_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9F5Q6_2_LC_4_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9F5Q6_2_LC_4_17_0  (
            .in0(N__35963),
            .in1(N__35991),
            .in2(N__36045),
            .in3(N__36227),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9F5Q6Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_4_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_4_17_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_4_17_1  (
            .in0(N__36324),
            .in1(N__36057),
            .in2(_gnd_net_),
            .in3(N__36085),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_4_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_4_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_4_17_2  (
            .in0(N__35964),
            .in1(_gnd_net_),
            .in2(N__35985),
            .in3(N__36228),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_17_3  (
            .in0(N__35953),
            .in1(N__36347),
            .in2(_gnd_net_),
            .in3(N__35933),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35955),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84059),
            .ce(N__37517),
            .sr(N__77312));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_17_5 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_17_5  (
            .in0(N__35954),
            .in1(N__36348),
            .in2(_gnd_net_),
            .in3(N__35934),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDJGT5_7_LC_4_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDJGT5_7_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDJGT5_7_LC_4_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDJGT5_7_LC_4_17_6  (
            .in0(N__35828),
            .in1(N__35840),
            .in2(N__35910),
            .in3(N__35867),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDJGT5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUOU2_7_LC_4_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUOU2_7_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRUOU2_7_LC_4_17_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIRUOU2_7_LC_4_17_7  (
            .in0(N__35868),
            .in1(_gnd_net_),
            .in2(N__35844),
            .in3(N__35829),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIRUOU2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_4_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_4_18_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_4_18_0  (
            .in0(N__36373),
            .in1(N__36190),
            .in2(_gnd_net_),
            .in3(N__36210),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_4_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_4_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_4_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_4_18_1  (
            .in0(N__36213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84077),
            .ce(N__37516),
            .sr(N__77318));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_4_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_4_18_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_4_18_2  (
            .in0(N__36374),
            .in1(N__36191),
            .in2(_gnd_net_),
            .in3(N__36211),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_4_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_4_18_3 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_4_18_3  (
            .in0(N__36219),
            .in1(N__36157),
            .in2(N__36231),
            .in3(N__36173),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_18_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_18_4  (
            .in0(N__36323),
            .in1(N__36056),
            .in2(_gnd_net_),
            .in3(N__36086),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_4_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_4_18_5 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_4_18_5  (
            .in0(N__36212),
            .in1(N__36192),
            .in2(N__36177),
            .in3(N__36375),
            .lcout(),
            .ltout(\pid_alt.un1_pid_prereg_16_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI32PN4_1_LC_4_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI32PN4_1_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI32PN4_1_LC_4_18_6 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI32PN4_1_LC_4_18_6  (
            .in0(N__36174),
            .in1(N__36161),
            .in2(N__36141),
            .in3(N__36138),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI32PN4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_4_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_4_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_4_18_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_4_18_7  (
            .in0(N__36087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84077),
            .ce(N__37516),
            .sr(N__77318));
    defparam \dron_frame_decoder_1.state_RNIRK8L_5_LC_4_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIRK8L_5_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIRK8L_5_LC_4_19_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \dron_frame_decoder_1.state_RNIRK8L_5_LC_4_19_1  (
            .in0(N__71893),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58037),
            .lcout(\dron_frame_decoder_1.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_1_LC_4_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_1_LC_4_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_1_LC_4_19_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_1_LC_4_19_2  (
            .in0(N__36455),
            .in1(N__52825),
            .in2(N__58484),
            .in3(N__57995),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84088),
            .ce(),
            .sr(N__77325));
    defparam \pid_alt.error_axb_1_LC_4_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_4_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36454),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_9_LC_4_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_9_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_9_LC_4_19_4 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_9_LC_4_19_4  (
            .in0(N__36416),
            .in1(N__52826),
            .in2(N__58485),
            .in3(N__57996),
            .lcout(drone_altitude_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84088),
            .ce(),
            .sr(N__77325));
    defparam \dron_frame_decoder_1.source_H_disp_side_1_LC_4_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_1_LC_4_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_1_LC_4_19_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_1_LC_4_19_5  (
            .in0(N__36426),
            .in1(N__58342),
            .in2(N__71911),
            .in3(N__57997),
            .lcout(drone_H_disp_side_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84088),
            .ce(),
            .sr(N__77325));
    defparam \pid_side.error_axb_1_LC_4_19_6 .C_ON=1'b0;
    defparam \pid_side.error_axb_1_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_1_LC_4_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_1_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36425),
            .lcout(\pid_side.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_RNID543_9_LC_4_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNID543_9_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNID543_9_LC_4_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNID543_9_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36415),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_1_LC_4_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_4_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_4_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36390),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84096),
            .ce(N__36278),
            .sr(N__82880));
    defparam \pid_alt.error_p_reg_esr_3_LC_4_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_4_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36360),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84096),
            .ce(N__36278),
            .sr(N__82880));
    defparam \pid_alt.error_p_reg_esr_2_LC_4_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_4_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_4_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36336),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84096),
            .ce(N__36278),
            .sr(N__82880));
    defparam \pid_alt.error_p_reg_esr_9_LC_4_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_4_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_4_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36306),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84105),
            .ce(N__36279),
            .sr(N__82872));
    defparam \pid_alt.state_RNICP2N1_0_LC_5_4_5 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_5_4_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__36636),
            .in2(_gnd_net_),
            .in3(N__83002),
            .lcout(\pid_alt.N_579_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_5_5_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_5_5_6 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_5_5_6  (
            .in0(N__37854),
            .in1(N__48349),
            .in2(N__37790),
            .in3(N__77662),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83875),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_5_5_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_5_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__37783),
            .in2(_gnd_net_),
            .in3(N__37853),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_6_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__36487),
            .in2(_gnd_net_),
            .in3(N__36501),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_5_6_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_5_6_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_5_6_3  (
            .in0(N__77614),
            .in1(N__36557),
            .in2(N__36507),
            .in3(N__38033),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83886),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_6_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_6_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_5_6_6  (
            .in0(N__38950),
            .in1(N__38095),
            .in2(N__36606),
            .in3(N__77612),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_5_6_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_5_6_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_5_6_7  (
            .in0(N__77613),
            .in1(N__36556),
            .in2(N__36504),
            .in3(N__36488),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83886),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_7_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_7_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_5_7_0  (
            .in0(N__36486),
            .in1(N__36500),
            .in2(N__36489),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_7_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__38192),
            .in2(_gnd_net_),
            .in3(N__36465),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_7_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__38144),
            .in2(_gnd_net_),
            .in3(N__36582),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_7_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__38102),
            .in2(_gnd_net_),
            .in3(N__36579),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_5_7_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_5_7_4 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.timer_Count_4_LC_5_7_4  (
            .in0(N__77640),
            .in1(N__36555),
            .in2(N__36576),
            .in3(N__38032),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83897),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_7_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_7_5 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_5_7_5  (
            .in0(N__38145),
            .in1(N__38906),
            .in2(N__37989),
            .in3(N__38101),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(\uart_pc.timer_Count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_5_7_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_5_7_6 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_pc.timer_Count_3_LC_5_7_6  (
            .in0(N__77639),
            .in1(N__36573),
            .in2(N__36567),
            .in3(N__38031),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83897),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_5_7_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_5_7_7 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.timer_Count_2_LC_5_7_7  (
            .in0(N__38030),
            .in1(N__36564),
            .in2(N__36558),
            .in3(N__77641),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83897),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_8_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__38188),
            .in2(_gnd_net_),
            .in3(N__38143),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_8_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_8_3 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_5_8_3  (
            .in0(N__38951),
            .in1(N__36537),
            .in2(N__36531),
            .in3(N__38910),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_5_8_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_5_8_4 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_5_8_4  (
            .in0(N__38222),
            .in1(N__39401),
            .in2(_gnd_net_),
            .in3(N__77634),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_5_8_5 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_5_8_5 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart_pc.state_0_LC_5_8_5  (
            .in0(N__38952),
            .in1(N__36602),
            .in2(N__36588),
            .in3(N__38103),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83911),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_10_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_10_1 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_10_1  (
            .in0(N__37086),
            .in1(N__37206),
            .in2(N__37160),
            .in3(N__37260),
            .lcout(\pid_alt.source_pid_9_0_tz_6 ),
            .ltout(\pid_alt.source_pid_9_0_tz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_11_LC_5_10_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_5_10_2 .LUT_INIT=16'b1101111110001010;
    LogicCell40 \pid_alt.source_pid_1_11_LC_5_10_2  (
            .in0(N__47701),
            .in1(N__36816),
            .in2(N__36585),
            .in3(N__50734),
            .lcout(throttle_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83935),
            .ce(),
            .sr(N__38481));
    defparam \pid_alt.source_pid_1_6_LC_5_10_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_5_10_3 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_6_LC_5_10_3  (
            .in0(N__38534),
            .in1(N__47699),
            .in2(N__50635),
            .in3(N__36831),
            .lcout(throttle_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83935),
            .ce(),
            .sr(N__38481));
    defparam \pid_alt.source_pid_1_7_LC_5_10_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_5_10_4 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_7_LC_5_10_4  (
            .in0(N__47697),
            .in1(N__38535),
            .in2(N__50827),
            .in3(N__36873),
            .lcout(throttle_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83935),
            .ce(),
            .sr(N__38481));
    defparam \pid_alt.source_pid_1_8_LC_5_10_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_5_10_5 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_8_LC_5_10_5  (
            .in0(N__38536),
            .in1(N__47700),
            .in2(N__54407),
            .in3(N__36891),
            .lcout(throttle_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83935),
            .ce(),
            .sr(N__38481));
    defparam \pid_alt.source_pid_1_9_LC_5_10_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_5_10_6 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_9_LC_5_10_6  (
            .in0(N__47698),
            .in1(N__38537),
            .in2(N__47111),
            .in3(N__36852),
            .lcout(throttle_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83935),
            .ce(),
            .sr(N__38481));
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_10_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIOVDUE_1_LC_5_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIOVDUE_1_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__47696),
            .in2(_gnd_net_),
            .in3(N__38461),
            .lcout(\pid_alt.N_76_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_11_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_5_11_0  (
            .in0(N__36692),
            .in1(N__36644),
            .in2(N__36681),
            .in3(N__36704),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_11_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_11_1 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG2382_12_LC_5_11_1  (
            .in0(N__36777),
            .in1(N__37192),
            .in2(_gnd_net_),
            .in3(N__37081),
            .lcout(\pid_alt.N_44 ),
            .ltout(\pid_alt.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_11_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_11_2 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__37383),
            .in2(N__36711),
            .in3(N__37346),
            .lcout(\pid_alt.N_46 ),
            .ltout(\pid_alt.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_1_LC_5_11_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_1_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_1_LC_5_11_3 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_1_LC_5_11_3  (
            .in0(N__37256),
            .in1(N__37155),
            .in2(N__36708),
            .in3(N__36705),
            .lcout(throttle_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83948),
            .ce(N__37055),
            .sr(N__38489));
    defparam \pid_alt.source_pid_1_esr_2_LC_5_11_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_2_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_2_LC_5_11_4 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_2_LC_5_11_4  (
            .in0(N__37154),
            .in1(N__36693),
            .in2(N__36665),
            .in3(N__37257),
            .lcout(throttle_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83948),
            .ce(N__37055),
            .sr(N__38489));
    defparam \pid_alt.source_pid_1_esr_3_LC_5_11_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_3_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_3_LC_5_11_5 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \pid_alt.source_pid_1_esr_3_LC_5_11_5  (
            .in0(N__37258),
            .in1(N__36680),
            .in2(N__36666),
            .in3(N__37159),
            .lcout(throttle_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83948),
            .ce(N__37055),
            .sr(N__38489));
    defparam \pid_alt.source_pid_1_esr_0_LC_5_11_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_0_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_0_LC_5_11_6 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_0_LC_5_11_6  (
            .in0(N__36658),
            .in1(N__36645),
            .in2(N__37161),
            .in3(N__37255),
            .lcout(throttle_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83948),
            .ce(N__37055),
            .sr(N__38489));
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_11_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_5_11_7 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_5_11_7  (
            .in0(N__67379),
            .in1(N__47686),
            .in2(N__50057),
            .in3(N__77589),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_12_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_12_0  (
            .in0(N__36612),
            .in1(N__36809),
            .in2(N__38513),
            .in3(N__47688),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_5_12_1  (
            .in0(N__36789),
            .in1(N__37382),
            .in2(N__36624),
            .in3(N__37345),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_12_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_12_2  (
            .in0(N__36830),
            .in1(N__36887),
            .in2(N__36872),
            .in3(N__36847),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_5_12_3  (
            .in0(N__36886),
            .in1(N__36865),
            .in2(N__36851),
            .in3(N__36829),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_4 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__36808),
            .in2(N__36795),
            .in3(N__38506),
            .lcout(\pid_alt.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_12_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__37077),
            .in2(_gnd_net_),
            .in3(N__36749),
            .lcout(\pid_alt.N_90 ),
            .ltout(\pid_alt.N_90_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_5_12_6  (
            .in0(N__37201),
            .in1(N__37344),
            .in2(N__36792),
            .in3(N__47687),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_5_12_7  (
            .in0(N__36788),
            .in1(N__37230),
            .in2(N__36780),
            .in3(N__36776),
            .lcout(\pid_alt.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_5_13_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_5_13_0  (
            .in0(N__37248),
            .in1(N__37320),
            .in2(N__37149),
            .in3(N__36756),
            .lcout(throttle_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83979),
            .ce(N__37056),
            .sr(N__38490));
    defparam \pid_alt.pid_prereg_esr_RNI7OVM_19_LC_5_13_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI7OVM_19_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI7OVM_19_LC_5_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI7OVM_19_LC_5_13_1  (
            .in0(N__36738),
            .in1(N__36732),
            .in2(N__36726),
            .in3(N__36717),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_5_13_2 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_5_13_2  (
            .in0(N__37246),
            .in1(_gnd_net_),
            .in2(N__37148),
            .in3(N__37199),
            .lcout(throttle_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83979),
            .ce(N__37056),
            .sr(N__38490));
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \pid_alt.source_pid_1_esr_RNO_0_4_LC_5_13_3  (
            .in0(N__37381),
            .in1(N__37125),
            .in2(N__37359),
            .in3(N__37245),
            .lcout(),
            .ltout(\pid_alt.source_pid_9_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_5_13_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_5_13_4  (
            .in0(N__37247),
            .in1(N__37358),
            .in2(N__37323),
            .in3(N__37319),
            .lcout(throttle_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83979),
            .ce(N__37056),
            .sr(N__38490));
    defparam \pid_alt.pid_prereg_esr_RNIFUTM_14_LC_5_13_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFUTM_14_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFUTM_14_LC_5_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFUTM_14_LC_5_13_5  (
            .in0(N__37308),
            .in1(N__37302),
            .in2(N__37296),
            .in3(N__37287),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_15_LC_5_13_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_15_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_15_LC_5_13_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT4CP1_15_LC_5_13_6  (
            .in0(N__37281),
            .in1(N__37275),
            .in2(N__37269),
            .in3(N__37266),
            .lcout(\pid_alt.N_216 ),
            .ltout(\pid_alt.N_216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_12_LC_5_13_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_5_13_7 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_5_13_7  (
            .in0(N__37200),
            .in1(N__37126),
            .in2(N__37089),
            .in3(N__37082),
            .lcout(throttle_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83979),
            .ce(N__37056),
            .sr(N__38490));
    defparam \pid_alt.error_i_acumm_esr_4_LC_5_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_5_14_0 .LUT_INIT=16'b1011101010111111;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_5_14_0  (
            .in0(N__37041),
            .in1(N__46640),
            .in2(N__46595),
            .in3(N__36996),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83995),
            .ce(N__36936),
            .sr(N__46514));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGJTE3_14_LC_5_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGJTE3_14_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGJTE3_14_LC_5_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGJTE3_14_LC_5_15_0  (
            .in0(N__36897),
            .in1(N__37631),
            .in2(N__37430),
            .in3(N__37760),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGJTE3Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_15_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_15_1  (
            .in0(N__37568),
            .in1(_gnd_net_),
            .in2(N__37545),
            .in3(N__37623),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICEFN1_14_LC_5_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICEFN1_14_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICEFN1_14_LC_5_15_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICEFN1_14_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__37632),
            .in2(N__37764),
            .in3(N__37761),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICEFN1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_15_3  (
            .in0(N__37715),
            .in1(N__37692),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_15_4  (
            .in0(N__37622),
            .in1(N__37541),
            .in2(_gnd_net_),
            .in3(N__37567),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK5TH3_13_LC_5_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK5TH3_13_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK5TH3_13_LC_5_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK5TH3_13_LC_5_15_5  (
            .in0(N__37605),
            .in1(N__37466),
            .in2(N__37584),
            .in3(N__37456),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK5TH3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37569),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84014),
            .ce(N__37519),
            .sr(N__77283));
    defparam \pid_alt.error_d_reg_prev_esr_RNI45EN1_13_LC_5_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI45EN1_13_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI45EN1_13_LC_5_15_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI45EN1_13_LC_5_15_7  (
            .in0(N__37473),
            .in1(N__37467),
            .in2(_gnd_net_),
            .in3(N__37457),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI45EN1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_5_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_5_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64985),
            .lcout(drone_H_disp_front_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84028),
            .ce(N__38628),
            .sr(N__77292));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_17_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__38400),
            .in2(_gnd_net_),
            .in3(N__77619),
            .lcout(\Commands_frame_decoder.source_CH1data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_0_LC_5_18_2 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_5_18_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_5_18_2  (
            .in0(N__50042),
            .in1(N__67378),
            .in2(_gnd_net_),
            .in3(N__47732),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84060),
            .ce(),
            .sr(N__77313));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_18_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_18_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_5_18_6  (
            .in0(N__37823),
            .in1(N__48348),
            .in2(N__39672),
            .in3(N__79277),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84060),
            .ce(),
            .sr(N__77313));
    defparam \reset_module_System.reset_LC_7_1_6 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_7_1_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_7_1_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_7_1_6  (
            .in0(N__40676),
            .in1(N__39015),
            .in2(_gnd_net_),
            .in3(N__38982),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83826),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_7_4_0 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40575),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83848),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_7_4_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_7_4_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI6QPK_14_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__37846),
            .in2(_gnd_net_),
            .in3(N__37922),
            .lcout(\Commands_frame_decoder.N_369_2 ),
            .ltout(\Commands_frame_decoder.N_369_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_4_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_7_4_3 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_7_4_3  (
            .in0(N__38064),
            .in1(N__37947),
            .in2(N__37809),
            .in3(N__37885),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_370_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_4_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_7_4_4 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_7_4_4  (
            .in0(N__38715),
            .in1(N__37940),
            .in2(N__37806),
            .in3(N__37803),
            .lcout(\Commands_frame_decoder.state_ns_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_4_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_4_7 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_4_7  (
            .in0(N__37847),
            .in1(N__48283),
            .in2(N__37797),
            .in3(N__38714),
            .lcout(\Commands_frame_decoder.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_7_5_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_7_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_7_5_1  (
            .in0(N__79198),
            .in1(N__73692),
            .in2(N__48316),
            .in3(N__38052),
            .lcout(\Commands_frame_decoder.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_7_5_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_7_5_4 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_7_5_4 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \Commands_frame_decoder.state_0_LC_7_5_4  (
            .in0(N__40202),
            .in1(N__37770),
            .in2(N__37923),
            .in3(N__37865),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83857),
            .ce(),
            .sr(N__77246));
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_7_5_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_7_5_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Commands_frame_decoder.state_RNO_4_0_LC_7_5_5  (
            .in0(N__80203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80413),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_7_5_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_7_5_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_7_5_6  (
            .in0(N__79864),
            .in1(N__80074),
            .in2(N__37950),
            .in3(N__37913),
            .lcout(\Commands_frame_decoder.N_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_7_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_7_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_1_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__79865),
            .in2(_gnd_net_),
            .in3(N__80432),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_7_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_7_6_1  (
            .in0(N__80044),
            .in1(N__37941),
            .in2(N__37929),
            .in3(N__80204),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_LC_7_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_7_6_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_7_6_2  (
            .in0(N__37918),
            .in1(N__37886),
            .in2(N__37926),
            .in3(N__40177),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83866),
            .ce(),
            .sr(N__77247));
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_7_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_2_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__79866),
            .in2(_gnd_net_),
            .in3(N__80433),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_6_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_7_6_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_2_LC_7_6_5  (
            .in0(N__80045),
            .in1(N__37917),
            .in2(N__37890),
            .in3(N__80205),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_2_LC_7_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_7_6_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_7_6_6  (
            .in0(N__38414),
            .in1(N__37887),
            .in2(N__37872),
            .in3(N__40178),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83866),
            .ce(),
            .sr(N__77247));
    defparam \Commands_frame_decoder.state_14_LC_7_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_14_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_14_LC_7_6_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_14_LC_7_6_7  (
            .in0(N__48333),
            .in1(N__38565),
            .in2(_gnd_net_),
            .in3(N__37869),
            .lcout(\Commands_frame_decoder.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83866),
            .ce(),
            .sr(N__77247));
    defparam \uart_pc.state_4_LC_7_7_0 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_7_7_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \uart_pc.state_4_LC_7_7_0  (
            .in0(N__38902),
            .in1(N__38007),
            .in2(N__38040),
            .in3(N__77660),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_7_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_7_7_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_7_7_1  (
            .in0(N__39281),
            .in1(N__38159),
            .in2(_gnd_net_),
            .in3(N__38111),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_7_7_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_7_7_2 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_drone.timer_Count_0_LC_7_7_2  (
            .in0(N__38831),
            .in1(N__42352),
            .in2(N__42324),
            .in3(N__77658),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_7_7_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_7_7_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_7_7_3  (
            .in0(N__38160),
            .in1(N__38901),
            .in2(N__37988),
            .in3(N__38112),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_7_7_4 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_7_7_4 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_pc.state_3_LC_7_7_4  (
            .in0(N__37984),
            .in1(N__38006),
            .in2(N__37998),
            .in3(N__77659),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_7_7_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_7_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__38830),
            .in2(_gnd_net_),
            .in3(N__38844),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_7_7_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_7_7_6 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_7_7_6  (
            .in0(N__42323),
            .in1(N__42353),
            .in2(N__37995),
            .in3(N__77661),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83876),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_7_7_7 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_7_7_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \reset_module_System.count_1_LC_7_7_7  (
            .in0(N__40686),
            .in1(N__39006),
            .in2(N__40677),
            .in3(N__38978),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_2_LC_7_8_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_7_8_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_7_8_0  (
            .in0(N__37980),
            .in1(N__39377),
            .in2(N__38211),
            .in3(N__77627),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_7_8_1 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_7_8_1 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_pc.state_2_LC_7_8_1  (
            .in0(N__38167),
            .in1(N__38209),
            .in2(N__37992),
            .in3(N__38115),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83887),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_7_8_2 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_7_8_2 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_7_8_2  (
            .in0(N__38210),
            .in1(N__39378),
            .in2(N__38229),
            .in3(N__77628),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83887),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_7_8_3  (
            .in0(N__38931),
            .in1(N__38196),
            .in2(N__38169),
            .in3(N__38113),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(\uart_pc.data_rdyc_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_8_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_7_8_4 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__39376),
            .in2(N__38172),
            .in3(N__77626),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_7_8_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_8_5 .LUT_INIT=16'b0101000100010001;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_7_8_5  (
            .in0(N__38930),
            .in1(N__38885),
            .in2(N__38168),
            .in3(N__38114),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_7_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_7_8_6  (
            .in0(N__80003),
            .in1(N__80187),
            .in2(N__79837),
            .in3(N__80395),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_7_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_7_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__80982),
            .in2(_gnd_net_),
            .in3(N__79630),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__39037),
            .in2(_gnd_net_),
            .in3(N__77625),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_7_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_7_9_1 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \uart_pc.data_3_LC_7_9_1  (
            .in0(N__39072),
            .in1(N__39200),
            .in2(N__38043),
            .in3(N__79684),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83898),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_7_9_2 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_7_9_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_2_LC_7_9_2  (
            .in0(N__39199),
            .in1(N__39167),
            .in2(N__39096),
            .in3(N__80199),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83898),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_9_4 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_7_9_4  (
            .in0(N__39583),
            .in1(N__39485),
            .in2(_gnd_net_),
            .in3(N__39528),
            .lcout(\uart_pc.N_152 ),
            .ltout(\uart_pc.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_7_9_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_7_9_5 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__38249),
            .in2(N__38268),
            .in3(N__38903),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_7_9_6 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_7_9_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_0_LC_7_9_6  (
            .in0(N__39198),
            .in1(N__39166),
            .in2(N__39141),
            .in3(N__80412),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83898),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_0_LC_7_10_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_7_10_1 .LUT_INIT=16'b0000111100100000;
    LogicCell40 \uart_pc.bit_Count_0_LC_7_10_1  (
            .in0(N__38905),
            .in1(N__39280),
            .in2(N__38262),
            .in3(N__39490),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83912),
            .ce(),
            .sr(N__77252));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_10_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_7_10_2  (
            .in0(N__39489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38257),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_7_10_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_7_10_3 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_7_10_3  (
            .in0(N__38238),
            .in1(N__39591),
            .in2(N__38265),
            .in3(N__39537),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83912),
            .ce(),
            .sr(N__77252));
    defparam \uart_pc.bit_Count_1_LC_7_10_4 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_7_10_4 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_1_LC_7_10_4  (
            .in0(N__39491),
            .in1(N__38261),
            .in2(N__39545),
            .in3(N__38237),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83912),
            .ce(),
            .sr(N__77252));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_7_10_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_7_10_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_7_10_5  (
            .in0(N__39585),
            .in1(N__39529),
            .in2(_gnd_net_),
            .in3(N__39486),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_7_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_7_10_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_7_10_6  (
            .in0(N__39487),
            .in1(_gnd_net_),
            .in2(N__39544),
            .in3(N__39586),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_7_10_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_7_10_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_7_10_7  (
            .in0(N__39584),
            .in1(N__39533),
            .in2(_gnd_net_),
            .in3(N__39488),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_rdy_LC_7_11_1 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_7_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__39405),
            .in2(_gnd_net_),
            .in3(N__39042),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83922),
            .ce(),
            .sr(N__77258));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__38415),
            .in2(_gnd_net_),
            .in3(N__48236),
            .lcout(\Commands_frame_decoder.source_CH1data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH1data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_3_LC_7_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_7_11_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_3_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__38382),
            .in2(N__38385),
            .in3(N__40221),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83922),
            .ce(),
            .sr(N__77258));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_11_6  (
            .in0(N__48237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38381),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \Commands_frame_decoder.state_4_LC_7_11_7  (
            .in0(N__40222),
            .in1(_gnd_net_),
            .in2(N__38373),
            .in3(N__39219),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83922),
            .ce(),
            .sr(N__77258));
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_4_LC_7_12_0  (
            .in0(N__48269),
            .in1(N__38341),
            .in2(N__41193),
            .in3(N__79227),
            .lcout(xy_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83936),
            .ce(),
            .sr(N__77266));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_12_3 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_7_12_3  (
            .in0(N__39654),
            .in1(_gnd_net_),
            .in2(N__77664),
            .in3(N__48266),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_7_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_7_12_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_7_12_4  (
            .in0(N__48268),
            .in1(N__77600),
            .in2(_gnd_net_),
            .in3(N__39703),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_7_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_7_12_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_7_12_5  (
            .in0(N__39718),
            .in1(_gnd_net_),
            .in2(N__77665),
            .in3(N__48267),
            .lcout(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_7_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_7_12_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_RNITUI31_13_LC_7_12_6  (
            .in0(N__48265),
            .in1(N__77593),
            .in2(_gnd_net_),
            .in3(N__38557),
            .lcout(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_13_LC_7_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_13_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_13_LC_7_12_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_13_LC_7_12_7  (
            .in0(N__38558),
            .in1(N__48168),
            .in2(_gnd_net_),
            .in3(N__40223),
            .lcout(\Commands_frame_decoder.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83936),
            .ce(),
            .sr(N__77266));
    defparam \pid_alt.source_pid_1_10_LC_7_13_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_7_13_5 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_10_LC_7_13_5  (
            .in0(N__38544),
            .in1(N__47683),
            .in2(N__50869),
            .in3(N__38517),
            .lcout(throttle_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83949),
            .ce(),
            .sr(N__38488));
    defparam \pid_front.error_p_reg_esr_0_LC_7_14_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_0_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_0_LC_7_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_0_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38445),
            .lcout(\pid_front.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83963),
            .ce(N__83106),
            .sr(N__82882));
    defparam \pid_front.error_p_reg_esr_3_LC_7_14_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_3_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_3_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_3_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38433),
            .lcout(\pid_front.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83963),
            .ce(N__83106),
            .sr(N__82882));
    defparam \dron_frame_decoder_1.WDT_RNIG3NH2_15_LC_7_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIG3NH2_15_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIG3NH2_15_LC_7_15_0 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIG3NH2_15_LC_7_15_0  (
            .in0(N__39633),
            .in1(N__41235),
            .in2(N__41439),
            .in3(N__41277),
            .lcout(\dron_frame_decoder_1.WDT10_0 ),
            .ltout(\dron_frame_decoder_1.WDT10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_0_LC_7_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_7_15_1 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_7_15_1 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_7_15_1  (
            .in0(N__58264),
            .in1(N__39752),
            .in2(N__38418),
            .in3(N__39849),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_7_LC_7_15_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_7_15_2 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_7_15_2  (
            .in0(N__71876),
            .in1(N__58276),
            .in2(N__38600),
            .in3(N__51406),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_6_LC_7_15_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_7_15_3 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_7_15_3  (
            .in0(N__51405),
            .in1(N__38593),
            .in2(N__58303),
            .in3(N__58389),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_4_LC_7_15_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_7_15_4 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_7_15_4  (
            .in0(N__71875),
            .in1(N__58269),
            .in2(N__58036),
            .in3(N__51403),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_5_LC_7_15_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_7_15_5 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_7_15_5  (
            .in0(N__51404),
            .in1(N__53235),
            .in2(N__58302),
            .in3(N__58029),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_2_LC_7_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_7_15_6 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_7_15_6  (
            .in0(N__53234),
            .in1(N__58265),
            .in2(N__53360),
            .in3(N__51402),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.state_3_LC_7_15_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_7_15_7 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_7_15_7  (
            .in0(N__51407),
            .in1(N__53355),
            .in2(N__58301),
            .in3(N__39861),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83980),
            .ce(),
            .sr(N__77284));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_7_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65211),
            .lcout(drone_H_disp_front_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83996),
            .ce(N__38624),
            .sr(N__77293));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_7_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57991),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83996),
            .ce(N__38624),
            .sr(N__77293));
    defparam \dron_frame_decoder_1.state_RNITC181_3_LC_7_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNITC181_3_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNITC181_3_LC_7_17_1 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \dron_frame_decoder_1.state_RNITC181_3_LC_7_17_1  (
            .in0(N__58312),
            .in1(N__53359),
            .in2(N__53265),
            .in3(N__77621),
            .lcout(\dron_frame_decoder_1.N_371_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_17_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__40241),
            .in2(_gnd_net_),
            .in3(N__77622),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_17_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_17_5  (
            .in0(N__58311),
            .in1(N__58401),
            .in2(N__38601),
            .in3(N__38577),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIM14N_0_LC_7_17_7 .C_ON=1'b0;
    defparam \pid_front.state_RNIM14N_0_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIM14N_0_LC_7_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.state_RNIM14N_0_LC_7_17_7  (
            .in0(N__46076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83003),
            .lcout(\pid_front.state_RNIM14NZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_7_18_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_7_18_0 .LUT_INIT=16'b1101000011111101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6B6F_6_LC_7_18_0  (
            .in0(N__40320),
            .in1(N__40291),
            .in2(N__38664),
            .in3(N__38670),
            .lcout(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_7_18_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_7_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__39962),
            .in2(_gnd_net_),
            .in3(N__39894),
            .lcout(\pid_front.N_1662_i ),
            .ltout(\pid_front.N_1662_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_7_18_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_7_18_2 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_7_18_2  (
            .in0(N__38660),
            .in1(N__40317),
            .in2(N__38643),
            .in3(N__40290),
            .lcout(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ),
            .ltout(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_7_18_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_7_18_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_7_18_3  (
            .in0(N__43811),
            .in1(_gnd_net_),
            .in2(N__38640),
            .in3(N__40038),
            .lcout(\pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_7_18_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_7_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIU9ST_6_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__43810),
            .in2(_gnd_net_),
            .in3(N__38637),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIHMAE2_5_LC_7_18_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIHMAE2_5_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIHMAE2_5_LC_7_18_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIHMAE2_5_LC_7_18_5  (
            .in0(N__40140),
            .in1(N__40037),
            .in2(N__38631),
            .in3(N__43855),
            .lcout(\pid_front.error_p_reg_esr_RNIHMAE2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_6_LC_7_18_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_7_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_6_LC_7_18_6  (
            .in0(N__39895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84029),
            .ce(N__52541),
            .sr(N__52428));
    defparam \pid_front.error_d_reg_prev_esr_5_LC_7_18_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_7_18_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_5_LC_7_18_7  (
            .in0(N__40292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84029),
            .ce(N__52541),
            .sr(N__52428));
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_7_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_7_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_13_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48054),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_7_19_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_12_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51925),
            .lcout(\pid_front.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_7_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_11_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51891),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_7_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_7_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_2_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49358),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_7_19_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_7_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_4_LC_7_19_4  (
            .in0(N__43887),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_7_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_7_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_5_LC_7_19_5  (
            .in0(N__43857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_7_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_6_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43815),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_7_19_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_7_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_7_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43782),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84045),
            .ce(N__46063),
            .sr(N__77319));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_7_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80467),
            .lcout(front_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_7_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73787),
            .lcout(front_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_7_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_7_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_7_20_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_7_20_2  (
            .in0(N__80262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(front_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_7_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_7_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79714),
            .lcout(front_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_7_20_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80105),
            .lcout(front_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_7_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_7_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81086),
            .lcout(front_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_7_20_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_7_20_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_7_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79891),
            .lcout(front_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84061),
            .ce(N__40448),
            .sr(N__77326));
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_7_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_7_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_8_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43746),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84078),
            .ce(N__46059),
            .sr(N__77333));
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_7_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_7_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_9_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47766),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84078),
            .ce(N__46059),
            .sr(N__77333));
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_7_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_7_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_10_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47919),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84078),
            .ce(N__46059),
            .sr(N__77333));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_7_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_7_22_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41694),
            .in3(N__41812),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_7_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_7_22_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_7_22_6  (
            .in0(N__41813),
            .in1(N__41689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_7_23_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_7_23_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_7_23_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__80463),
            .in2(_gnd_net_),
            .in3(N__83014),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84097),
            .ce(N__38750),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_7_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_7_23_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__80104),
            .in2(_gnd_net_),
            .in3(N__83013),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84097),
            .ce(N__38750),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_3_LC_7_23_7 .C_ON=1'b0;
    defparam \pid_side.error_axb_3_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_3_LC_7_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_3_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40463),
            .lcout(\pid_side.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_7_24_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_7_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49723),
            .lcout(drone_H_disp_front_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_8_4_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_8_4_7 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_8_4_7  (
            .in0(N__42432),
            .in1(N__42393),
            .in2(N__48347),
            .in3(N__38697),
            .lcout(\Commands_frame_decoder.N_364_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_5_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state57_i_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__48332),
            .in2(_gnd_net_),
            .in3(N__77630),
            .lcout(\Commands_frame_decoder.un1_state57_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_8_5_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_8_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_4_LC_8_5_3  (
            .in0(N__42170),
            .in1(N__42152),
            .in2(N__42135),
            .in3(N__42110),
            .lcout(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_8_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_8_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIHV6P_11_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__42490),
            .in2(_gnd_net_),
            .in3(N__42469),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_8_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_8_6_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_8_6_1  (
            .in0(N__38850),
            .in1(N__38706),
            .in2(N__38700),
            .in3(N__38856),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(\Commands_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_8_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_8_6_2 .LUT_INIT=16'b0001000100010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_8_6_2  (
            .in0(N__48331),
            .in1(N__42427),
            .in2(N__38688),
            .in3(N__42390),
            .lcout(\Commands_frame_decoder.N_402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_8_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_8_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNITK4L_8_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__42556),
            .in2(_gnd_net_),
            .in3(N__42604),
            .lcout(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_6 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_6  (
            .in0(N__42512),
            .in1(N__42491),
            .in2(N__42581),
            .in3(N__42470),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_8_7_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_8_7_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_8_7_0  (
            .in0(N__38829),
            .in1(N__38843),
            .in2(N__38832),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_8_7_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_8_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__40637),
            .in2(_gnd_net_),
            .in3(N__38811),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_8_7_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__42995),
            .in2(_gnd_net_),
            .in3(N__38808),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_8_7_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_8_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__42951),
            .in2(_gnd_net_),
            .in3(N__38805),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_8_7_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_8_7_4 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_2_LC_8_7_4  (
            .in0(N__38802),
            .in1(N__42348),
            .in2(N__77666),
            .in3(N__42318),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83867),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_8_7_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_8_7_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_8_7_5  (
            .in0(N__40831),
            .in1(N__40875),
            .in2(N__41070),
            .in3(N__40752),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_8_7_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_8_7_7 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart_drone.timer_Count_4_LC_8_7_7  (
            .in0(N__42319),
            .in1(N__77642),
            .in2(N__42354),
            .in3(N__38796),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83867),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_8_8_0 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_8_8_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \uart_pc.data_4_LC_8_8_0  (
            .in0(N__39041),
            .in1(N__39197),
            .in2(N__39612),
            .in3(N__79197),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83877),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI53692_14_LC_8_8_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI53692_14_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI53692_14_LC_8_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI53692_14_LC_8_8_2  (
            .in0(N__42669),
            .in1(N__40857),
            .in2(N__40911),
            .in3(N__39843),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_12_LC_8_8_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_8_8_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_12_LC_8_8_3  (
            .in0(N__40944),
            .in1(N__40809),
            .in2(N__39021),
            .in3(N__38958),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_8_8_4 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_8_8_4 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_8_8_4  (
            .in0(N__40810),
            .in1(N__40671),
            .in2(N__39018),
            .in3(N__39010),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83877),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_8_8_6 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_8_8_6 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \reset_module_System.count_2_LC_8_8_6  (
            .in0(N__40776),
            .in1(N__40672),
            .in2(N__39014),
            .in3(N__38977),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83877),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_8_8_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_8_8_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_8_8_7  (
            .in0(N__40733),
            .in1(N__40766),
            .in2(N__41028),
            .in3(N__40787),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_8_9_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_8_9_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_8_9_0  (
            .in0(N__38949),
            .in1(N__38904),
            .in2(_gnd_net_),
            .in3(N__77620),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_8_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_8_9_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_1_4_LC_8_9_1  (
            .in0(N__39201),
            .in1(N__39168),
            .in2(N__39057),
            .in3(N__80037),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83888),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_9_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_8_9_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_8_9_2  (
            .in0(N__39543),
            .in1(N__39587),
            .in2(_gnd_net_),
            .in3(N__39495),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_9_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_8_9_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_8_9_3  (
            .in0(N__39494),
            .in1(N__39590),
            .in2(_gnd_net_),
            .in3(N__39542),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_8_9_4 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_8_9_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_5_LC_8_9_4  (
            .in0(N__39170),
            .in1(N__39203),
            .in2(N__39441),
            .in3(N__81010),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83888),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_8_9_6 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_8_9_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_LC_8_9_6  (
            .in0(N__39169),
            .in1(N__39202),
            .in2(N__39120),
            .in3(N__73662),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83888),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_8_9_7 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_8_9_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_6_LC_8_9_7  (
            .in0(N__39204),
            .in1(N__39171),
            .in2(N__39258),
            .in3(N__79857),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83888),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_8_10_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_8_10_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uart_pc.data_Aux_0_LC_8_10_0  (
            .in0(N__39137),
            .in1(N__39147),
            .in2(N__39423),
            .in3(N__39311),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_1_LC_8_10_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_8_10_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_1_LC_8_10_1  (
            .in0(N__39312),
            .in1(N__39113),
            .in2(N__39421),
            .in3(N__39126),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_2_LC_8_10_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_8_10_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_8_10_2  (
            .in0(N__39102),
            .in1(N__39408),
            .in2(N__39095),
            .in3(N__39313),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_3_LC_8_10_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_8_10_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_3_LC_8_10_3  (
            .in0(N__39314),
            .in1(N__39071),
            .in2(N__39422),
            .in3(N__39078),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_8_10_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_8_10_4  (
            .in0(N__39493),
            .in1(_gnd_net_),
            .in2(N__39546),
            .in3(N__39589),
            .lcout(),
            .ltout(\uart_pc.data_Auxce_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_5_LC_8_10_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_8_10_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uart_pc.data_Aux_5_LC_8_10_5  (
            .in0(N__39316),
            .in1(N__39419),
            .in2(N__39060),
            .in3(N__39053),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_4_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_8_10_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_8_10_6  (
            .in0(N__39618),
            .in1(N__39409),
            .in2(N__39608),
            .in3(N__39315),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83899),
            .ce(),
            .sr(N__39236));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_8_10_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_8_10_7  (
            .in0(N__39588),
            .in1(N__39538),
            .in2(_gnd_net_),
            .in3(N__39492),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_6_LC_8_11_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_8_11_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \uart_pc.data_Aux_6_LC_8_11_0  (
            .in0(N__39317),
            .in1(N__39434),
            .in2(N__39450),
            .in3(N__39407),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83913),
            .ce(),
            .sr(N__39237));
    defparam \uart_pc.data_Aux_7_LC_8_11_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_8_11_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \uart_pc.data_Aux_7_LC_8_11_1  (
            .in0(N__39406),
            .in1(N__39318),
            .in2(N__39254),
            .in3(N__39282),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83913),
            .ce(),
            .sr(N__39237));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_8_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_8_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__48247),
            .in2(_gnd_net_),
            .in3(N__39218),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_8_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_8_11_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_8_11_5  (
            .in0(N__48248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40155),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_8_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_8_11_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39207),
            .in3(N__77608),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_12_LC_8_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_8_12_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_12_LC_8_12_1  (
            .in0(N__48276),
            .in1(N__48365),
            .in2(N__39723),
            .in3(N__40205),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_11_LC_8_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_8_12_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_8_12_2  (
            .in0(N__40204),
            .in1(N__39705),
            .in2(N__48346),
            .in3(N__39722),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_8_12_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_10_LC_8_12_3  (
            .in0(N__39704),
            .in1(N__44609),
            .in2(_gnd_net_),
            .in3(N__40203),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_8_LC_8_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_8_12_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_8_12_4  (
            .in0(N__40208),
            .in1(N__48278),
            .in2(N__41192),
            .in3(N__39689),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_9_LC_8_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_8_12_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_9_LC_8_12_5  (
            .in0(N__48277),
            .in1(N__41205),
            .in2(N__39690),
            .in3(N__40209),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_7_LC_8_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_8_12_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_8_12_6  (
            .in0(N__40207),
            .in1(N__41188),
            .in2(N__39665),
            .in3(N__48279),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \Commands_frame_decoder.state_6_LC_8_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_8_12_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_6_LC_8_12_7  (
            .in0(N__39661),
            .in1(N__39678),
            .in2(_gnd_net_),
            .in3(N__40206),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83923),
            .ce(),
            .sr(N__77273));
    defparam \dron_frame_decoder_1.WDT_RNISF2A1_10_LC_8_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNISF2A1_10_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNISF2A1_10_LC_8_13_0 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNISF2A1_10_LC_8_13_0  (
            .in0(N__39774),
            .in1(N__41299),
            .in2(N__41343),
            .in3(N__41321),
            .lcout(\dron_frame_decoder_1.WDT10lt13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIBAK71_10_LC_8_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIBAK71_10_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIBAK71_10_LC_8_13_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIBAK71_10_LC_8_13_1  (
            .in0(N__41320),
            .in1(_gnd_net_),
            .in2(N__41301),
            .in3(N__41338),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10_0_icf0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIVT8F2_15_LC_8_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIVT8F2_15_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIVT8F2_15_LC_8_13_2 .LUT_INIT=16'b0101010111110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIVT8F2_15_LC_8_13_2  (
            .in0(N__41428),
            .in1(N__41272),
            .in2(N__39624),
            .in3(N__41227),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10_0_icf0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIN9PJ4_15_LC_8_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIN9PJ4_15_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIN9PJ4_15_LC_8_13_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIN9PJ4_15_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__39783),
            .in2(N__39621),
            .in3(N__39773),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIJIDQ_11_LC_8_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIJIDQ_11_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIJIDQ_11_LC_8_13_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIJIDQ_11_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__41295),
            .in2(_gnd_net_),
            .in3(N__41319),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10_0_icf1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI76222_15_LC_8_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI76222_15_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI76222_15_LC_8_13_5 .LUT_INIT=16'b0111001101110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI76222_15_LC_8_13_5  (
            .in0(N__41226),
            .in1(N__41427),
            .in2(N__39786),
            .in3(N__41254),
            .lcout(\dron_frame_decoder_1.WDT10_0_icf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIB571_5_LC_8_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIB571_5_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIB571_5_LC_8_13_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIB571_5_LC_8_13_6  (
            .in0(N__41357),
            .in1(N__41372),
            .in2(_gnd_net_),
            .in3(N__41099),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10lto9_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIH5E2_4_LC_8_13_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIH5E2_4_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIH5E2_4_LC_8_13_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIH5E2_4_LC_8_13_7  (
            .in0(N__41387),
            .in1(N__41084),
            .in2(N__39777),
            .in3(N__41114),
            .lcout(\dron_frame_decoder_1.WDT10lt10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_3_1_LC_8_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_3_1_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_3_1_LC_8_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_3_1_LC_8_14_0  (
            .in0(N__64966),
            .in1(N__65201),
            .in2(N__58280),
            .in3(N__57979),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIMEKA3_1_LC_8_14_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIMEKA3_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIMEKA3_1_LC_8_14_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIMEKA3_1_LC_8_14_1  (
            .in0(N__64967),
            .in1(N__39765),
            .in2(N__51381),
            .in3(N__39759),
            .lcout(\dron_frame_decoder_1.N_127_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.m34_2_LC_8_14_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.m34_2_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.m34_2_LC_8_14_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \dron_frame_decoder_1.m34_2_LC_8_14_2  (
            .in0(N__68542),
            .in1(N__65200),
            .in2(_gnd_net_),
            .in3(N__57978),
            .lcout(\dron_frame_decoder_1.m34Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.m15_LC_8_14_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.m15_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.m15_LC_8_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.m15_LC_8_14_3  (
            .in0(N__68632),
            .in1(N__71798),
            .in2(N__65126),
            .in3(N__72025),
            .lcout(\dron_frame_decoder_1.N_123_mux ),
            .ltout(\dron_frame_decoder_1.N_123_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIUS6K3_0_LC_8_14_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIUS6K3_0_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIUS6K3_0_LC_8_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIUS6K3_0_LC_8_14_4  (
            .in0(N__68543),
            .in1(N__39751),
            .in2(N__39732),
            .in3(N__39729),
            .lcout(\dron_frame_decoder_1.N_186 ),
            .ltout(\dron_frame_decoder_1.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_8_14_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_8_14_5 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_8_14_5  (
            .in0(N__51379),
            .in1(N__39879),
            .in2(N__39864),
            .in3(N__39860),
            .lcout(\dron_frame_decoder_1.state_ns_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_rdy_LC_8_14_7 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_8_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.data_rdy_LC_8_14_7  (
            .in0(N__43179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42630),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83950),
            .ce(),
            .sr(N__77285));
    defparam \pid_side.state_RNINK4U_0_0_LC_8_15_0 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_0_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_0_LC_8_15_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNINK4U_0_0_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__67218),
            .in2(_gnd_net_),
            .in3(N__77602),
            .lcout(\pid_side.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_15_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__40965),
            .in2(_gnd_net_),
            .in3(N__40986),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_15_3 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_8_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79870),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83964),
            .ce(N__42891),
            .sr(N__77294));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_4 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__47421),
            .in2(_gnd_net_),
            .in3(N__44588),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_8_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_8_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39834),
            .lcout(drone_H_disp_front_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_8_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_8_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39828),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_8_16_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_8_16_0 .LUT_INIT=16'b0101100110100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_8_16_0  (
            .in0(N__41475),
            .in1(N__41594),
            .in2(N__41619),
            .in3(N__41481),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ),
            .ltout(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_8_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIS0F23_7_LC_8_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIS0F23_7_LC_8_16_1  (
            .in0(N__45272),
            .in1(N__39947),
            .in2(N__40029),
            .in3(N__43744),
            .lcout(\pid_front.error_p_reg_esr_RNIS0F23Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_8_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_8_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3K9L1_6_LC_8_16_2  (
            .in0(N__43781),
            .in1(_gnd_net_),
            .in2(N__40014),
            .in3(N__40020),
            .lcout(\pid_front.error_p_reg_esr_RNI3K9L1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_8_16_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_8_16_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_8_16_3  (
            .in0(N__40026),
            .in1(N__39948),
            .in2(_gnd_net_),
            .in3(N__43745),
            .lcout(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_8_16_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_8_16_4 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_8_16_4  (
            .in0(N__39897),
            .in1(N__39990),
            .in2(N__39972),
            .in3(N__39996),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ),
            .ltout(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_8_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_8_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3K9L1_0_6_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__40010),
            .in2(N__39999),
            .in3(N__43780),
            .lcout(\pid_front.error_p_reg_esr_RNI3K9L1_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_8_16_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_8_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__41593),
            .in2(_gnd_net_),
            .in3(N__41613),
            .lcout(\pid_front.N_1668_i ),
            .ltout(\pid_front.N_1668_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_8_16_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_8_16_7 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_7_LC_8_16_7  (
            .in0(N__39989),
            .in1(N__39968),
            .in2(N__39951),
            .in3(N__39896),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_5_LC_8_17_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_5_LC_8_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_5_LC_8_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_5_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39939),
            .lcout(\pid_front.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83997),
            .ce(N__83090),
            .sr(N__82877));
    defparam \pid_front.error_d_reg_esr_6_LC_8_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_6_LC_8_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_6_LC_8_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_6_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39915),
            .lcout(\pid_front.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83997),
            .ce(N__83090),
            .sr(N__82877));
    defparam \pid_front.error_d_reg_esr_7_LC_8_17_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_7_LC_8_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_7_LC_8_17_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_7_LC_8_17_2  (
            .in0(N__40125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83997),
            .ce(N__83090),
            .sr(N__82877));
    defparam \pid_front.error_p_reg_esr_10_LC_8_17_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_10_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_10_LC_8_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_10_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40110),
            .lcout(\pid_front.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83997),
            .ce(N__83090),
            .sr(N__82877));
    defparam \pid_front.error_p_reg_esr_11_LC_8_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_11_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_11_LC_8_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_11_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40095),
            .lcout(\pid_front.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83997),
            .ce(N__83090),
            .sr(N__82877));
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_8_18_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_8_18_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIMI772_3_LC_8_18_0  (
            .in0(N__40080),
            .in1(N__47454),
            .in2(N__45458),
            .in3(N__43883),
            .lcout(\pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_8_18_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_8_18_1 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_8_18_1  (
            .in0(N__40050),
            .in1(N__75860),
            .in2(N__40071),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ),
            .ltout(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI4U472_3_LC_8_18_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI4U472_3_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI4U472_3_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI4U472_3_LC_8_18_2  (
            .in0(N__47532),
            .in1(N__47453),
            .in2(N__40074),
            .in3(N__43882),
            .lcout(\pid_front.error_p_reg_esr_RNI4U472Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_4_LC_8_18_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_8_18_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_4_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__75861),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84015),
            .ce(N__52527),
            .sr(N__52429));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_8_18_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_8_18_4 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_4_LC_8_18_4  (
            .in0(N__75859),
            .in1(N__40067),
            .in2(_gnd_net_),
            .in3(N__40049),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ),
            .ltout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_8_18_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_8_18_5 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_5_LC_8_18_5  (
            .in0(N__40299),
            .in1(N__40274),
            .in2(N__40041),
            .in3(N__40319),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_8_18_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_8_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_8_18_6  (
            .in0(N__40318),
            .in1(N__40298),
            .in2(N__40275),
            .in3(N__40254),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ),
            .ltout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKJHV_0_5_LC_8_18_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKJHV_0_5_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKJHV_0_5_LC_8_18_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKJHV_0_5_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40248),
            .in3(N__43848),
            .lcout(\pid_front.error_p_reg_esr_RNIKJHV_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_5_LC_8_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_8_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_8_19_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_5_LC_8_19_0  (
            .in0(N__40154),
            .in1(N__40245),
            .in2(_gnd_net_),
            .in3(N__40224),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84030),
            .ce(),
            .sr(N__77327));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_8_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_8_19_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__51618),
            .in2(_gnd_net_),
            .in3(N__78749),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIUO6U_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIFM151_0_LC_8_19_4 .C_ON=1'b0;
    defparam \pid_front.state_RNIFM151_0_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIFM151_0_LC_8_19_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNIFM151_0_LC_8_19_4  (
            .in0(N__52378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46077),
            .lcout(\pid_front.N_404_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKJHV_5_LC_8_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKJHV_5_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKJHV_5_LC_8_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKJHV_5_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__40139),
            .in2(_gnd_net_),
            .in3(N__43856),
            .lcout(\pid_front.error_p_reg_esr_RNIKJHVZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNISV141_0_LC_8_19_6 .C_ON=1'b0;
    defparam \pid_front.state_RNISV141_0_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNISV141_0_LC_8_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNISV141_0_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__52047),
            .in2(_gnd_net_),
            .in3(N__83005),
            .lcout(\pid_front.N_429_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_8_20_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_8_20_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_8_20_0  (
            .in0(N__41747),
            .in1(N__42083),
            .in2(N__41732),
            .in3(N__51725),
            .lcout(\pid_front.un10lt9_1 ),
            .ltout(\pid_front.un10lt9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_8_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_8_20_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_8_20_1  (
            .in0(N__41893),
            .in1(N__41644),
            .in2(N__40128),
            .in3(N__41666),
            .lcout(),
            .ltout(\pid_front.error_i_acumm16lt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_8_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_8_20_2 .LUT_INIT=16'b0100010001001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_8_20_2  (
            .in0(N__40362),
            .in1(N__42272),
            .in2(N__40353),
            .in3(N__40341),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_8_20_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_8_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_8_20_3  (
            .in0(N__41645),
            .in1(N__41665),
            .in2(N__41897),
            .in3(N__40350),
            .lcout(),
            .ltout(\pid_front.un10lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_8_20_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_8_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_8_20_4  (
            .in0(N__41573),
            .in1(N__41764),
            .in2(N__40344),
            .in3(N__41552),
            .lcout(\pid_front.un10lt11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_8_20_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_8_20_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_8_20_5  (
            .in0(N__41765),
            .in1(N__41551),
            .in2(_gnd_net_),
            .in3(N__41572),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_8_20_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_8_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_8_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_3_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47559),
            .lcout(\pid_front.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84046),
            .ce(N__46064),
            .sr(N__77334));
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_8_20_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_8_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_8_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_1_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52273),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84046),
            .ce(N__46064),
            .sr(N__77334));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_8_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_8_21_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_8_21_0  (
            .in0(N__42033),
            .in1(N__41990),
            .in2(N__42015),
            .in3(N__42024),
            .lcout(\pid_front.error_i_acumm16lto27_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_8_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_8_21_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_8_21_1  (
            .in0(N__41870),
            .in1(_gnd_net_),
            .in2(N__44196),
            .in3(N__40410),
            .lcout(),
            .ltout(\pid_front.error_i_acumm16lto27_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_8_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_8_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_8_21_2  (
            .in0(N__40422),
            .in1(N__40326),
            .in2(N__40335),
            .in3(N__40332),
            .lcout(\pid_front.error_i_acumm16lto27_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_8_21_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_8_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_8_21_3  (
            .in0(N__40487),
            .in1(N__40374),
            .in2(N__42066),
            .in3(N__40385),
            .lcout(\pid_front.error_i_acumm16lto27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_8_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_8_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_8_21_4  (
            .in0(N__42003),
            .in1(N__40476),
            .in2(N__42048),
            .in3(N__40505),
            .lcout(\pid_front.error_i_acumm16lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_8_21_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_8_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_8_21_5  (
            .in0(N__42023),
            .in1(N__42011),
            .in2(N__41991),
            .in3(N__42032),
            .lcout(),
            .ltout(\pid_front.un10lto27_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_8_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_8_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_8_21_6  (
            .in0(N__40409),
            .in1(N__41869),
            .in2(N__40413),
            .in3(N__44192),
            .lcout(\pid_front.un10lto27_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_8_21_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_8_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_8_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_26_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48657),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84062),
            .ce(N__46061),
            .sr(N__77341));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_8_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_8_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_8_22_0  (
            .in0(N__40491),
            .in1(N__40373),
            .in2(N__42065),
            .in3(N__40386),
            .lcout(),
            .ltout(\pid_front.un10lto27_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_8_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_8_22_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__40392),
            .in2(N__40401),
            .in3(N__40398),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_8_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_8_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_8_22_2  (
            .in0(N__42002),
            .in1(N__40475),
            .in2(N__40506),
            .in3(N__42044),
            .lcout(\pid_front.un10lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_8_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_8_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_8_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_18_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49059),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84079),
            .ce(N__46060),
            .sr(N__77345));
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_8_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_8_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_8_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_19_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48966),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84079),
            .ce(N__46060),
            .sr(N__77345));
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_8_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_8_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_8_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_14_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43962),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84079),
            .ce(N__46060),
            .sr(N__77345));
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_8_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_8_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_8_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_20_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46338),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84079),
            .ce(N__46060),
            .sr(N__77345));
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_8_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_8_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_8_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_15_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48456),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84079),
            .ce(N__46060),
            .sr(N__77345));
    defparam \dron_frame_decoder_1.source_H_disp_front_1_LC_8_23_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_1_LC_8_23_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_1_LC_8_23_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_1_LC_8_23_1  (
            .in0(N__58338),
            .in1(N__58004),
            .in2(N__53326),
            .in3(N__42222),
            .lcout(drone_H_disp_front_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84089),
            .ce(),
            .sr(N__77349));
    defparam \dron_frame_decoder_1.source_H_disp_front_3_LC_8_23_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_3_LC_8_23_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_3_LC_8_23_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_3_LC_8_23_3  (
            .in0(N__58339),
            .in1(N__64994),
            .in2(N__53327),
            .in3(N__42210),
            .lcout(drone_H_disp_front_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84089),
            .ce(),
            .sr(N__77349));
    defparam \dron_frame_decoder_1.source_H_disp_front_4_LC_8_23_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_4_LC_8_23_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_4_LC_8_23_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_4_LC_8_23_5  (
            .in0(N__58340),
            .in1(N__65235),
            .in2(N__53328),
            .in3(N__41979),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84089),
            .ce(),
            .sr(N__77349));
    defparam \dron_frame_decoder_1.source_H_disp_side_3_LC_8_23_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_3_LC_8_23_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_3_LC_8_23_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_3_LC_8_23_7  (
            .in0(N__58341),
            .in1(N__64995),
            .in2(N__71956),
            .in3(N__40464),
            .lcout(drone_H_disp_side_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84089),
            .ce(),
            .sr(N__77349));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_8_24_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_8_24_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_8_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_8_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79289),
            .lcout(front_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84098),
            .ce(N__40452),
            .sr(N__77354));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_3_1 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_3_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_3_1  (
            .in0(N__40431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83827),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40581),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83827),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_9_4_0 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_9_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40548),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83832),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_9_4_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_9_4_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_9_4_5  (
            .in0(N__40566),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83832),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_9_4_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40554),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83832),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__40542),
            .in2(N__42530),
            .in3(N__42531),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__40536),
            .in2(_gnd_net_),
            .in3(N__40530),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__40527),
            .in2(_gnd_net_),
            .in3(N__40521),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__40518),
            .in2(_gnd_net_),
            .in3(N__40512),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__42111),
            .in2(_gnd_net_),
            .in3(N__40509),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__42153),
            .in2(_gnd_net_),
            .in3(N__40608),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__42171),
            .in2(_gnd_net_),
            .in3(N__40605),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__42133),
            .in2(_gnd_net_),
            .in3(N__40602),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__83840),
            .ce(),
            .sr(N__40703));
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__42606),
            .in2(_gnd_net_),
            .in3(N__40599),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__42558),
            .in2(_gnd_net_),
            .in3(N__40596),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__42580),
            .in2(_gnd_net_),
            .in3(N__40593),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__42471),
            .in2(_gnd_net_),
            .in3(N__40590),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__42492),
            .in2(_gnd_net_),
            .in3(N__40587),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__42513),
            .in2(_gnd_net_),
            .in3(N__40584),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__42391),
            .in2(_gnd_net_),
            .in3(N__40710),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__42428),
            .in2(_gnd_net_),
            .in3(N__40707),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83849),
            .ce(),
            .sr(N__40704));
    defparam \uart_drone.state_RNO_0_3_LC_9_7_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_9_7_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_9_7_0  (
            .in0(N__42989),
            .in1(N__42932),
            .in2(N__43064),
            .in3(N__42731),
            .lcout(\uart_drone.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_9_7_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__40811),
            .in2(_gnd_net_),
            .in3(N__40838),
            .lcout(\reset_module_System.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_9_7_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_9_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_9_7_3  (
            .in0(N__40893),
            .in1(N__41046),
            .in2(N__41004),
            .in3(N__40929),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_7_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_9_7_4 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_9_7_4  (
            .in0(N__42987),
            .in1(N__42826),
            .in2(N__40638),
            .in3(N__42930),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__40636),
            .in2(_gnd_net_),
            .in3(N__42988),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_9_7_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_9_7_6  (
            .in0(N__42830),
            .in1(N__42931),
            .in2(N__40620),
            .in3(N__77623),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_9_7_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_9_7_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_9_7_7  (
            .in0(N__77624),
            .in1(N__42307),
            .in2(N__40617),
            .in3(N__40614),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83858),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_9_8_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__40839),
            .in2(N__40812),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_9_8_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_9_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__40788),
            .in2(_gnd_net_),
            .in3(N__40770),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_9_8_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_9_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__40767),
            .in2(_gnd_net_),
            .in3(N__40755),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_9_8_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_9_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__40751),
            .in2(_gnd_net_),
            .in3(N__40740),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_9_8_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_9_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__42681),
            .in2(_gnd_net_),
            .in3(N__40737),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_9_8_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_9_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__40734),
            .in2(_gnd_net_),
            .in3(N__40722),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_9_8_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_9_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__42708),
            .in2(_gnd_net_),
            .in3(N__40719),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_9_8_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_9_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__42720),
            .in2(_gnd_net_),
            .in3(N__40716),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__83868),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_9_9_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_9_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__42695),
            .in2(_gnd_net_),
            .in3(N__40713),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_9_9_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_9_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__40982),
            .in2(_gnd_net_),
            .in3(N__40968),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_9_9_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_9_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__40961),
            .in2(_gnd_net_),
            .in3(N__40947),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_9_9_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_9_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__40943),
            .in2(_gnd_net_),
            .in3(N__40932),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_9_9_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_9_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__40925),
            .in2(_gnd_net_),
            .in3(N__40914),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_9_9_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_9_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__40910),
            .in2(_gnd_net_),
            .in3(N__40896),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_9_9_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_9_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__40889),
            .in2(_gnd_net_),
            .in3(N__40878),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_9_9_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_9_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__40871),
            .in2(_gnd_net_),
            .in3(N__40860),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__83878),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_9_10_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_9_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__40856),
            .in2(_gnd_net_),
            .in3(N__40842),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__83889),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_9_10_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_9_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__41063),
            .in2(_gnd_net_),
            .in3(N__41049),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__83889),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_9_10_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_9_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__41045),
            .in2(_gnd_net_),
            .in3(N__41031),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__83889),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_9_10_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_9_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__41024),
            .in2(_gnd_net_),
            .in3(N__41010),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__83889),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_9_10_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_9_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__41000),
            .in2(_gnd_net_),
            .in3(N__41007),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83889),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_11_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_9_11_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_9_11_1  (
            .in0(N__44904),
            .in1(_gnd_net_),
            .in2(N__44855),
            .in3(N__44793),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_11_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_9_11_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_9_11_4  (
            .in0(N__44794),
            .in1(N__44841),
            .in2(_gnd_net_),
            .in3(N__44905),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_9_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_9_11_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_9_11_5  (
            .in0(N__44906),
            .in1(_gnd_net_),
            .in2(N__44856),
            .in3(N__44795),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_9_11_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_9_11_7  (
            .in0(N__44907),
            .in1(_gnd_net_),
            .in2(N__44857),
            .in3(N__44796),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_12_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_9_12_0 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_9_12_0  (
            .in0(N__44797),
            .in1(_gnd_net_),
            .in2(N__44858),
            .in3(N__44913),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_9_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_9_12_2  (
            .in0(N__41204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48320),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_9_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_9_12_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_9_12_6  (
            .in0(N__41184),
            .in1(N__48321),
            .in2(_gnd_net_),
            .in3(N__77631),
            .lcout(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_9_13_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_9_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__41148),
            .in2(N__41163),
            .in3(N__41162),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_1_LC_9_13_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__41142),
            .in2(_gnd_net_),
            .in3(N__41136),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_2_LC_9_13_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_9_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__41133),
            .in2(_gnd_net_),
            .in3(N__41127),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_3_LC_9_13_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__41124),
            .in2(_gnd_net_),
            .in3(N__41118),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_4_LC_9_13_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__41115),
            .in2(_gnd_net_),
            .in3(N__41103),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_5_LC_9_13_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_9_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__41100),
            .in2(_gnd_net_),
            .in3(N__41088),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_6_LC_9_13_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__41085),
            .in2(_gnd_net_),
            .in3(N__41073),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_7_LC_9_13_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__41388),
            .in2(_gnd_net_),
            .in3(N__41376),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__83924),
            .ce(),
            .sr(N__58551));
    defparam \dron_frame_decoder_1.WDT_8_LC_9_14_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__41373),
            .in2(_gnd_net_),
            .in3(N__41361),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_9_LC_9_14_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__41358),
            .in2(_gnd_net_),
            .in3(N__41346),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_10_LC_9_14_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__41342),
            .in2(_gnd_net_),
            .in3(N__41325),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_11_LC_9_14_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__41322),
            .in2(_gnd_net_),
            .in3(N__41304),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_12_LC_9_14_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__41300),
            .in2(_gnd_net_),
            .in3(N__41280),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_13_LC_9_14_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__41276),
            .in2(_gnd_net_),
            .in3(N__41238),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_14_LC_9_14_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__41231),
            .in2(_gnd_net_),
            .in3(N__41208),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \dron_frame_decoder_1.WDT_15_LC_9_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_9_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__41432),
            .in2(_gnd_net_),
            .in3(N__41442),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83937),
            .ce(),
            .sr(N__58550));
    defparam \pid_front.pid_prereg_14_LC_9_15_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_14_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_14_LC_9_15_0 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_front.pid_prereg_14_LC_9_15_0  (
            .in0(N__41409),
            .in1(N__45651),
            .in2(N__52184),
            .in3(N__45639),
            .lcout(\pid_front.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83951),
            .ce(),
            .sr(N__77303));
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_9_15_1 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_9_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_RNO_LC_9_15_1  (
            .in0(N__41407),
            .in1(N__45692),
            .in2(N__45624),
            .in3(N__45743),
            .lcout(\pid_front.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_4_c_RNO_LC_9_15_2 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_4_c_RNO_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_4_c_RNO_LC_9_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_4_c_RNO_LC_9_15_2  (
            .in0(N__45578),
            .in1(N__45545),
            .in2(N__45945),
            .in3(N__45602),
            .lcout(\pid_front.un11lto30_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIQ6EV_17_LC_9_15_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIQ6EV_17_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIQ6EV_17_LC_9_15_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIQ6EV_17_LC_9_15_3  (
            .in0(N__45546),
            .in1(N__45944),
            .in2(_gnd_net_),
            .in3(N__45579),
            .lcout(),
            .ltout(\pid_front.pid_prereg_esr_RNIQ6EVZ0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_9_15_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_9_15_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI295P1_15_LC_9_15_4  (
            .in0(N__41408),
            .in1(N__45603),
            .in2(N__41394),
            .in3(N__45623),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ),
            .ltout(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_9_15_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_9_15_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIUHO16_12_LC_9_15_5  (
            .in0(N__45744),
            .in1(N__45693),
            .in2(N__41391),
            .in3(N__43470),
            .lcout(\pid_front.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_0_LC_9_15_7 .C_ON=1'b0;
    defparam \pid_front.state_0_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_0_LC_9_15_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_0_LC_9_15_7  (
            .in0(N__52110),
            .in1(N__67377),
            .in2(_gnd_net_),
            .in3(N__52169),
            .lcout(\pid_front.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83951),
            .ce(),
            .sr(N__77303));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_9_16_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_9_16_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_9_16_0  (
            .in0(N__84133),
            .in1(N__41504),
            .in2(_gnd_net_),
            .in3(N__41489),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_9_16_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_9_16_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_9_16_1  (
            .in0(N__51610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78766),
            .lcout(\pid_front.N_1698_i ),
            .ltout(\pid_front.N_1698_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_9_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_9_16_2 .LUT_INIT=16'b1010111110001110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIROQ33_12_LC_9_16_2  (
            .in0(N__43559),
            .in1(N__43595),
            .in2(N__41529),
            .in3(N__43618),
            .lcout(\pid_front.error_p_reg_esr_RNIROQ33Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_9_16_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_9_16_3 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVTNC2_13_LC_9_16_3  (
            .in0(N__48837),
            .in1(N__78697),
            .in2(N__48878),
            .in3(N__47960),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIVTNC2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_9_16_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_9_16_4 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_9_16_4  (
            .in0(N__48005),
            .in1(N__41526),
            .in2(N__41514),
            .in3(N__41511),
            .lcout(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_14_LC_9_16_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_9_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_14_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84135),
            .lcout(\pid_front.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83965),
            .ce(N__52542),
            .sr(N__52448));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_16_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_16_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_16_6  (
            .in0(N__84134),
            .in1(N__41505),
            .in2(_gnd_net_),
            .in3(N__41490),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_9_16_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_9_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_9_16_7  (
            .in0(N__48836),
            .in1(N__48871),
            .in2(_gnd_net_),
            .in3(N__78696),
            .lcout(\pid_front.error_p_reg_esr_RNIETB61_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_17_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_9_17_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_8_LC_9_17_0  (
            .in0(N__82298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83981),
            .ce(N__52540),
            .sr(N__52444));
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_9_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_9_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__47828),
            .in2(_gnd_net_),
            .in3(N__82297),
            .lcout(\pid_front.N_1674_i ),
            .ltout(\pid_front.N_1674_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_9_17_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_9_17_2 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_8_LC_9_17_2  (
            .in0(N__41474),
            .in1(N__41595),
            .in2(N__41445),
            .in3(N__41614),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_9_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_9_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI873N_11_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__48916),
            .in2(_gnd_net_),
            .in3(N__48895),
            .lcout(\pid_front.un1_pid_prereg_79 ),
            .ltout(\pid_front.un1_pid_prereg_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIROQ33_0_12_LC_9_17_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_0_12_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_0_12_LC_9_17_4 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIROQ33_0_12_LC_9_17_4  (
            .in0(N__43560),
            .in1(N__43502),
            .in2(N__41622),
            .in3(N__43594),
            .lcout(\pid_front.error_p_reg_esr_RNIROQ33_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_7_LC_9_17_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_9_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_7_LC_9_17_5  (
            .in0(N__41615),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83981),
            .ce(N__52540),
            .sr(N__52444));
    defparam \pid_front.error_d_reg_prev_esr_11_LC_9_17_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_9_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_11_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75731),
            .lcout(\pid_front.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83981),
            .ce(N__52540),
            .sr(N__52444));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_17_7 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_11_LC_9_17_7  (
            .in0(N__75730),
            .in1(N__48917),
            .in2(_gnd_net_),
            .in3(N__48896),
            .lcout(\pid_front.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_7_LC_9_18_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_7_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_7_LC_9_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_acumm_7_LC_9_18_0  (
            .in0(N__51705),
            .in1(N__41782),
            .in2(_gnd_net_),
            .in3(N__41580),
            .lcout(\pid_front.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_9_18_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_9_18_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_9_18_1  (
            .in0(N__52137),
            .in1(N__43994),
            .in2(_gnd_net_),
            .in3(N__77629),
            .lcout(\pid_front.error_i_acumm_3_sqmuxa ),
            .ltout(\pid_front.error_i_acumm_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_12_LC_9_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_12_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_12_LC_9_18_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \pid_front.error_i_acumm_12_LC_9_18_2  (
            .in0(N__51702),
            .in1(N__42271),
            .in2(N__41559),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_8_LC_9_18_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_8_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_8_LC_9_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_front.error_i_acumm_8_LC_9_18_3  (
            .in0(N__41783),
            .in1(N__41556),
            .in2(_gnd_net_),
            .in3(N__51706),
            .lcout(\pid_front.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_9_LC_9_18_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_9_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_9_LC_9_18_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_acumm_9_LC_9_18_4  (
            .in0(N__51707),
            .in1(N__41784),
            .in2(_gnd_net_),
            .in3(N__41772),
            .lcout(\pid_front.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_1_LC_9_18_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_1_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_1_LC_9_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_i_acumm_1_LC_9_18_5  (
            .in0(N__41751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51703),
            .lcout(\pid_front.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_2_LC_9_18_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_2_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_2_LC_9_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_i_acumm_2_LC_9_18_6  (
            .in0(N__51704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41736),
            .lcout(\pid_front.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_0_LC_9_18_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_0_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_0_LC_9_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_i_acumm_0_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__42084),
            .in2(_gnd_net_),
            .in3(N__51701),
            .lcout(\pid_front.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83998),
            .ce(N__51647),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_9_19_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_9_19_0 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_9_19_0  (
            .in0(N__41715),
            .in1(N__41706),
            .in2(N__43995),
            .in3(N__54982),
            .lcout(\pid_front.error_i_acumm_2_sqmuxa_1 ),
            .ltout(\pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_9_19_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_9_19_1 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_9_19_1  (
            .in0(N__52130),
            .in1(N__43993),
            .in2(N__41700),
            .in3(N__42231),
            .lcout(\pid_front.error_i_acumm_2_sqmuxa ),
            .ltout(\pid_front.error_i_acumm_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_11_LC_9_19_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_11_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_11_LC_9_19_2 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \pid_front.error_i_acumm_11_LC_9_19_2  (
            .in0(N__41840),
            .in1(N__52132),
            .in2(N__41697),
            .in3(N__41693),
            .lcout(\pid_front.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_4_LC_9_19_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_4_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_4_LC_9_19_3 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_front.error_i_acumm_4_LC_9_19_3  (
            .in0(N__52134),
            .in1(N__41844),
            .in2(N__41670),
            .in3(N__51698),
            .lcout(\pid_front.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_5_LC_9_19_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_5_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_5_LC_9_19_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_front.error_i_acumm_5_LC_9_19_4  (
            .in0(N__51699),
            .in1(N__52135),
            .in2(N__41850),
            .in3(N__41646),
            .lcout(\pid_front.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_6_LC_9_19_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_6_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_6_LC_9_19_5 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_front.error_i_acumm_6_LC_9_19_5  (
            .in0(N__52136),
            .in1(N__41848),
            .in2(N__41898),
            .in3(N__51700),
            .lcout(\pid_front.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_13_LC_9_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_13_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_13_LC_9_19_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_front.error_i_acumm_13_LC_9_19_6  (
            .in0(N__51697),
            .in1(N__52133),
            .in2(N__41849),
            .in3(N__41871),
            .lcout(\pid_front.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_10_LC_9_19_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_10_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_10_LC_9_19_7 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_front.error_i_acumm_10_LC_9_19_7  (
            .in0(N__52131),
            .in1(N__41839),
            .in2(N__41823),
            .in3(N__51696),
            .lcout(\pid_front.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84016),
            .ce(N__51651),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_20_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_20_0  (
            .in0(N__48674),
            .in1(N__41793),
            .in2(N__41964),
            .in3(N__48697),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_9_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_9_20_1 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_9_20_1  (
            .in0(N__84289),
            .in1(N__48610),
            .in2(N__49170),
            .in3(N__46376),
            .lcout(\pid_front.un1_pid_prereg_0_24 ),
            .ltout(\pid_front.un1_pid_prereg_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_9_20_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_9_20_2 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_9_20_2  (
            .in0(N__49215),
            .in1(N__41915),
            .in2(N__41799),
            .in3(N__49197),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_9_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_9_20_3 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_9_20_3  (
            .in0(N__84287),
            .in1(N__48608),
            .in2(N__49169),
            .in3(N__46007),
            .lcout(\pid_front.un1_pid_prereg_0_16 ),
            .ltout(\pid_front.un1_pid_prereg_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_20_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_20_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_20_4  (
            .in0(N__41959),
            .in1(N__45990),
            .in2(N__41796),
            .in3(N__46659),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_20_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_20_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_20_5  (
            .in0(N__41792),
            .in1(N__41960),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_20_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_20_6 .LUT_INIT=16'b0001111010000111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_20_6  (
            .in0(N__48609),
            .in1(N__84288),
            .in2(N__48728),
            .in3(N__49162),
            .lcout(\pid_front.un1_pid_prereg_0_19 ),
            .ltout(\pid_front.un1_pid_prereg_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_20_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_20_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_20_7  (
            .in0(N__48698),
            .in1(_gnd_net_),
            .in2(N__41967),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .LUT_INIT=16'b0101011010010101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0  (
            .in0(N__44120),
            .in1(N__84291),
            .in2(N__48622),
            .in3(N__49152),
            .lcout(\pid_front.un1_pid_prereg_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_9_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_9_21_1 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_9_21_1  (
            .in0(N__84293),
            .in1(N__48603),
            .in2(N__49167),
            .in3(N__44008),
            .lcout(\pid_front.un1_pid_prereg_0_25 ),
            .ltout(\pid_front.un1_pid_prereg_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_9_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_9_21_2 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__41945),
            .in2(N__41949),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_9_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_9_21_3 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_9_21_3  (
            .in0(N__84294),
            .in1(N__48604),
            .in2(N__49168),
            .in3(N__44009),
            .lcout(\pid_front.un1_pid_prereg_0_26 ),
            .ltout(\pid_front.un1_pid_prereg_0_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_9_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_9_21_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_9_21_4  (
            .in0(N__41946),
            .in1(N__41919),
            .in2(N__41934),
            .in3(N__41916),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_5  (
            .in0(N__84292),
            .in1(N__48599),
            .in2(N__49166),
            .in3(N__44119),
            .lcout(\pid_front.un1_pid_prereg_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_9_21_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_9_21_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_front.pid_prereg_esr_RNO_0_30_LC_9_21_6  (
            .in0(N__41927),
            .in1(N__41917),
            .in2(N__41931),
            .in3(N__41918),
            .lcout(\pid_front.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_9_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_9_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_9_21_7  (
            .in0(N__49148),
            .in1(N__84290),
            .in2(_gnd_net_),
            .in3(N__48598),
            .lcout(\pid_front.un1_pid_prereg_370_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_9_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_9_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_0_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__44249),
            .in2(_gnd_net_),
            .in3(N__43656),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_9_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_9_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_9_22_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_21_LC_9_22_1  (
            .in0(N__46452),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_9_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_9_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_9_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_17_LC_9_22_2  (
            .in0(N__43926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_9_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_9_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_22_LC_9_22_3  (
            .in0(N__46677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_9_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_9_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_23_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46011),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_9_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_9_22_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_24_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__44121),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_9_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_9_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_16_LC_9_22_6  (
            .in0(N__48815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_9_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_9_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_25_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48727),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84063),
            .ce(N__46062),
            .sr(N__77350));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIB9VA_4_LC_9_23_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIB9VA_4_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIB9VA_4_LC_9_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIB9VA_4_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41978),
            .lcout(drone_H_disp_front_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_9_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_9_23_4 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_9_23_4  (
            .in0(N__42294),
            .in1(N__42282),
            .in2(N__42273),
            .in3(N__42237),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_1_LC_9_23_5 .C_ON=1'b0;
    defparam \pid_front.error_axb_1_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_1_LC_9_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_1_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42221),
            .lcout(\pid_front.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_3_LC_9_23_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_3_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_3_LC_9_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_3_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42209),
            .lcout(\pid_front.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIPKTD_0_LC_9_28_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIPKTD_0_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIPKTD_0_LC_9_28_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIPKTD_0_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__52185),
            .in2(_gnd_net_),
            .in3(N__77588),
            .lcout(\pid_front.state_RNIPKTDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_10_4_0 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_10_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42177),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83824),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_10_4_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_10_4_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_10_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_10_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42183),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83824),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_10_5_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_10_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_10_5_0  (
            .in0(N__42169),
            .in1(N__42151),
            .in2(N__42134),
            .in3(N__42109),
            .lcout(\Commands_frame_decoder.WDT8lto9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_10_5_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_10_5_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_10_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_10_5_6  (
            .in0(N__48350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42449),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83829),
            .ce(),
            .sr(N__77248));
    defparam \Commands_frame_decoder.source_data_valid_LC_10_5_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_10_5_7 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_10_5_7  (
            .in0(N__42450),
            .in1(N__42093),
            .in2(N__44408),
            .in3(N__48351),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83829),
            .ce(),
            .sr(N__77248));
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_10_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_10_6_2 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \Commands_frame_decoder.preinit_RNIR9JL1_LC_10_6_2  (
            .in0(N__42511),
            .in1(N__42448),
            .in2(N__42392),
            .in3(N__42423),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_10_6_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_10_6_3 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \Commands_frame_decoder.WDT_RNII01C2_8_LC_10_6_3  (
            .in0(N__42605),
            .in1(N__42588),
            .in2(N__42582),
            .in3(N__42557),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lt12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_10_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_10_6_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__42540),
            .in2(N__42534),
            .in3(N__42360),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_6 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_6  (
            .in0(N__42510),
            .in1(N__42489),
            .in2(_gnd_net_),
            .in3(N__42468),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_7 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_7  (
            .in0(N__42447),
            .in1(N__42422),
            .in2(N__42396),
            .in3(N__42383),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_10_7_1 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_10_7_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_drone.state_1_LC_10_7_1  (
            .in0(N__42770),
            .in1(N__43142),
            .in2(N__42645),
            .in3(N__77638),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83842),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_10_7_2 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_10_7_2 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \uart_drone.state_4_LC_10_7_2  (
            .in0(N__77636),
            .in1(N__42903),
            .in2(N__43063),
            .in3(N__42342),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83842),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_10_7_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_10_7_3 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_10_7_3  (
            .in0(N__43049),
            .in1(N__42996),
            .in2(N__42746),
            .in3(N__42949),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_7_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_10_7_4 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_10_7_4  (
            .in0(N__43050),
            .in1(N__42659),
            .in2(N__42783),
            .in3(N__42831),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_10_7_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_10_7_5 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_10_7_5  (
            .in0(N__42742),
            .in1(N__43141),
            .in2(N__42771),
            .in3(N__77635),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_10_7_6 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_10_7_6 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_drone.state_2_LC_10_7_6  (
            .in0(N__42950),
            .in1(N__42769),
            .in2(N__42756),
            .in3(N__42997),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83842),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_10_7_7 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_10_7_7 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \uart_drone.state_3_LC_10_7_7  (
            .in0(N__42902),
            .in1(N__42753),
            .in2(N__42747),
            .in3(N__77637),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83842),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_10_8_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_10_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_10_8_0  (
            .in0(N__42719),
            .in1(N__42707),
            .in2(N__42696),
            .in3(N__42680),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_10_8_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_10_8_1 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_10_8_1  (
            .in0(N__43134),
            .in1(N__42641),
            .in2(_gnd_net_),
            .in3(N__77611),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_10_8_2 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_10_8_2 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_10_8_2  (
            .in0(N__42957),
            .in1(N__42660),
            .in2(N__42648),
            .in3(N__42833),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83850),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_10_8_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_10_8_3  (
            .in0(N__43133),
            .in1(N__42622),
            .in2(_gnd_net_),
            .in3(N__77609),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_8_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_10_8_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_10_8_4  (
            .in0(N__42623),
            .in1(_gnd_net_),
            .in2(N__42609),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_10_8_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_10_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_10_8_5  (
            .in0(N__42855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83850),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_10_8_6 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_10_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42846),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83850),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_10_8_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_10_8_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_10_8_7  (
            .in0(N__43054),
            .in1(N__42832),
            .in2(_gnd_net_),
            .in3(N__77610),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_0 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_10_9_0  (
            .in0(N__44819),
            .in1(N__44773),
            .in2(_gnd_net_),
            .in3(N__44883),
            .lcout(\uart_drone.N_152 ),
            .ltout(\uart_drone.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_9_1 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_10_9_1  (
            .in0(N__43061),
            .in1(_gnd_net_),
            .in2(N__42840),
            .in3(N__43009),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(\uart_drone.un1_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_10_9_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_10_9_2 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \uart_drone.bit_Count_1_LC_10_9_2  (
            .in0(N__43013),
            .in1(N__44774),
            .in2(N__42837),
            .in3(N__44886),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83860),
            .ce(),
            .sr(N__77259));
    defparam \uart_drone.state_RNI62411_4_LC_10_9_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_10_9_3 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_10_9_3  (
            .in0(N__42998),
            .in1(N__42834),
            .in2(N__43065),
            .in3(N__42955),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(\uart_drone.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_9_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42795),
            .in3(N__44884),
            .lcout(),
            .ltout(\uart_drone.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_2_LC_10_9_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_10_9_5 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uart_drone.bit_Count_2_LC_10_9_5  (
            .in0(N__44775),
            .in1(N__42792),
            .in2(N__42786),
            .in3(N__44820),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83860),
            .ce(),
            .sr(N__77259));
    defparam \uart_drone.bit_Count_0_LC_10_9_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_10_9_6 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \uart_drone.bit_Count_0_LC_10_9_6  (
            .in0(N__43202),
            .in1(N__43062),
            .in2(N__43014),
            .in3(N__44885),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83860),
            .ce(),
            .sr(N__77259));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_9_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_10_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_10_9_7  (
            .in0(N__42999),
            .in1(N__43201),
            .in2(_gnd_net_),
            .in3(N__42956),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80481),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73717),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80258),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79713),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_10_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79242),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_10_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_10_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80099),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81059),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83870),
            .ce(N__42887),
            .sr(N__77267));
    defparam \uart_drone.data_Aux_0_LC_10_11_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_10_11_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_0_LC_10_11_0  (
            .in0(N__42864),
            .in1(N__43091),
            .in2(N__43183),
            .in3(N__43229),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_1_LC_10_11_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_10_11_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_10_11_1  (
            .in0(N__43230),
            .in1(N__44571),
            .in2(N__43080),
            .in3(N__43173),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_2_LC_10_11_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_10_11_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_10_11_2  (
            .in0(N__43260),
            .in1(N__43177),
            .in2(N__43374),
            .in3(N__43231),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_3_LC_10_11_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_10_11_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_10_11_3  (
            .in0(N__43232),
            .in1(N__43254),
            .in2(N__43359),
            .in3(N__43174),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_4_LC_10_11_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_10_11_4 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uart_drone.data_Aux_4_LC_10_11_4  (
            .in0(N__43343),
            .in1(N__43248),
            .in2(N__43184),
            .in3(N__43233),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_5_LC_10_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_10_11_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_5_LC_10_11_5  (
            .in0(N__43234),
            .in1(N__44751),
            .in2(N__43332),
            .in3(N__43175),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_6_LC_10_11_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_10_11_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_10_11_6  (
            .in0(N__43242),
            .in1(N__43178),
            .in2(N__43317),
            .in3(N__43235),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_Aux_7_LC_10_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_10_11_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_10_11_7  (
            .in0(N__43236),
            .in1(N__43206),
            .in2(N__43302),
            .in3(N__43176),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83880),
            .ce(),
            .sr(N__43104));
    defparam \uart_drone.data_esr_0_LC_10_12_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43092),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_1_LC_10_12_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43079),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_2_LC_10_12_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43373),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_3_LC_10_12_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43358),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_4_LC_10_12_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43344),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_5_LC_10_12_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_10_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43331),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_6_LC_10_12_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43316),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \uart_drone.data_esr_7_LC_10_12_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43301),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83891),
            .ce(N__43287),
            .sr(N__43275));
    defparam \pid_front.un11lto30_i_a2_0_c_LC_10_13_0 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__44937),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\pid_front.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_LC_10_13_1 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_10_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__43380),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2 ),
            .carryout(\pid_front.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_2_c_LC_10_13_2 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_10_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__45132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_0 ),
            .carryout(\pid_front.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_3_c_LC_10_13_3 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_10_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__43401),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_1 ),
            .carryout(\pid_front.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_4_c_LC_10_13_4 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_10_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_4_c_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__43392),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_2 ),
            .carryout(\pid_front.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_5_c_LC_10_13_5 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_10_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_5_c_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__43464),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_3 ),
            .carryout(\pid_front.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_6_c_LC_10_13_6 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_10_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_6_c_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__43432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_4 ),
            .carryout(\pid_front.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_LC_10_13_7 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_10_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__43447),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_5 ),
            .carryout(\pid_front.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_10_14_0 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_10_14_0 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_10_14_0  (
            .in0(N__45691),
            .in1(N__45740),
            .in2(N__46151),
            .in3(N__43383),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_o2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_10_14_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_10_14_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIN7IV_28_LC_10_14_1  (
            .in0(N__46197),
            .in1(N__46118),
            .in2(_gnd_net_),
            .in3(N__46239),
            .lcout(\pid_front.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_10_14_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_10_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_10_14_2  (
            .in0(N__45789),
            .in1(N__45819),
            .in2(N__46269),
            .in3(N__45861),
            .lcout(\pid_front.un11lto30_i_a2_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_10_14_6 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_10_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_RNO_LC_10_14_6  (
            .in0(N__45361),
            .in1(N__45480),
            .in2(N__45422),
            .in3(N__45313),
            .lcout(\pid_front.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIROQ33_1_12_LC_10_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_1_12_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_1_12_LC_10_15_0 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIROQ33_1_12_LC_10_15_0  (
            .in0(N__43596),
            .in1(N__43555),
            .in2(N__43503),
            .in3(N__43619),
            .lcout(\pid_front.un1_pid_prereg_167_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_12_LC_10_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_12_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_12_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_12_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43488),
            .lcout(\pid_front.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83926),
            .ce(N__83132),
            .sr(N__82875));
    defparam \pid_front.pid_prereg_esr_RNIBQKJ3_20_LC_10_15_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIBQKJ3_20_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIBQKJ3_20_LC_10_15_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIBQKJ3_20_LC_10_15_2  (
            .in0(N__43449),
            .in1(N__43434),
            .in2(_gnd_net_),
            .in3(N__43463),
            .lcout(\pid_front.pid_prereg_esr_RNIBQKJ3Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_10_15_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_10_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNI211A1_20_LC_10_15_3  (
            .in0(N__45885),
            .in1(N__45897),
            .in2(N__45924),
            .in3(N__45909),
            .lcout(\pid_front.un11lto30_i_a2_4_and ),
            .ltout(\pid_front.un11lto30_i_a2_4_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_10_15_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_10_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNID3QC5_15_LC_10_15_4  (
            .in0(N__43448),
            .in1(N__43433),
            .in2(N__43419),
            .in3(N__43416),
            .lcout(\pid_front.N_98 ),
            .ltout(\pid_front.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_10_15_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_10_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIA6N08_0_LC_10_15_5  (
            .in0(N__45153),
            .in1(N__44949),
            .in2(N__43410),
            .in3(N__44931),
            .lcout(),
            .ltout(\pid_front.N_389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIH9GOH_1_LC_10_15_6 .C_ON=1'b0;
    defparam \pid_front.state_RNIH9GOH_1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIH9GOH_1_LC_10_15_6 .LUT_INIT=16'b1110101011101110;
    LogicCell40 \pid_front.state_RNIH9GOH_1_LC_10_15_6  (
            .in0(N__54973),
            .in1(N__52109),
            .in2(N__43407),
            .in3(N__45159),
            .lcout(\pid_front.un1_reset_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNII9PE6_12_LC_10_16_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNII9PE6_12_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNII9PE6_12_LC_10_16_0 .LUT_INIT=16'b1101001000101101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNII9PE6_12_LC_10_16_0  (
            .in0(N__51617),
            .in1(N__78770),
            .in2(N__48020),
            .in3(N__48077),
            .lcout(\pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNII9PE6Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_0_12_LC_10_16_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_0_12_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_0_12_LC_10_16_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUBM0G_0_12_LC_10_16_1  (
            .in0(N__48056),
            .in1(N__43960),
            .in2(N__43404),
            .in3(N__43523),
            .lcout(\pid_front.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJ1FT1_12_LC_10_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJ1FT1_12_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJ1FT1_12_LC_10_16_2 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJ1FT1_12_LC_10_16_2  (
            .in0(N__43554),
            .in1(N__78768),
            .in2(N__43620),
            .in3(N__51612),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIJ1FT1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6J6A4_12_LC_10_16_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6J6A4_12_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6J6A4_12_LC_10_16_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6J6A4_12_LC_10_16_3  (
            .in0(N__43593),
            .in1(N__43530),
            .in2(N__43569),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNI6J6A4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI7FD85_12_LC_10_16_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI7FD85_12_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI7FD85_12_LC_10_16_4 .LUT_INIT=16'b1111010100110001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI7FD85_12_LC_10_16_4  (
            .in0(N__43566),
            .in1(N__51613),
            .in2(N__48019),
            .in3(N__78769),
            .lcout(\pid_front.un1_pid_prereg_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_10_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_10_16_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNICIRCD_14_LC_10_16_5  (
            .in0(N__43688),
            .in1(N__48762),
            .in2(N__48786),
            .in3(N__43671),
            .lcout(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_10_16_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBQB61_12_LC_10_16_6 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBQB61_12_LC_10_16_6  (
            .in0(N__43553),
            .in1(N__51611),
            .in2(_gnd_net_),
            .in3(N__78767),
            .lcout(\pid_front.error_p_reg_esr_RNIBQB61Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_12_LC_10_16_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_12_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUBM0G_12_LC_10_16_7 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUBM0G_12_LC_10_16_7  (
            .in0(N__48057),
            .in1(N__43524),
            .in2(N__43515),
            .in3(N__43961),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIUBM0GZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKGIG5_13_LC_10_17_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKGIG5_13_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKGIG5_13_LC_10_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKGIG5_13_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__48015),
            .in2(_gnd_net_),
            .in3(N__48073),
            .lcout(\pid_front.un1_pid_prereg_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_10_17_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_10_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_10_17_1  (
            .in0(N__49412),
            .in1(N__52640),
            .in2(_gnd_net_),
            .in3(N__43924),
            .lcout(\pid_front.un1_pid_prereg_0_3 ),
            .ltout(\pid_front.un1_pid_prereg_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_10_17_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_10_17_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43506),
            .in3(N__43669),
            .lcout(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_10_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_10_17_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_16_LC_10_17_3  (
            .in0(N__49413),
            .in1(N__52641),
            .in2(_gnd_net_),
            .in3(N__43925),
            .lcout(\pid_front.un1_pid_prereg_0_4 ),
            .ltout(\pid_front.un1_pid_prereg_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_10_17_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_10_17_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNICN0DD_15_LC_10_17_4  (
            .in0(N__43689),
            .in1(N__49025),
            .in2(N__43677),
            .in3(N__43670),
            .lcout(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_10_17_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_10_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_10_17_5  (
            .in0(N__49074),
            .in1(N__49383),
            .in2(_gnd_net_),
            .in3(N__49054),
            .lcout(\pid_front.un1_pid_prereg_0_5 ),
            .ltout(\pid_front.un1_pid_prereg_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_10_17_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_10_17_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43674),
            .in3(N__49007),
            .lcout(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_10_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_10_17_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_10_17_7  (
            .in0(N__51990),
            .in1(N__52692),
            .in2(_gnd_net_),
            .in3(N__48814),
            .lcout(\pid_front.un1_pid_prereg_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_10_18_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_10_18_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNII1MD_0_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__43652),
            .in2(N__44250),
            .in3(_gnd_net_),
            .lcout(\pid_front.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_10_18_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__43641),
            .in2(N__44223),
            .in3(N__43635),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_10_18_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__43632),
            .in2(N__44322),
            .in3(N__43626),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_10_18_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_10_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__51660),
            .in2(N__55413),
            .in3(N__43623),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_10_18_4 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_10_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI9CPM_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__43893),
            .in2(N__55617),
            .in3(N__43866),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNI9CPM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNILQKE_LC_10_18_5 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNILQKE_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNILQKE_LC_10_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNILQKE_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__43863),
            .in2(N__59448),
            .in3(N__43824),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNILQKE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_10_18_6 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__43821),
            .in2(N__59010),
            .in3(N__43794),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_10_18_7 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_10_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIIOSM_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__46758),
            .in2(N__43791),
            .in3(N__43755),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIIOSM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_10_19_0 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__43752),
            .in2(N__58938),
            .in3(N__43719),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_10_19_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__43716),
            .in2(N__44265),
            .in3(N__43710),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_10_19_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__43707),
            .in2(N__50241),
            .in3(N__43701),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_10_19_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__43698),
            .in2(N__55539),
            .in3(N__43692),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_10_19_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIV4AU_12_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__43974),
            .in2(N__55875),
            .in3(N__43968),
            .lcout(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_10_19_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI29BU_13_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__44047),
            .in2(N__47010),
            .in3(N__43965),
            .lcout(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_10_19_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4CCU_14_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__55965),
            .in2(N__44079),
            .in3(N__43935),
            .lcout(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_10_19_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6FDU_15_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__44051),
            .in2(N__53058),
            .in3(N__43932),
            .lcout(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_10_20_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8IEU_16_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__44052),
            .in2(N__44346),
            .in3(N__43929),
            .lcout(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_10_20_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIALFU_17_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__46881),
            .in2(N__44080),
            .in3(N__43905),
            .lcout(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_10_20_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNICOGU_18_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__44056),
            .in2(N__53721),
            .in3(N__43902),
            .lcout(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_10_20_3 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_10_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIERHU_19_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__46836),
            .in2(N__44081),
            .in3(N__43899),
            .lcout(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_10_20_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_10_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI7MJU_20_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__44060),
            .in2(N__55938),
            .in3(N__43896),
            .lcout(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_10_20_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_10_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI08DV_21_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__44172),
            .in2(N__44082),
            .in3(N__44130),
            .lcout(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_10_20_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_10_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI2BEV_22_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__44064),
            .in2(N__56334),
            .in3(N__44127),
            .lcout(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_10_20_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_10_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4EFV_23_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__44142),
            .in2(N__44083),
            .in3(N__44124),
            .lcout(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_10_21_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6HGV_24_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__44084),
            .in2(N__53661),
            .in3(N__44106),
            .lcout(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_10_21_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8KHV_25_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__44280),
            .in2(N__44093),
            .in3(N__44103),
            .lcout(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_10_21_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIANIV_26_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__44088),
            .in2(N__53685),
            .in3(N__44100),
            .lcout(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_10_21_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__44150),
            .in2(N__44094),
            .in3(N__44097),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_10_21_4 .C_ON=1'b0;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_10_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_10_21_4  (
            .in0(N__44151),
            .in1(N__44092),
            .in2(_gnd_net_),
            .in3(N__44013),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_10_21_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_10_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_28_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44010),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84018),
            .ce(N__46065),
            .sr(N__77346));
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_10_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_10_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_27_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46377),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84018),
            .ce(N__46065),
            .sr(N__77346));
    defparam \pid_front.error_i_reg_esr_RNO_7_21_LC_10_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_7_21_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_7_21_LC_10_22_0 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_7_21_LC_10_22_0  (
            .in0(N__71586),
            .in1(N__55822),
            .in2(N__73600),
            .in3(N__53824),
            .lcout(),
            .ltout(\pid_front.g0_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_10_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_10_22_1 .LUT_INIT=16'b1011000010110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_21_LC_10_22_1  (
            .in0(N__73593),
            .in1(N__56157),
            .in2(N__44181),
            .in3(N__55741),
            .lcout(),
            .ltout(\pid_front.N_88_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_10_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_10_22_2 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_21_LC_10_22_2  (
            .in0(N__44163),
            .in1(N__69661),
            .in2(N__44178),
            .in3(N__65751),
            .lcout(),
            .ltout(\pid_front.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_21_LC_10_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_21_LC_10_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_21_LC_10_22_3 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \pid_front.error_i_reg_esr_21_LC_10_22_3  (
            .in0(N__69970),
            .in1(N__44157),
            .in2(N__44175),
            .in3(N__49899),
            .lcout(\pid_front.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84032),
            .ce(N__59377),
            .sr(N__77351));
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_10_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_10_22_4 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_21_LC_10_22_4  (
            .in0(N__71160),
            .in1(N__56512),
            .in2(N__73599),
            .in3(N__56089),
            .lcout(\pid_front.N_126_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_10_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_10_22_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_21_LC_10_22_5  (
            .in0(N__56513),
            .in1(N__69655),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_27_LC_10_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_27_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_27_LC_10_22_6 .LUT_INIT=16'b0100000011100000;
    LogicCell40 \pid_front.error_i_reg_esr_27_LC_10_22_6  (
            .in0(N__69656),
            .in1(N__56514),
            .in2(N__69978),
            .in3(N__55550),
            .lcout(\pid_front.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84032),
            .ce(N__59377),
            .sr(N__77351));
    defparam \pid_front.error_i_reg_esr_23_LC_10_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_23_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_23_LC_10_22_7 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_23_LC_10_22_7  (
            .in0(N__69662),
            .in1(N__46863),
            .in2(N__69977),
            .in3(N__46767),
            .lcout(\pid_front.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84032),
            .ce(N__59377),
            .sr(N__77351));
    defparam \pid_front.error_cry_1_c_RNIT3DD1_LC_10_23_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIT3DD1_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIT3DD1_LC_10_23_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_1_c_RNIT3DD1_LC_10_23_0  (
            .in0(N__71398),
            .in1(N__49973),
            .in2(_gnd_net_),
            .in3(N__50203),
            .lcout(),
            .ltout(\pid_front.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI1VBE3_LC_10_23_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI1VBE3_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI1VBE3_LC_10_23_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_1_c_RNI1VBE3_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__72994),
            .in2(N__44229),
            .in3(N__44211),
            .lcout(\pid_front.N_12_1 ),
            .ltout(\pid_front.N_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_10_23_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_10_23_2 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_17_LC_10_23_2  (
            .in0(N__61672),
            .in1(N__70525),
            .in2(N__44226),
            .in3(N__58912),
            .lcout(\pid_front.m5_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_1_LC_10_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_1_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_1_LC_10_23_3 .LUT_INIT=16'b1000000010110000;
    LogicCell40 \pid_front.error_i_reg_esr_1_LC_10_23_3  (
            .in0(N__58913),
            .in1(N__70748),
            .in2(N__62166),
            .in3(N__44307),
            .lcout(\pid_front.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84048),
            .ce(N__59422),
            .sr(N__77355));
    defparam \pid_front.error_cry_0_0_c_RNI1I0I1_LC_10_23_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI1I0I1_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI1I0I1_LC_10_23_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI1I0I1_LC_10_23_4  (
            .in0(N__71397),
            .in1(N__50356),
            .in2(_gnd_net_),
            .in3(N__50134),
            .lcout(\pid_front.N_9_1 ),
            .ltout(\pid_front.N_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNID6LS3_LC_10_23_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNID6LS3_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNID6LS3_LC_10_23_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNID6LS3_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__72993),
            .in2(N__44205),
            .in3(N__46959),
            .lcout(\pid_front.N_39_0 ),
            .ltout(\pid_front.N_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_10_23_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_10_23_6 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_19_LC_10_23_6  (
            .in0(N__61671),
            .in1(N__55507),
            .in2(N__44202),
            .in3(N__70526),
            .lcout(),
            .ltout(\pid_front.m7_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_10_23_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_10_23_7 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_19_LC_10_23_7  (
            .in0(N__69956),
            .in1(N__69657),
            .in2(N__44199),
            .in3(N__56515),
            .lcout(\pid_front.error_i_reg_9_rn_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNI42002_LC_10_24_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI42002_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI42002_LC_10_24_0 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \pid_front.error_cry_0_c_RNI42002_LC_10_24_0  (
            .in0(N__70517),
            .in1(N__66067),
            .in2(N__69680),
            .in3(N__58911),
            .lcout(\pid_front.un4_error_i_reg_23_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNI7LQG2_LC_10_24_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNI7LQG2_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNI7LQG2_LC_10_24_1 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \pid_front.error_cry_9_c_RNI7LQG2_LC_10_24_1  (
            .in0(N__72982),
            .in1(N__56480),
            .in2(N__71165),
            .in3(N__56078),
            .lcout(\pid_front.N_126 ),
            .ltout(\pid_front.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_10_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_10_24_2 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_25_LC_10_24_2  (
            .in0(N__56481),
            .in1(N__70521),
            .in2(N__44310),
            .in3(N__66066),
            .lcout(\pid_front.m29_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIHILH1_LC_10_24_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIHILH1_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIHILH1_LC_10_24_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \pid_front.error_cry_0_c_RNIHILH1_LC_10_24_3  (
            .in0(N__72981),
            .in1(N__71156),
            .in2(N__61834),
            .in3(N__49630),
            .lcout(\pid_front.m1_0_03 ),
            .ltout(\pid_front.m1_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIM3445_LC_10_24_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIM3445_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIM3445_LC_10_24_4 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \pid_front.error_cry_0_c_RNIM3445_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__44306),
            .in2(N__44295),
            .in3(N__66065),
            .lcout(\pid_front.N_93_0 ),
            .ltout(\pid_front.N_93_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_10_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_10_24_5 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_25_LC_10_24_5  (
            .in0(N__69957),
            .in1(N__69666),
            .in2(N__44292),
            .in3(N__44289),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_25_LC_10_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_25_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_25_LC_10_24_6 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_25_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__59240),
            .in2(N__44283),
            .in3(N__46904),
            .lcout(\pid_front.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84064),
            .ce(N__59424),
            .sr(N__77361));
    defparam \pid_front.error_i_reg_esr_9_LC_10_24_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_9_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_9_LC_10_24_7 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \pid_front.error_i_reg_esr_9_LC_10_24_7  (
            .in0(N__46905),
            .in1(N__65458),
            .in2(N__70530),
            .in3(N__44271),
            .lcout(\pid_front.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84064),
            .ce(N__59424),
            .sr(N__77361));
    defparam \pid_front.error_i_reg_esr_0_LC_10_25_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_0_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_0_LC_10_25_0 .LUT_INIT=16'b1100000001000100;
    LogicCell40 \pid_front.error_i_reg_esr_0_LC_10_25_0  (
            .in0(N__58987),
            .in1(N__62152),
            .in2(N__61749),
            .in3(N__70737),
            .lcout(\pid_front.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84080),
            .ce(N__59423),
            .sr(N__77366));
    defparam \pid_front.error_cry_0_c_RNI634G3_LC_10_25_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI634G3_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI634G3_LC_10_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_front.error_cry_0_c_RNI634G3_LC_10_25_1  (
            .in0(N__50091),
            .in1(N__55994),
            .in2(_gnd_net_),
            .in3(N__72908),
            .lcout(\pid_front.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_10_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_10_25_2 .LUT_INIT=16'b1000111100000111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_16_LC_10_25_2  (
            .in0(N__73601),
            .in1(N__66069),
            .in2(N__56527),
            .in3(N__56034),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_2Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_10_25_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_10_25_3 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_16_LC_10_25_3  (
            .in0(N__69915),
            .in1(N__69659),
            .in2(N__44352),
            .in3(N__44334),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_16_LC_10_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_16_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_16_LC_10_25_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_16_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__61914),
            .in2(N__44349),
            .in3(N__44328),
            .lcout(\pid_front.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84080),
            .ce(N__59423),
            .sr(N__77366));
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_10_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_10_25_5 .LUT_INIT=16'b0000100000001101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_16_LC_10_25_5  (
            .in0(N__66068),
            .in1(N__61745),
            .in2(N__70529),
            .in3(N__58986),
            .lcout(\pid_front.m4_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_10_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_10_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_16_LC_10_25_6  (
            .in0(N__70733),
            .in1(N__53616),
            .in2(_gnd_net_),
            .in3(N__55907),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_2_LC_10_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_2_LC_10_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_2_LC_10_26_3 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_2_LC_10_26_3  (
            .in0(N__70741),
            .in1(N__59202),
            .in2(N__62165),
            .in3(N__56382),
            .lcout(\pid_front.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84090),
            .ce(N__59427),
            .sr(N__77372));
    defparam \ppm_encoder_1.throttle_4_LC_11_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_11_7_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_11_7_2  (
            .in0(N__47181),
            .in1(N__47214),
            .in2(N__62674),
            .in3(N__59152),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83834),
            .ce(),
            .sr(N__77253));
    defparam \ppm_encoder_1.throttle_5_LC_11_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_11_7_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_11_7_3  (
            .in0(N__47136),
            .in1(N__47169),
            .in2(N__57001),
            .in3(N__62604),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83834),
            .ce(),
            .sr(N__77253));
    defparam \ppm_encoder_1.throttle_9_LC_11_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_11_7_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_11_7_4  (
            .in0(N__47115),
            .in1(N__47085),
            .in2(N__62675),
            .in3(N__56914),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83834),
            .ce(),
            .sr(N__77253));
    defparam \scaler_4.source_data_1_4_LC_11_7_5 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_11_7_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \scaler_4.source_data_1_4_LC_11_7_5  (
            .in0(N__44404),
            .in1(N__44535),
            .in2(N__47289),
            .in3(N__47390),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83834),
            .ce(),
            .sr(N__77253));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_7_6 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_7_6  (
            .in0(N__44498),
            .in1(N__47285),
            .in2(_gnd_net_),
            .in3(N__44534),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_11_7_7 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_11_7_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \scaler_4.source_data_1_esr_ctle_14_LC_11_7_7  (
            .in0(N__44403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77615),
            .lcout(\scaler_4.debug_CH3_20A_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_11_8_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_11_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__44494),
            .in2(N__44379),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_11_8_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__44459),
            .in2(N__44499),
            .in3(N__44370),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_7_LC_11_8_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__44435),
            .in2(N__44463),
            .in3(N__44367),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_8_LC_11_8_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__44741),
            .in2(N__44439),
            .in3(N__44364),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_9_LC_11_8_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_11_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__44717),
            .in2(N__44745),
            .in3(N__44361),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_10_LC_11_8_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__44693),
            .in2(N__44721),
            .in3(N__44358),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_11_LC_11_8_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_11_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__44660),
            .in2(N__44697),
            .in3(N__44355),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_12_LC_11_8_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_11_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__44645),
            .in2(N__44664),
            .in3(N__44565),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__83843),
            .ce(N__44549),
            .sr(N__77260));
    defparam \scaler_4.source_data_1_esr_13_LC_11_9_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__44646),
            .in2(N__44625),
            .in3(N__44562),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__83851),
            .ce(N__44556),
            .sr(N__77268));
    defparam \scaler_4.source_data_1_esr_14_LC_11_9_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44559),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83851),
            .ce(N__44556),
            .sr(N__77268));
    defparam \scaler_4.source_data_1_esr_5_LC_11_9_3 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_11_9_3  (
            .in0(N__44493),
            .in1(N__47284),
            .in2(_gnd_net_),
            .in3(N__44527),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83851),
            .ce(N__44556),
            .sr(N__77268));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_10_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__44521),
            .in2(N__47278),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_10_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__44505),
            .in2(N__47256),
            .in3(N__44472),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_10_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__44469),
            .in2(N__47247),
            .in3(N__44448),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_10_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__44445),
            .in2(N__47238),
            .in3(N__44424),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_10_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__44421),
            .in2(N__47229),
            .in3(N__44730),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_10_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__44727),
            .in2(N__47439),
            .in3(N__44706),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_10_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__44703),
            .in2(N__47430),
            .in3(N__44682),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_10_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__44679),
            .in2(_gnd_net_),
            .in3(N__44649),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_11_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__44577),
            .in2(N__60526),
            .in3(N__44631),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_11_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44628),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__44613),
            .in2(_gnd_net_),
            .in3(N__77633),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_2232_i_l_ofx_LC_11_11_4 .C_ON=1'b0;
    defparam \scaler_4.N_2232_i_l_ofx_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_2232_i_l_ofx_LC_11_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_2232_i_l_ofx_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__47417),
            .in2(_gnd_net_),
            .in3(N__44595),
            .lcout(\scaler_4.N_2232_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_11_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_11_11_5  (
            .in0(N__44798),
            .in1(N__44851),
            .in2(_gnd_net_),
            .in3(N__44911),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_11_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_11_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_11_11_6  (
            .in0(N__44912),
            .in1(_gnd_net_),
            .in2(N__44859),
            .in3(N__44799),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_12_LC_11_12_0 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_12_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_12_LC_11_12_0 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \pid_front.source_pid_1_esr_12_LC_11_12_0  (
            .in0(N__45742),
            .in1(N__46157),
            .in2(N__45699),
            .in3(N__45185),
            .lcout(front_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_13_LC_11_12_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_13_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_13_LC_11_12_1 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \pid_front.source_pid_1_esr_13_LC_11_12_1  (
            .in0(N__45186),
            .in1(_gnd_net_),
            .in2(N__46167),
            .in3(N__45695),
            .lcout(front_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_10_LC_11_12_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_10_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_10_LC_11_12_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_10_LC_11_12_2  (
            .in0(N__45109),
            .in1(N__46154),
            .in2(_gnd_net_),
            .in3(N__45210),
            .lcout(front_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_11_LC_11_12_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_11_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_11_LC_11_12_3 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \pid_front.source_pid_1_esr_11_LC_11_12_3  (
            .in0(N__45772),
            .in1(_gnd_net_),
            .in2(N__46166),
            .in3(N__45114),
            .lcout(front_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_6_LC_11_12_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_6_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_6_LC_11_12_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_6_LC_11_12_4  (
            .in0(N__45110),
            .in1(N__46155),
            .in2(_gnd_net_),
            .in3(N__45366),
            .lcout(front_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_7_LC_11_12_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_7_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_7_LC_11_12_5 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_7_LC_11_12_5  (
            .in0(N__46152),
            .in1(N__45112),
            .in2(_gnd_net_),
            .in3(N__45315),
            .lcout(front_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_8_LC_11_12_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_8_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_8_LC_11_12_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_8_LC_11_12_6  (
            .in0(N__45111),
            .in1(N__46156),
            .in2(_gnd_net_),
            .in3(N__45258),
            .lcout(front_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.source_pid_1_esr_9_LC_11_12_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_9_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_9_LC_11_12_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_9_LC_11_12_7  (
            .in0(N__46153),
            .in1(N__45113),
            .in2(_gnd_net_),
            .in3(N__45234),
            .lcout(front_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83881),
            .ce(N__47321),
            .sr(N__47364));
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_11_13_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_11_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIVFPG_1_LC_11_13_1  (
            .in0(N__44966),
            .in1(N__45423),
            .in2(N__45525),
            .in3(N__44984),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_11_13_2 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_11_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_RNO_LC_11_13_2  (
            .in0(N__44983),
            .in1(N__44965),
            .in2(N__45524),
            .in3(N__45001),
            .lcout(\pid_front.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_11_13_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_11_13_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI6TRI_0_LC_11_13_3  (
            .in0(N__45002),
            .in1(N__45741),
            .in2(_gnd_net_),
            .in3(N__45486),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_1_LC_11_13_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_1_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_1_LC_11_13_4 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_front.source_pid_1_esr_1_LC_11_13_4  (
            .in0(N__44985),
            .in1(N__45056),
            .in2(N__45125),
            .in3(N__46149),
            .lcout(front_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83892),
            .ce(N__47320),
            .sr(N__47358));
    defparam \pid_front.source_pid_1_esr_2_LC_11_13_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_2_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_2_LC_11_13_5 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_front.source_pid_1_esr_2_LC_11_13_5  (
            .in0(N__44967),
            .in1(N__45062),
            .in2(N__46165),
            .in3(N__45124),
            .lcout(front_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83892),
            .ce(N__47320),
            .sr(N__47358));
    defparam \pid_front.source_pid_1_esr_3_LC_11_13_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_3_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_3_LC_11_13_6 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_front.source_pid_1_esr_3_LC_11_13_6  (
            .in0(N__45520),
            .in1(N__45057),
            .in2(N__45126),
            .in3(N__46150),
            .lcout(front_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83892),
            .ce(N__47320),
            .sr(N__47358));
    defparam \pid_front.source_pid_1_esr_0_LC_11_13_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_0_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_0_LC_11_13_7 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_front.source_pid_1_esr_0_LC_11_13_7  (
            .in0(N__45003),
            .in1(N__45061),
            .in2(N__46164),
            .in3(N__45123),
            .lcout(front_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83892),
            .ce(N__47320),
            .sr(N__47358));
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_11_14_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_11_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI4ABT_6_LC_11_14_0  (
            .in0(N__45314),
            .in1(N__45209),
            .in2(N__45774),
            .in3(N__45362),
            .lcout(),
            .ltout(\pid_front.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_14_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_11_14_1  (
            .in0(N__45257),
            .in1(N__45694),
            .in2(N__44919),
            .in3(N__45233),
            .lcout(\pid_front.N_99 ),
            .ltout(\pid_front.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_14_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_14_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI3Q532_4_LC_11_14_2  (
            .in0(N__46122),
            .in1(N__45420),
            .in2(N__44916),
            .in3(N__45484),
            .lcout(\pid_front.N_75 ),
            .ltout(\pid_front.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_11_14_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_11_14_3 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \pid_front.pid_prereg_esr_RNIDDR99_30_LC_11_14_3  (
            .in0(N__45179),
            .in1(N__45168),
            .in2(N__45162),
            .in3(N__46123),
            .lcout(\pid_front.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_5_LC_11_14_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_5_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_5_LC_11_14_5 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \pid_front.source_pid_1_esr_5_LC_11_14_5  (
            .in0(N__45421),
            .in1(N__45116),
            .in2(N__45152),
            .in3(N__46125),
            .lcout(front_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83901),
            .ce(N__47322),
            .sr(N__47363));
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_14_6 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_RNO_LC_11_14_6  (
            .in0(N__45232),
            .in1(N__45208),
            .in2(N__45773),
            .in3(N__45256),
            .lcout(\pid_front.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_4_LC_11_14_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_4_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_4_LC_11_14_7 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \pid_front.source_pid_1_esr_4_LC_11_14_7  (
            .in0(N__45485),
            .in1(N__45115),
            .in2(N__45063),
            .in3(N__46124),
            .lcout(front_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83901),
            .ce(N__47322),
            .sr(N__47363));
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_11_15_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__45029),
            .in2(N__45033),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_0_LC_11_15_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_0_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_0_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__52929),
            .in2(N__52976),
            .in3(N__44988),
            .lcout(\pid_front.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_1_LC_11_15_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_1_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_1_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_1_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__52236),
            .in2(N__52277),
            .in3(N__44970),
            .lcout(\pid_front.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_1 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_2_LC_11_15_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_2_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_2_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_2_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__49320),
            .in2(N__49357),
            .in3(N__44952),
            .lcout(\pid_front.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_2 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_3_LC_11_15_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_3_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_3_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_3_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__49280),
            .in2(N__47580),
            .in3(N__45501),
            .lcout(\pid_front.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_3 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_4_LC_11_15_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_4_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_4_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_4_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__45498),
            .in2(N__47525),
            .in3(N__45462),
            .lcout(\pid_front.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_4 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_5_LC_11_15_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_5_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_5_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_5_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__45459),
            .in2(N__45438),
            .in3(N__45396),
            .lcout(\pid_front.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_5 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_6_LC_11_15_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_6_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_6_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_6_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__45393),
            .in2(N__45381),
            .in3(N__45345),
            .lcout(\pid_front.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_6 ),
            .clk(N__83914),
            .ce(N__46069),
            .sr(N__77314));
    defparam \pid_front.pid_prereg_esr_7_LC_11_16_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_7_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_7_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_7_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__45342),
            .in2(N__45333),
            .in3(N__45291),
            .lcout(\pid_front.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_7 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_8_LC_11_16_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_8_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_8_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_8_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__45288),
            .in2(N__45279),
            .in3(N__45237),
            .lcout(\pid_front.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_8 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_9_LC_11_16_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_9_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_9_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_9_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__47739),
            .in2(N__47789),
            .in3(N__45213),
            .lcout(\pid_front.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_9 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_10_LC_11_16_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_10_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_10_LC_11_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_10_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__47892),
            .in2(N__47886),
            .in3(N__45189),
            .lcout(\pid_front.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_10 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_11_LC_11_16_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_11_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_11_LC_11_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_11_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__48107),
            .in2(N__47940),
            .in3(N__45747),
            .lcout(\pid_front.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_11 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_12_LC_11_16_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_12_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_12_LC_11_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_12_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__51855),
            .in2(N__48096),
            .in3(N__45702),
            .lcout(\pid_front.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_12 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.pid_prereg_esr_13_LC_11_16_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_13_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_13_LC_11_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_13_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__51968),
            .in2(N__51954),
            .in3(N__45654),
            .lcout(\pid_front.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_13 ),
            .clk(N__83927),
            .ce(N__46068),
            .sr(N__77320));
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_11_16_7 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_11_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__45650),
            .in2(_gnd_net_),
            .in3(N__45627),
            .lcout(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_15_LC_11_17_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_15_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_15_LC_11_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_15_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__48504),
            .in2(N__48521),
            .in3(N__45606),
            .lcout(\pid_front.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_15 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_16_LC_11_17_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_16_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_16_LC_11_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_16_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__48498),
            .in2(N__48480),
            .in3(N__45588),
            .lcout(\pid_front.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_16 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_17_LC_11_17_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_17_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_17_LC_11_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_17_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__45585),
            .in2(N__48744),
            .in3(N__45564),
            .lcout(\pid_front.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_17 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_18_LC_11_17_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_18_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_18_LC_11_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_18_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__45561),
            .in2(N__45555),
            .in3(N__45528),
            .lcout(\pid_front.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_18 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_19_LC_11_17_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_19_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_19_LC_11_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_19_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__45951),
            .in2(N__48993),
            .in3(N__45927),
            .lcout(\pid_front.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_19 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_20_LC_11_17_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_20_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_20_LC_11_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_20_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__46395),
            .in2(N__49449),
            .in3(N__45912),
            .lcout(\pid_front.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_20 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_21_LC_11_17_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_21_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_21_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_21_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__46278),
            .in2(N__45963),
            .in3(N__45900),
            .lcout(\pid_front.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_21 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_22_LC_11_17_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_22_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_22_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_22_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__46347),
            .in2(N__46710),
            .in3(N__45888),
            .lcout(\pid_front.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_22 ),
            .clk(N__83939),
            .ce(N__46067),
            .sr(N__77328));
    defparam \pid_front.pid_prereg_esr_23_LC_11_18_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_23_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_23_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_23_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__45969),
            .in2(N__46386),
            .in3(N__45876),
            .lcout(\pid_front.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_23 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_24_LC_11_18_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_24_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_24_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_24_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__45873),
            .in2(N__46020),
            .in3(N__45849),
            .lcout(\pid_front.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_24 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_25_LC_11_18_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_25_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_25_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_25_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__45846),
            .in2(N__45834),
            .in3(N__45807),
            .lcout(\pid_front.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_25 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_26_LC_11_18_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_26_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_26_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_26_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__48663),
            .in2(N__45804),
            .in3(N__45777),
            .lcout(\pid_front.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_26 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_27_LC_11_18_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_27_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_27_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_27_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__49254),
            .in2(N__49224),
            .in3(N__46254),
            .lcout(\pid_front.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_27 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_28_LC_11_18_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_28_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_28_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_28_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__46251),
            .in2(N__49179),
            .in3(N__46227),
            .lcout(\pid_front.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_28 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_29_LC_11_18_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_29_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_29_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_29_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__46224),
            .in2(N__46212),
            .in3(N__46185),
            .lcout(\pid_front.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_29 ),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.pid_prereg_esr_30_LC_11_18_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_30_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_30_LC_11_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.pid_prereg_esr_30_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__46182),
            .in2(_gnd_net_),
            .in3(N__46170),
            .lcout(\pid_front.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83953),
            .ce(N__46066),
            .sr(N__77335));
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_11_19_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_11_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__45983),
            .in2(_gnd_net_),
            .in3(N__46654),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_11_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_11_19_1 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_11_19_1  (
            .in0(N__84302),
            .in1(N__48611),
            .in2(N__49144),
            .in3(N__46006),
            .lcout(\pid_front.un1_pid_prereg_0_15 ),
            .ltout(\pid_front.un1_pid_prereg_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_11_19_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_11_19_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_11_19_2  (
            .in0(N__46359),
            .in1(N__46431),
            .in2(N__45972),
            .in3(N__46655),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_11_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_11_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__46292),
            .in2(_gnd_net_),
            .in3(N__46310),
            .lcout(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_11_19_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_11_19_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_11_19_4  (
            .in0(N__48980),
            .in1(N__52599),
            .in2(_gnd_net_),
            .in3(N__48955),
            .lcout(\pid_front.un1_pid_prereg_0_8 ),
            .ltout(\pid_front.un1_pid_prereg_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_11_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_11_19_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI80EDD_17_LC_11_19_5  (
            .in0(N__49461),
            .in1(N__48936),
            .in2(N__46398),
            .in3(N__46309),
            .lcout(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_11_19_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_11_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_11_19_6  (
            .in0(N__46791),
            .in1(N__48380),
            .in2(_gnd_net_),
            .in3(N__46330),
            .lcout(\pid_front.un1_pid_prereg_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_11_19_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_11_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNID7NO6_20_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__46358),
            .in2(_gnd_net_),
            .in3(N__46430),
            .lcout(\pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_11_20_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_11_20_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_11_20_0  (
            .in0(N__84301),
            .in1(N__48631),
            .in2(N__49147),
            .in3(N__46375),
            .lcout(\pid_front.un1_pid_prereg_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_11_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_11_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_11_20_1  (
            .in0(N__46823),
            .in1(N__46694),
            .in2(_gnd_net_),
            .in3(N__46672),
            .lcout(\pid_front.un1_pid_prereg_0_13 ),
            .ltout(\pid_front.un1_pid_prereg_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_11_20_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_11_20_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_11_20_2  (
            .in0(N__46725),
            .in1(N__46737),
            .in2(N__46350),
            .in3(N__46423),
            .lcout(\pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_11_20_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_11_20_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_11_20_3  (
            .in0(N__46790),
            .in1(N__48387),
            .in2(_gnd_net_),
            .in3(N__46331),
            .lcout(\pid_front.un1_pid_prereg_0_10 ),
            .ltout(\pid_front.un1_pid_prereg_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_11_20_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_11_20_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNISOJED_18_LC_11_20_4  (
            .in0(N__46314),
            .in1(N__46296),
            .in2(N__46281),
            .in3(N__46736),
            .lcout(\pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_11_20_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_11_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_11_20_5  (
            .in0(N__46410),
            .in1(N__46461),
            .in2(_gnd_net_),
            .in3(N__46448),
            .lcout(\pid_front.un1_pid_prereg_0_11 ),
            .ltout(\pid_front.un1_pid_prereg_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_11_20_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_11_20_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI20QN6_19_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46728),
            .in3(N__46721),
            .lcout(\pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_11_20_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_11_20_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_11_20_7  (
            .in0(N__46824),
            .in1(N__46695),
            .in2(_gnd_net_),
            .in3(N__46673),
            .lcout(\pid_front.un1_pid_prereg_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_5_LC_11_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_11_21_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_11_21_0  (
            .in0(N__46641),
            .in1(N__46532),
            .in2(N__46602),
            .in3(N__47684),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84000),
            .ce(),
            .sr(N__46518));
    defparam \pid_front.error_cry_0_c_RNIPTAD1_LC_11_21_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIPTAD1_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIPTAD1_LC_11_21_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_0_c_RNIPTAD1_LC_11_21_1  (
            .in0(N__71447),
            .in1(N__49620),
            .in2(_gnd_net_),
            .in3(N__49960),
            .lcout(\pid_front.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIFP1H1_LC_11_21_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_8_c_RNIFP1H1_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIFP1H1_LC_11_21_2 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \pid_front.error_cry_8_c_RNIFP1H1_LC_11_21_2  (
            .in0(N__55723),
            .in1(_gnd_net_),
            .in2(N__56158),
            .in3(N__71154),
            .lcout(\pid_front.N_45_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_21_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_21_3  (
            .in0(N__48632),
            .in1(N__51554),
            .in2(_gnd_net_),
            .in3(N__84349),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_21_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__46409),
            .in2(N__46455),
            .in3(N__46447),
            .lcout(\pid_front.un1_pid_prereg_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_21_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_21_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_21_5  (
            .in0(N__46815),
            .in1(N__51576),
            .in2(_gnd_net_),
            .in3(N__84395),
            .lcout(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_21_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_21_6  (
            .in0(N__84350),
            .in1(_gnd_net_),
            .in2(N__51558),
            .in3(N__48633),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_21_7  (
            .in0(N__46814),
            .in1(N__51575),
            .in2(_gnd_net_),
            .in3(N__84394),
            .lcout(\pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNID0MD1_LC_11_22_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNID0MD1_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNID0MD1_LC_11_22_0 .LUT_INIT=16'b0001100101011101;
    LogicCell40 \pid_front.error_cry_0_c_RNID0MD1_LC_11_22_0  (
            .in0(N__71454),
            .in1(N__73308),
            .in2(N__61814),
            .in3(N__49609),
            .lcout(),
            .ltout(\pid_front.m14_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIS4023_LC_11_22_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIS4023_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIS4023_LC_11_22_1 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_front.error_cry_1_c_RNIS4023_LC_11_22_1  (
            .in0(N__72972),
            .in1(N__49959),
            .in2(N__46776),
            .in3(N__50193),
            .lcout(\pid_front.N_15_1 ),
            .ltout(\pid_front.N_15_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI7L6B3_LC_11_22_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI7L6B3_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI7L6B3_LC_11_22_2 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \pid_front.error_cry_1_c_RNI7L6B3_LC_11_22_2  (
            .in0(N__70492),
            .in1(_gnd_net_),
            .in2(N__46773),
            .in3(N__66042),
            .lcout(),
            .ltout(\pid_front.m104_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI6I86D_LC_11_22_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI6I86D_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI6I86D_LC_11_22_3 .LUT_INIT=16'b1101000011010011;
    LogicCell40 \pid_front.error_cry_1_c_RNI6I86D_LC_11_22_3  (
            .in0(N__53112),
            .in1(N__70493),
            .in2(N__46770),
            .in3(N__55429),
            .lcout(\pid_front.m11_2_03_3_i_0 ),
            .ltout(\pid_front.m11_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_7_LC_11_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_7_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_7_LC_11_22_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \pid_front.error_i_reg_7_LC_11_22_4  (
            .in0(N__55583),
            .in1(N__65441),
            .in2(N__46761),
            .in3(N__46754),
            .lcout(\pid_front.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84019),
            .ce(),
            .sr(N__77356));
    defparam \pid_front.error_cry_1_c_RNI3KQB7_LC_11_22_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI3KQB7_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI3KQB7_LC_11_22_5 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_1_c_RNI3KQB7_LC_11_22_5  (
            .in0(N__61655),
            .in1(N__55506),
            .in2(N__70516),
            .in3(N__55428),
            .lcout(),
            .ltout(\pid_front.m53_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIDC92H_LC_11_22_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIDC92H_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIDC92H_LC_11_22_6 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_front.error_cry_1_c_RNIDC92H_LC_11_22_6  (
            .in0(N__70491),
            .in1(N__53111),
            .in2(N__46740),
            .in3(N__53080),
            .lcout(\pid_front.N_54_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_11_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_11_23_0 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_17_LC_11_23_0  (
            .in0(N__69658),
            .in1(N__46851),
            .in2(N__69969),
            .in3(N__46890),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_17_LC_11_23_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_17_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_17_LC_11_23_1 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_17_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__61912),
            .in2(N__46884),
            .in3(N__46965),
            .lcout(\pid_front.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84033),
            .ce(N__59345),
            .sr(N__77362));
    defparam \pid_front.error_cry_9_c_RNI4CS12_LC_11_23_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNI4CS12_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNI4CS12_LC_11_23_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_9_c_RNI4CS12_LC_11_23_2  (
            .in0(N__71155),
            .in1(N__56440),
            .in2(_gnd_net_),
            .in3(N__56062),
            .lcout(\pid_front.N_44_1 ),
            .ltout(\pid_front.N_44_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIO12O3_LC_11_23_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_8_c_RNIO12O3_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIO12O3_LC_11_23_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_front.error_cry_8_c_RNIO12O3_LC_11_23_3  (
            .in0(N__73567),
            .in1(_gnd_net_),
            .in2(N__46869),
            .in3(N__46947),
            .lcout(\pid_front.N_46_1 ),
            .ltout(\pid_front.N_46_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_11_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_11_23_4 .LUT_INIT=16'b1000000011110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_23_LC_11_23_4  (
            .in0(N__70747),
            .in1(N__70513),
            .in2(N__46866),
            .in3(N__56441),
            .lcout(\pid_front.m27_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_11_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_11_23_5 .LUT_INIT=16'b1011001100010011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_17_LC_11_23_5  (
            .in0(N__73568),
            .in1(N__56467),
            .in2(N__66064),
            .in3(N__46857),
            .lcout(\pid_front.error_i_reg_esr_RNO_2Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_11_23_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_11_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_19_LC_11_23_6  (
            .in0(N__65743),
            .in1(N__53110),
            .in2(_gnd_net_),
            .in3(N__53081),
            .lcout(),
            .ltout(\pid_front.N_50_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_19_LC_11_23_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_19_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_19_LC_11_23_7 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \pid_front.error_i_reg_esr_19_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(N__61913),
            .in2(N__46845),
            .in3(N__46842),
            .lcout(\pid_front.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84033),
            .ce(N__59345),
            .sr(N__77362));
    defparam \pid_front.error_i_reg_esr_RNO_12_21_LC_11_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_12_21_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_12_21_LC_11_24_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_12_21_LC_11_24_0  (
            .in0(N__73286),
            .in1(N__50282),
            .in2(N__71467),
            .in3(N__53492),
            .lcout(\pid_front.g0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_11_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_11_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_17_LC_11_24_1  (
            .in0(N__65735),
            .in1(N__46923),
            .in2(_gnd_net_),
            .in3(N__46914),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNI9BMR1_LC_11_24_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNI9BMR1_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNI9BMR1_LC_11_24_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_1_0_c_RNI9BMR1_LC_11_24_2  (
            .in0(N__72675),
            .in1(N__50281),
            .in2(_gnd_net_),
            .in3(N__53493),
            .lcout(\pid_front.N_51_1 ),
            .ltout(\pid_front.N_51_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNITD7Q3_LC_11_24_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNITD7Q3_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNITD7Q3_LC_11_24_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNITD7Q3_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__73574),
            .in2(N__46953),
            .in3(N__53043),
            .lcout(\pid_front.N_89_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIRFVG1_LC_11_24_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIRFVG1_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIRFVG1_LC_11_24_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_5_c_RNIRFVG1_LC_11_24_4  (
            .in0(N__72676),
            .in1(N__55797),
            .in2(_gnd_net_),
            .in3(N__53804),
            .lcout(),
            .ltout(\pid_front.N_47_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIF5573_LC_11_24_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIF5573_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIF5573_LC_11_24_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_5_c_RNIF5573_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__73573),
            .in2(N__46950),
            .in3(N__46946),
            .lcout(\pid_front.N_88_0 ),
            .ltout(\pid_front.N_88_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_11_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_11_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_13_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__46932),
            .in2(N__46926),
            .in3(N__65734),
            .lcout(\pid_front.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIH9L97_LC_11_24_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIH9L97_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIH9L97_LC_11_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIH9L97_LC_11_24_7  (
            .in0(N__65733),
            .in1(N__46922),
            .in2(_gnd_net_),
            .in3(N__46913),
            .lcout(\pid_front.N_90_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIH0F73_LC_11_25_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIH0F73_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIH0F73_LC_11_25_0 .LUT_INIT=16'b1010001010100111;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIH0F73_LC_11_25_0  (
            .in0(N__46896),
            .in1(N__50354),
            .in2(N__73306),
            .in3(N__50132),
            .lcout(\pid_front.N_12_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIFDEL1_LC_11_25_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIFDEL1_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIFDEL1_LC_11_25_1 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_front.error_cry_1_c_RNIFDEL1_LC_11_25_1  (
            .in0(N__73287),
            .in1(N__49974),
            .in2(N__71468),
            .in3(N__50195),
            .lcout(\pid_front.g0_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIATU12_LC_11_25_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIATU12_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIATU12_LC_11_25_2 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIATU12_LC_11_25_2  (
            .in0(N__73295),
            .in1(N__50296),
            .in2(N__71469),
            .in3(N__53508),
            .lcout(),
            .ltout(\pid_front.g0_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI9DJP3_LC_11_25_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI9DJP3_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI9DJP3_LC_11_25_3 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_front.error_cry_4_c_RNI9DJP3_LC_11_25_3  (
            .in0(N__73288),
            .in1(N__53568),
            .in2(N__47043),
            .in3(N__53866),
            .lcout(),
            .ltout(\pid_front.N_89_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIDO397_LC_11_25_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIDO397_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIDO397_LC_11_25_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIDO397_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__61673),
            .in2(N__47040),
            .in3(N__47037),
            .lcout(\pid_front.N_116_0 ),
            .ltout(\pid_front.N_116_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_11_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_11_25_5 .LUT_INIT=16'b0101010100000101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_13_LC_11_25_5  (
            .in0(N__69660),
            .in1(_gnd_net_),
            .in2(N__47031),
            .in3(N__47027),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_13_LC_11_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_13_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_13_LC_11_25_6 .LUT_INIT=16'b0100100011001000;
    LogicCell40 \pid_front.error_i_reg_esr_13_LC_11_25_6  (
            .in0(N__47028),
            .in1(N__69872),
            .in2(N__47019),
            .in3(N__47016),
            .lcout(\pid_front.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84065),
            .ce(N__59346),
            .sr(N__77373));
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_5_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_5_2 .LUT_INIT=16'b1010101011001110;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_12_5_2  (
            .in0(N__46985),
            .in1(N__46974),
            .in2(N__56316),
            .in3(N__50391),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83821),
            .ce(),
            .sr(N__77250));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__56720),
            .in2(_gnd_net_),
            .in3(N__56264),
            .lcout(\ppm_encoder_1.N_134_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_7_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__62414),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_7_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__50531),
            .in2(_gnd_net_),
            .in3(N__46968),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_7_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__50960),
            .in2(_gnd_net_),
            .in3(N__47073),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_7_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__50921),
            .in2(_gnd_net_),
            .in3(N__47070),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_7_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__50459),
            .in2(_gnd_net_),
            .in3(N__47067),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_7_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__51038),
            .in2(_gnd_net_),
            .in3(N__47064),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_7_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__50978),
            .in2(_gnd_net_),
            .in3(N__47061),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_7_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__50444),
            .in2(N__60586),
            .in3(N__47058),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__47055),
            .in2(_gnd_net_),
            .in3(N__47049),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83835),
            .ce(N__60713),
            .sr(N__77269));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__59537),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__50904),
            .in2(N__60537),
            .in3(N__47046),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__62810),
            .in2(_gnd_net_),
            .in3(N__47220),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__59663),
            .in2(N__60538),
            .in3(N__47217),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__47210),
            .in2(_gnd_net_),
            .in3(N__47172),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__47165),
            .in2(_gnd_net_),
            .in3(N__47127),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__60484),
            .in2(N__50648),
            .in3(N__47124),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__50834),
            .in2(_gnd_net_),
            .in3(N__47121),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__54403),
            .in2(_gnd_net_),
            .in3(N__47118),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__47107),
            .in2(_gnd_net_),
            .in3(N__47076),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__50876),
            .in2(_gnd_net_),
            .in3(N__47304),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__50741),
            .in2(_gnd_net_),
            .in3(N__47301),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__54686),
            .in2(_gnd_net_),
            .in3(N__47298),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__57287),
            .in2(N__60536),
            .in3(N__47295),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47292),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83852),
            .ce(N__60724),
            .sr(N__77278));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_12_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80505),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_12_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_12_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_12_11_1  (
            .in0(N__73721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_12_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_12_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80238),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_12_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_12_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79725),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_12_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79268),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_12_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_12_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__80107),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_12_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_12_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81075),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_12_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_12_11_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_12_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79888),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83861),
            .ce(N__47403),
            .sr(N__77286));
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47397),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83871),
            .ce(N__60725),
            .sr(N__77295));
    defparam \ppm_encoder_1.rudder_esr_5_LC_12_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_12_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47379),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83871),
            .ce(N__60725),
            .sr(N__77295));
    defparam \pid_front.state_1_LC_12_13_0 .C_ON=1'b0;
    defparam \pid_front.state_1_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_1_LC_12_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.state_1_LC_12_13_0  (
            .in0(N__52194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83882),
            .ce(),
            .sr(N__77304));
    defparam \pid_front.state_RNI26LH_0_LC_12_13_1 .C_ON=1'b0;
    defparam \pid_front.state_RNI26LH_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI26LH_0_LC_12_13_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_RNI26LH_0_LC_12_13_1  (
            .in0(N__52080),
            .in1(N__67367),
            .in2(_gnd_net_),
            .in3(N__52193),
            .lcout(\pid_front.state_ns_0 ),
            .ltout(\pid_front.state_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIVIRQ_0_0_LC_12_13_2 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_0_LC_12_13_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.state_RNIVIRQ_0_0_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47367),
            .in3(N__77601),
            .lcout(\pid_front.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIEI7TH_1_LC_12_13_3 .C_ON=1'b0;
    defparam \pid_front.state_RNIEI7TH_1_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIEI7TH_1_LC_12_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNIEI7TH_1_LC_12_13_3  (
            .in0(N__52081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47362),
            .lcout(\pid_front.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_1_LC_12_13_5 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50073),
            .lcout(\pid_alt.N_76_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83882),
            .ce(),
            .sr(N__77304));
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_14_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_14_0  (
            .in0(N__47568),
            .in1(N__47557),
            .in2(N__49287),
            .in3(N__47507),
            .lcout(\pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_14_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_14_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_14_1  (
            .in0(N__47499),
            .in1(N__47484),
            .in2(_gnd_net_),
            .in3(N__75827),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ),
            .ltout(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_14_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_14_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__47508),
            .in2(N__47562),
            .in3(N__47558),
            .lcout(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_14_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_14_3  (
            .in0(N__47474),
            .in1(N__47462),
            .in2(_gnd_net_),
            .in3(N__75685),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_14_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_2_LC_12_14_4  (
            .in0(N__75828),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83893),
            .ce(N__52572),
            .sr(N__52467));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_14_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_14_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_14_5  (
            .in0(N__47498),
            .in1(N__47483),
            .in2(_gnd_net_),
            .in3(N__75826),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_14_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_3_LC_12_14_6  (
            .in0(N__75687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83893),
            .ce(N__52572),
            .sr(N__52467));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_14_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_14_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_14_7  (
            .in0(N__47475),
            .in1(N__47463),
            .in2(_gnd_net_),
            .in3(N__75686),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_12_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_12_15_0 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_12_15_0  (
            .in0(N__48108),
            .in1(N__47868),
            .in2(N__47931),
            .in3(N__47918),
            .lcout(\pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_12_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_12_15_1 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_12_15_1  (
            .in0(N__75792),
            .in1(N__48087),
            .in2(N__51792),
            .in3(N__51771),
            .lcout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ),
            .ltout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_12_15_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_12_15_2  (
            .in0(N__47885),
            .in1(N__47867),
            .in2(N__47922),
            .in3(N__47917),
            .lcout(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_12_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_12_15_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_12_15_3  (
            .in0(N__47805),
            .in1(N__47811),
            .in2(_gnd_net_),
            .in3(N__47765),
            .lcout(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_12_15_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_12_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__51788),
            .in2(_gnd_net_),
            .in3(N__75791),
            .lcout(\pid_front.N_1680_i ),
            .ltout(\pid_front.N_1680_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_12_15_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_12_15_5 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_9_LC_12_15_5  (
            .in0(N__47858),
            .in1(N__47837),
            .in2(N__47871),
            .in3(N__82307),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_12_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_12_15_6 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_12_15_6  (
            .in0(N__82308),
            .in1(N__47859),
            .in2(N__47841),
            .in3(N__47817),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ),
            .ltout(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_12_15_7  (
            .in0(N__47804),
            .in1(N__47790),
            .in2(N__47769),
            .in3(N__47764),
            .lcout(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_12_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_12_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIVGCQ_12_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__48369),
            .in2(_gnd_net_),
            .in3(N__48340),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_12_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_12_16_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNISTI31_12_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48156),
            .in3(N__77603),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_7_LC_12_16_4 .C_ON=1'b0;
    defparam \pid_front.error_axb_7_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_7_LC_12_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_axb_7_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__48152),
            .in2(_gnd_net_),
            .in3(N__48126),
            .lcout(\pid_front.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_12_16_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_12_16_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__51892),
            .in2(_gnd_net_),
            .in3(N__51805),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_12_16_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_12_16_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_12_16_6  (
            .in0(N__51806),
            .in1(_gnd_net_),
            .in2(N__51899),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_12_16_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_12_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__51833),
            .in2(_gnd_net_),
            .in3(N__78830),
            .lcout(\pid_front.N_1686_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI4CD85_12_LC_12_17_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4CD85_12_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4CD85_12_LC_12_17_0 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4CD85_12_LC_12_17_0  (
            .in0(N__51609),
            .in1(N__78771),
            .in2(_gnd_net_),
            .in3(N__48081),
            .lcout(),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI4CD85Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIKI4D7_12_LC_12_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIKI4D7_12_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIKI4D7_12_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIKI4D7_12_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__48055),
            .in2(N__48024),
            .in3(N__48021),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIKI4D7Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQTN5D_13_LC_12_17_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQTN5D_13_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQTN5D_13_LC_12_17_2 .LUT_INIT=16'b1111110011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQTN5D_13_LC_12_17_2  (
            .in0(N__47979),
            .in1(N__47967),
            .in2(N__48846),
            .in3(N__47949),
            .lcout(\pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13 ),
            .ltout(\pid_front.error_p_reg_esr_RNIQTN5DZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3TJH01_13_LC_12_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3TJH01_13_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3TJH01_13_LC_12_17_3 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3TJH01_13_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__48427),
            .in2(N__48528),
            .in3(N__48525),
            .lcout(\pid_front.error_p_reg_esr_RNI3TJH01Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI5HTGG_13_LC_12_17_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI5HTGG_13_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI5HTGG_13_LC_12_17_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI5HTGG_13_LC_12_17_4  (
            .in0(N__48428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48491),
            .lcout(\pid_front.error_p_reg_esr_RNI5HTGGZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_12_17_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_12_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_12_17_5  (
            .in0(N__48471),
            .in1(N__52032),
            .in2(_gnd_net_),
            .in3(N__48455),
            .lcout(\pid_front.un1_pid_prereg_0_0 ),
            .ltout(\pid_front.un1_pid_prereg_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI31A7N_13_LC_12_17_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI31A7N_13_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI31A7N_13_LC_12_17_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI31A7N_13_LC_12_17_6  (
            .in0(N__48429),
            .in1(N__48492),
            .in2(N__48483),
            .in3(N__48776),
            .lcout(\pid_front.error_p_reg_esr_RNI31A7NZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_12_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_12_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_12_17_7  (
            .in0(N__48470),
            .in1(N__52031),
            .in2(_gnd_net_),
            .in3(N__48454),
            .lcout(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_12_18_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_12_18_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_12_18_0  (
            .in0(N__48416),
            .in1(N__48395),
            .in2(_gnd_net_),
            .in3(N__84433),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_19_LC_12_18_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_12_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_19_LC_12_18_1  (
            .in0(N__84435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83940),
            .ce(N__52569),
            .sr(N__52445));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_12_18_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_12_18_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_19_LC_12_18_2  (
            .in0(N__48417),
            .in1(N__48396),
            .in2(_gnd_net_),
            .in3(N__84434),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_12_18_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_12_18_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_12_18_3  (
            .in0(N__75732),
            .in1(N__48924),
            .in2(_gnd_net_),
            .in3(N__48903),
            .lcout(\pid_front.error_p_reg_esr_RNI8NB61_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_12_18_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_12_18_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_13_LC_12_18_4  (
            .in0(N__48882),
            .in1(N__48830),
            .in2(_gnd_net_),
            .in3(N__78698),
            .lcout(\pid_front.error_p_reg_esr_RNIETB61Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_13_LC_12_18_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_12_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_13_LC_12_18_5  (
            .in0(N__78699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83940),
            .ce(N__52569),
            .sr(N__52445));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_12_18_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_12_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_12_18_6  (
            .in0(N__48816),
            .in1(N__51986),
            .in2(_gnd_net_),
            .in3(N__52685),
            .lcout(\pid_front.un1_pid_prereg_0_1 ),
            .ltout(\pid_front.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_12_18_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_12_18_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48765),
            .in3(N__48755),
            .lcout(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_12_19_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_12_19_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_12_19_0  (
            .in0(N__48628),
            .in1(N__84296),
            .in2(N__49146),
            .in3(N__48655),
            .lcout(\pid_front.un1_pid_prereg_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_12_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_12_19_1 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_12_19_1  (
            .in0(N__84295),
            .in1(N__48629),
            .in2(N__49145),
            .in3(N__48732),
            .lcout(\pid_front.un1_pid_prereg_0_20 ),
            .ltout(\pid_front.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_12_19_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_12_19_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_12_19_2  (
            .in0(N__49247),
            .in1(N__48705),
            .in2(N__48684),
            .in3(N__48681),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_12_19_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_12_19_3 .LUT_INIT=16'b1010100011101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_12_19_3  (
            .in0(N__48656),
            .in1(N__48630),
            .in2(N__84303),
            .in3(N__49122),
            .lcout(\pid_front.un1_pid_prereg_0_22 ),
            .ltout(\pid_front.un1_pid_prereg_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_12_19_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_12_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_12_19_4  (
            .in0(N__49233),
            .in1(N__49248),
            .in2(N__49257),
            .in3(N__49192),
            .lcout(\pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_12_19_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_12_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__49246),
            .in2(_gnd_net_),
            .in3(N__49232),
            .lcout(\pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_12_19_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_12_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__49208),
            .in2(_gnd_net_),
            .in3(N__49193),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_22_LC_12_19_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_22_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_22_LC_12_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_22_LC_12_19_7  (
            .in0(N__84300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83954),
            .ce(N__52543),
            .sr(N__52446));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_20_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_20_0 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_20_0  (
            .in0(N__82259),
            .in1(_gnd_net_),
            .in2(N__49395),
            .in3(N__49434),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ),
            .ltout(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_20_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_20_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__49379),
            .in2(N__49062),
            .in3(N__49055),
            .lcout(\pid_front.un1_pid_prereg_0_6 ),
            .ltout(\pid_front.un1_pid_prereg_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_20_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_20_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_20_2  (
            .in0(N__49032),
            .in1(N__49014),
            .in2(N__48996),
            .in3(N__48935),
            .lcout(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_20_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_20_3  (
            .in0(N__52595),
            .in1(N__48981),
            .in2(_gnd_net_),
            .in3(N__48959),
            .lcout(\pid_front.un1_pid_prereg_0_7 ),
            .ltout(\pid_front.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_20_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_20_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49464),
            .in3(N__49460),
            .lcout(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_20_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_20_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_20_5  (
            .in0(N__49433),
            .in1(N__49391),
            .in2(_gnd_net_),
            .in3(N__82258),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_20_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_20_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_17_LC_12_20_6  (
            .in0(N__82260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83967),
            .ce(N__52558),
            .sr(N__52465));
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_20_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_20_7  (
            .in0(N__52583),
            .in1(N__52622),
            .in2(_gnd_net_),
            .in3(N__82228),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_21_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_21_0 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_21_0  (
            .in0(N__52945),
            .in1(N__52998),
            .in2(N__52299),
            .in3(N__52899),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_21_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_21_1  (
            .in0(N__52315),
            .in1(_gnd_net_),
            .in2(N__49365),
            .in3(N__49263),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_21_2  (
            .in0(N__49362),
            .in1(N__49307),
            .in2(N__49323),
            .in3(N__49482),
            .lcout(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_21_3 .LUT_INIT=16'b1110111110001010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_21_3  (
            .in0(N__49308),
            .in1(N__53006),
            .in2(N__52320),
            .in3(N__49293),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_21_4 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_21_4  (
            .in0(N__52944),
            .in1(N__52997),
            .in2(N__52298),
            .in3(N__52898),
            .lcout(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_21_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_0_LC_12_21_5  (
            .in0(N__52900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83983),
            .ce(N__52570),
            .sr(N__52466));
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_21_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__52314),
            .in2(_gnd_net_),
            .in3(N__52999),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_1_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53007),
            .lcout(\pid_front.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83983),
            .ce(N__52570),
            .sr(N__52466));
    defparam \dron_frame_decoder_1.source_H_disp_front_0_LC_12_22_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_0_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_0_LC_12_22_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_0_LC_12_22_0  (
            .in0(N__53310),
            .in1(N__61810),
            .in2(N__72072),
            .in3(N__53200),
            .lcout(drone_H_disp_front_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84001),
            .ce(),
            .sr(N__77363));
    defparam \pid_front.error_i_reg_esr_RNO_10_21_LC_12_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_10_21_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_10_21_LC_12_22_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_10_21_LC_12_22_1  (
            .in0(N__61809),
            .in1(N__71584),
            .in2(_gnd_net_),
            .in3(N__49616),
            .lcout(),
            .ltout(\pid_front.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_6_21_LC_12_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_6_21_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_6_21_LC_12_22_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_6_21_LC_12_22_2  (
            .in0(N__61674),
            .in1(_gnd_net_),
            .in2(N__49476),
            .in3(N__73580),
            .lcout(\pid_front.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_8_LC_12_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_8_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_8_LC_12_22_3 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_8_LC_12_22_3  (
            .in0(N__49473),
            .in1(N__53311),
            .in2(N__53210),
            .in3(N__72071),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84001),
            .ce(),
            .sr(N__77363));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIFDVA_8_LC_12_22_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIFDVA_8_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIFDVA_8_LC_12_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIFDVA_8_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49472),
            .lcout(drone_H_disp_front_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_0_LC_12_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_0_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_0_LC_12_22_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_fast_0_LC_12_22_5  (
            .in0(N__53315),
            .in1(N__72070),
            .in2(N__53211),
            .in3(N__49674),
            .lcout(dron_frame_decoder_1_source_H_disp_front_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84001),
            .ce(),
            .sr(N__77363));
    defparam \dron_frame_decoder_1.source_H_disp_front_2_LC_12_22_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_2_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_2_LC_12_22_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_2_LC_12_22_6  (
            .in0(N__49683),
            .in1(N__53201),
            .in2(N__53325),
            .in3(N__71837),
            .lcout(drone_H_disp_front_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84001),
            .ce(),
            .sr(N__77363));
    defparam \pid_front.error_axb_2_LC_12_22_7 .C_ON=1'b0;
    defparam \pid_front.error_axb_2_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_2_LC_12_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_2_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49682),
            .lcout(\pid_front.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_inv_LC_12_23_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_inv_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_inv_LC_12_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_cry_0_c_inv_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__49662),
            .in2(_gnd_net_),
            .in3(N__49673),
            .lcout(\pid_front.error_axb_0 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\pid_front.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNI39KI_LC_12_23_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_RNI39KI_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI39KI_LC_12_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_0_c_RNI39KI_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__49656),
            .in2(_gnd_net_),
            .in3(N__49578),
            .lcout(\pid_front.error_1 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0 ),
            .carryout(\pid_front.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI5CLI_LC_12_23_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_c_RNI5CLI_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI5CLI_LC_12_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_1_c_RNI5CLI_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__49575),
            .in2(_gnd_net_),
            .in3(N__49569),
            .lcout(\pid_front.error_2 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1 ),
            .carryout(\pid_front.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNI7FMI_LC_12_23_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_c_RNI7FMI_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNI7FMI_LC_12_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_2_c_RNI7FMI_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__49566),
            .in2(_gnd_net_),
            .in3(N__49557),
            .lcout(\pid_front.error_3 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2 ),
            .carryout(\pid_front.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNI1DAN_LC_12_23_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_c_RNI1DAN_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNI1DAN_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_c_RNI1DAN_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__49554),
            .in2(N__49545),
            .in3(N__49527),
            .lcout(\pid_front.error_4 ),
            .ltout(),
            .carryin(\pid_front.error_cry_3 ),
            .carryout(\pid_front.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIFSKI_LC_12_23_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_0_c_RNIFSKI_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIFSKI_LC_12_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIFSKI_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__53409),
            .in2(N__49524),
            .in3(N__49506),
            .lcout(\pid_front.error_5 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0_0 ),
            .carryout(\pid_front.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNII2RM_LC_12_23_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_0_c_RNII2RM_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNII2RM_LC_12_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNII2RM_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__53394),
            .in2(N__49503),
            .in3(N__49485),
            .lcout(\pid_front.error_6 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1_0 ),
            .carryout(\pid_front.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIL81R_LC_12_23_7 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_0_c_RNIL81R_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIL81R_LC_12_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIL81R_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__52698),
            .in2(N__49875),
            .in3(N__49857),
            .lcout(\pid_front.error_7 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2_0 ),
            .carryout(\pid_front.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIOE7V_LC_12_24_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_0_c_RNIOE7V_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIOE7V_LC_12_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIOE7V_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__49854),
            .in2(N__49845),
            .in3(N__49830),
            .lcout(\pid_front.error_8 ),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\pid_front.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_24_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_12_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_4_c_RNILNBG_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(N__49827),
            .in2(N__49809),
            .in3(N__49791),
            .lcout(\pid_front.error_9 ),
            .ltout(),
            .carryin(\pid_front.error_cry_4 ),
            .carryout(\pid_front.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIMGHM_LC_12_24_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_5_c_RNIMGHM_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIMGHM_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_5_c_RNIMGHM_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__53130),
            .in2(N__49788),
            .in3(N__49770),
            .lcout(\pid_front.error_10 ),
            .ltout(),
            .carryin(\pid_front.error_cry_5 ),
            .carryout(\pid_front.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_24_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_12_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_6_c_RNI3VJG_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__49767),
            .in2(_gnd_net_),
            .in3(N__49755),
            .lcout(\pid_front.error_11 ),
            .ltout(),
            .carryin(\pid_front.error_cry_6 ),
            .carryout(\pid_front.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_24_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_12_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_7_c_RNIAPPM_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__49752),
            .in2(N__49737),
            .in3(N__49701),
            .lcout(\pid_front.error_12 ),
            .ltout(),
            .carryin(\pid_front.error_cry_7 ),
            .carryout(\pid_front.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNI154L_LC_12_24_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_8_c_RNI154L_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNI154L_LC_12_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_8_c_RNI154L_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__49698),
            .in2(N__53445),
            .in3(N__49689),
            .lcout(\pid_front.error_13 ),
            .ltout(),
            .carryin(\pid_front.error_cry_8 ),
            .carryout(\pid_front.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIR17S_LC_12_24_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_9_c_RNIR17S_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIR17S_LC_12_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_9_c_RNIR17S_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__53424),
            .in2(N__53388),
            .in3(N__49686),
            .lcout(\pid_front.error_14 ),
            .ltout(),
            .carryin(\pid_front.error_cry_9 ),
            .carryout(\pid_front.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNI5FH01_LC_12_24_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNI5FH01_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNI5FH01_LC_12_24_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_cry_10_c_RNI5FH01_LC_12_24_7  (
            .in0(N__52728),
            .in1(N__53387),
            .in2(_gnd_net_),
            .in3(N__50001),
            .lcout(\pid_front.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNI1ADU1_LC_12_25_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNI1ADU1_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNI1ADU1_LC_12_25_0 .LUT_INIT=16'b1010111110111011;
    LogicCell40 \pid_front.error_cry_7_c_RNI1ADU1_LC_12_25_0  (
            .in0(N__72885),
            .in1(N__55710),
            .in2(N__55804),
            .in3(N__71462),
            .lcout(\pid_front.error_cry_7_c_RNI1ADUZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNI1ADU1_0_LC_12_25_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNI1ADU1_0_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNI1ADU1_0_LC_12_25_1 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \pid_front.error_cry_7_c_RNI1ADU1_0_LC_12_25_1  (
            .in0(N__71461),
            .in1(N__55784),
            .in2(N__55727),
            .in3(N__72884),
            .lcout(\pid_front.error_cry_7_c_RNI1ADU1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_12_25_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_12_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73771),
            .lcout(xy_ki_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84049),
            .ce(N__73402),
            .sr(N__77379));
    defparam \pid_front.error_i_reg_esr_RNO_11_21_LC_12_25_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_11_21_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_11_21_LC_12_25_3 .LUT_INIT=16'b0001100101011101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_11_21_LC_12_25_3  (
            .in0(N__71463),
            .in1(N__72886),
            .in2(N__49984),
            .in3(N__50196),
            .lcout(),
            .ltout(\pid_front.g0_11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_8_21_LC_12_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_8_21_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_8_21_LC_12_25_4 .LUT_INIT=16'b1011000010110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_8_21_LC_12_25_4  (
            .in0(N__72887),
            .in1(N__50355),
            .in2(N__49920),
            .in3(N__50133),
            .lcout(),
            .ltout(\pid_front.N_12_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_12_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_21_LC_12_25_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_21_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(N__61669),
            .in2(N__49917),
            .in3(N__49881),
            .lcout(),
            .ltout(\pid_front.N_116_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_12_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_12_25_6 .LUT_INIT=16'b0011000110111001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_21_LC_12_25_6  (
            .in0(N__69667),
            .in1(N__70453),
            .in2(N__49914),
            .in3(N__49911),
            .lcout(\pid_front.un4_error_i_reg_31_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_9_21_LC_12_25_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_9_21_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_9_21_LC_12_25_7 .LUT_INIT=16'b1010000110101011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_9_21_LC_12_25_7  (
            .in0(N__49887),
            .in1(N__53567),
            .in2(N__73307),
            .in3(N__53865),
            .lcout(\pid_front.N_89_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_12_26_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_12_26_0 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_26_LC_12_26_0  (
            .in0(N__69688),
            .in1(N__56504),
            .in2(N__69955),
            .in3(N__50250),
            .lcout(\pid_front.error_i_reg_9_rn_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_12_26_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_12_26_1 .LUT_INIT=16'b0000100000001101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_18_LC_12_26_1  (
            .in0(N__65747),
            .in1(N__59201),
            .in2(N__70515),
            .in3(N__56377),
            .lcout(),
            .ltout(\pid_front.m6_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_12_26_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_12_26_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_18_LC_12_26_2  (
            .in0(N__69933),
            .in1(N__69679),
            .in2(N__50373),
            .in3(N__56505),
            .lcout(\pid_front.error_i_reg_9_rn_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNII7HH1_LC_12_26_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNII7HH1_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNII7HH1_LC_12_26_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_0_0_c_RNII7HH1_LC_12_26_3  (
            .in0(N__71451),
            .in1(N__50353),
            .in2(_gnd_net_),
            .in3(N__50295),
            .lcout(\pid_front.N_27_1 ),
            .ltout(\pid_front.N_27_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIVCAK3_LC_12_26_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIVCAK3_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIVCAK3_LC_12_26_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIVCAK3_LC_12_26_4  (
            .in0(_gnd_net_),
            .in1(N__72907),
            .in2(N__50256),
            .in3(N__50087),
            .lcout(\pid_front.N_63 ),
            .ltout(\pid_front.N_63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIO7KH6_LC_12_26_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIO7KH6_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIO7KH6_LC_12_26_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIO7KH6_LC_12_26_5  (
            .in0(N__61664),
            .in1(_gnd_net_),
            .in2(N__50253),
            .in3(N__59200),
            .lcout(\pid_front.N_41_0 ),
            .ltout(\pid_front.N_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_10_LC_12_26_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_10_LC_12_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_10_LC_12_26_6 .LUT_INIT=16'b1100000001000100;
    LogicCell40 \pid_front.error_i_reg_esr_10_LC_12_26_6  (
            .in0(N__53697),
            .in1(N__65459),
            .in2(N__50244),
            .in3(N__70466),
            .lcout(\pid_front.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84066),
            .ce(N__59327),
            .sr(N__77384));
    defparam \pid_front.error_cry_3_c_RNIASQJ1_LC_12_26_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_c_RNIASQJ1_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNIASQJ1_LC_12_26_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_3_c_RNIASQJ1_LC_12_26_7  (
            .in0(N__72664),
            .in1(N__50194),
            .in2(_gnd_net_),
            .in3(N__50131),
            .lcout(\pid_front.N_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIH1EN_0_LC_12_30_2 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_30_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_30_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_12_30_2  (
            .in0(_gnd_net_),
            .in1(N__50072),
            .in2(_gnd_net_),
            .in3(N__77606),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_13_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_13_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_13_2_2  (
            .in0(N__54025),
            .in1(N__53947),
            .in2(N__54006),
            .in3(N__53974),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_13_LC_13_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_13_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_13_LC_13_2_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_13_LC_13_2_3  (
            .in0(N__66307),
            .in1(N__50421),
            .in2(N__50424),
            .in3(N__54244),
            .lcout(\ppm_encoder_1.N_139_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIV5A8_8_LC_13_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIV5A8_8_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIV5A8_8_LC_13_2_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIV5A8_8_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(N__54208),
            .in2(_gnd_net_),
            .in3(N__54586),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_13_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_13_3_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_13_3_0  (
            .in0(N__56274),
            .in1(N__50381),
            .in2(N__50412),
            .in3(N__50399),
            .lcout(\ppm_encoder_1.N_232 ),
            .ltout(\ppm_encoder_1.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_3_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_3_1  (
            .in0(N__56721),
            .in1(N__54972),
            .in2(N__50415),
            .in3(N__56265),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_13_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_13_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_13_3_3  (
            .in0(N__66346),
            .in1(N__62365),
            .in2(N__62391),
            .in3(N__56684),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_13_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_13_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_13_3_4  (
            .in0(N__56217),
            .in1(N__50382),
            .in2(N__50403),
            .in3(N__50400),
            .lcout(\ppm_encoder_1.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_13_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_13_3_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_13_3_6  (
            .in0(N__54633),
            .in1(N__53911),
            .in2(N__54107),
            .in3(N__56606),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_13_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_13_4_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_13_4_2  (
            .in0(N__53952),
            .in1(N__50505),
            .in2(N__50499),
            .in3(N__53976),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_13_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_13_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_13_4_6  (
            .in0(N__74759),
            .in1(N__66744),
            .in2(_gnd_net_),
            .in3(N__51018),
            .lcout(),
            .ltout(\ppm_encoder_1.N_313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_13_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_13_4_7 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_13_4_7  (
            .in0(_gnd_net_),
            .in1(N__56808),
            .in2(N__50508),
            .in3(N__74873),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_13_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_13_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_13_5_1  (
            .in0(N__78186),
            .in1(N__57219),
            .in2(_gnd_net_),
            .in3(N__50550),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83817),
            .ce(N__65866),
            .sr(N__77254));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_13_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_13_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_13_5_2  (
            .in0(N__78183),
            .in1(N__56976),
            .in2(_gnd_net_),
            .in3(N__66189),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83817),
            .ce(N__65866),
            .sr(N__77254));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_13_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_13_5_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_13_5_3  (
            .in0(N__59811),
            .in1(N__78184),
            .in2(_gnd_net_),
            .in3(N__54123),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83817),
            .ce(N__65866),
            .sr(N__77254));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_13_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_13_5_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_13_5_4  (
            .in0(N__53913),
            .in1(N__50478),
            .in2(N__54108),
            .in3(N__50490),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_13_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_13_5_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_13_5_5  (
            .in0(N__50787),
            .in1(N__78185),
            .in2(_gnd_net_),
            .in3(N__50484),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83817),
            .ce(N__65866),
            .sr(N__77254));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_13_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_13_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_13_5_6  (
            .in0(N__78182),
            .in1(N__54759),
            .in2(_gnd_net_),
            .in3(N__54114),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83817),
            .ce(N__65866),
            .sr(N__77254));
    defparam \ppm_encoder_1.rudder_10_LC_13_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_13_6_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_13_6_1  (
            .in0(N__50472),
            .in1(N__50466),
            .in2(N__62712),
            .in3(N__59980),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83820),
            .ce(),
            .sr(N__77261));
    defparam \ppm_encoder_1.rudder_13_LC_13_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_13_6_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_13_6_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_13_6_3  (
            .in0(N__50448),
            .in1(N__50430),
            .in2(N__62713),
            .in3(N__57052),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83820),
            .ce(),
            .sr(N__77261));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_13_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_13_6_4 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_13_6_4  (
            .in0(N__74855),
            .in1(N__76323),
            .in2(N__74766),
            .in3(N__54342),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_6_5 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_6_5  (
            .in0(N__74748),
            .in1(N__73878),
            .in2(N__50595),
            .in3(N__74856),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_7_LC_13_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_13_6_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_13_6_6  (
            .in0(N__50593),
            .in1(N__50544),
            .in2(N__62714),
            .in3(N__50538),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83820),
            .ce(),
            .sr(N__77261));
    defparam \ppm_encoder_1.aileron_1_LC_13_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_1_LC_13_6_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_1_LC_13_6_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_1_LC_13_6_7  (
            .in0(N__59760),
            .in1(N__66912),
            .in2(N__62711),
            .in3(N__57100),
            .lcout(\ppm_encoder_1.aileronZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83820),
            .ce(),
            .sr(N__77261));
    defparam \ppm_encoder_1.throttle_RNIB03T2_6_LC_13_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIB03T2_6_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIB03T2_6_LC_13_7_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIB03T2_6_LC_13_7_0  (
            .in0(N__66149),
            .in1(N__59935),
            .in2(N__50610),
            .in3(N__63250),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI1T1M6_6_LC_13_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI1T1M6_6_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI1T1M6_6_LC_13_7_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNI1T1M6_6_LC_13_7_1  (
            .in0(N__66168),
            .in1(_gnd_net_),
            .in2(N__50520),
            .in3(N__50517),
            .lcout(\ppm_encoder_1.throttle_RNI1T1M6Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_13_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_13_7_2 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNIAH7O2_6_LC_13_7_2  (
            .in0(N__50686),
            .in1(N__63148),
            .in2(N__50676),
            .in3(N__63327),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_13_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_13_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_13_7_3  (
            .in0(N__63504),
            .in1(N__50608),
            .in2(_gnd_net_),
            .in3(N__50674),
            .lcout(),
            .ltout(\ppm_encoder_1.N_292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_13_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_13_7_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_13_7_4  (
            .in0(N__50687),
            .in1(_gnd_net_),
            .in2(N__50511),
            .in3(N__63044),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_13_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_13_7_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_13_7_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_13_7_5  (
            .in0(N__60120),
            .in1(N__50688),
            .in2(N__60147),
            .in3(N__62671),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83823),
            .ce(),
            .sr(N__77270));
    defparam \ppm_encoder_1.elevator_6_LC_13_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_13_7_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_13_7_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_13_7_6  (
            .in0(N__50675),
            .in1(N__51135),
            .in2(N__62715),
            .in3(N__51159),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83823),
            .ce(),
            .sr(N__77270));
    defparam \ppm_encoder_1.throttle_6_LC_13_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_13_7_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_13_7_7 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_13_7_7  (
            .in0(N__50661),
            .in1(N__50609),
            .in2(N__50652),
            .in3(N__62672),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83823),
            .ce(),
            .sr(N__77270));
    defparam \ppm_encoder_1.throttle_RNID23T2_7_LC_13_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNID23T2_7_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNID23T2_7_LC_13_8_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNID23T2_7_LC_13_8_0  (
            .in0(N__50594),
            .in1(N__59951),
            .in2(N__54187),
            .in3(N__63265),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI622M6_7_LC_13_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI622M6_7_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI622M6_7_LC_13_8_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNI622M6_7_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__63534),
            .in2(N__50571),
            .in3(N__50568),
            .lcout(\ppm_encoder_1.throttle_RNI622M6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_13_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_13_8_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNICJ7O2_7_LC_13_8_2  (
            .in0(N__50560),
            .in1(N__63163),
            .in2(N__54160),
            .in3(N__63364),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_13_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_13_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_13_8_4  (
            .in0(N__50561),
            .in1(N__63045),
            .in2(_gnd_net_),
            .in3(N__54135),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_13_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_13_8_5 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_13_8_5  (
            .in0(N__60078),
            .in1(N__50562),
            .in2(N__60105),
            .in3(N__62678),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83828),
            .ce(),
            .sr(N__77274));
    defparam \ppm_encoder_1.elevator_7_LC_13_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_13_8_6 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_13_8_6  (
            .in0(N__62676),
            .in1(N__54162),
            .in2(N__51099),
            .in3(N__51123),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83828),
            .ce(),
            .sr(N__77274));
    defparam \ppm_encoder_1.throttle_7_LC_13_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_13_8_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_13_8_7  (
            .in0(N__50838),
            .in1(N__50805),
            .in2(N__54189),
            .in3(N__62677),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83828),
            .ce(),
            .sr(N__77274));
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_13_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_13_9_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI24LH2_11_LC_13_9_0  (
            .in0(N__50773),
            .in1(N__63164),
            .in2(N__50760),
            .in3(N__63362),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIT4BA6_11_LC_13_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIT4BA6_11_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIT4BA6_11_LC_13_9_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIT4BA6_11_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__66768),
            .in2(N__50799),
            .in3(N__50796),
            .lcout(\ppm_encoder_1.elevator_RNIT4BA6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI332R2_11_LC_13_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI332R2_11_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI332R2_11_LC_13_9_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNI332R2_11_LC_13_9_2  (
            .in0(N__51013),
            .in1(N__59934),
            .in2(N__50708),
            .in3(N__63266),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_13_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_13_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_13_9_3  (
            .in0(N__63490),
            .in1(N__50704),
            .in2(_gnd_net_),
            .in3(N__50758),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_9_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_9_4  (
            .in0(N__50774),
            .in1(_gnd_net_),
            .in2(N__50790),
            .in3(N__63046),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_13_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_13_9_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_13_9_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_13_9_5  (
            .in0(N__60804),
            .in1(N__60783),
            .in2(N__50778),
            .in3(N__62682),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83833),
            .ce(),
            .sr(N__77279));
    defparam \ppm_encoder_1.elevator_11_LC_13_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_13_9_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_13_9_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_13_9_6  (
            .in0(N__50759),
            .in1(N__51354),
            .in2(N__62716),
            .in3(N__51333),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83833),
            .ce(),
            .sr(N__77279));
    defparam \ppm_encoder_1.throttle_11_LC_13_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_13_9_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_13_9_7  (
            .in0(N__50745),
            .in1(N__50715),
            .in2(N__50709),
            .in3(N__62683),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83833),
            .ce(),
            .sr(N__77279));
    defparam \ppm_encoder_1.elevator_9_LC_13_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_13_10_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_13_10_0  (
            .in0(N__51081),
            .in1(N__51057),
            .in2(N__54558),
            .in3(N__62568),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.rudder_11_LC_13_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_13_10_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_13_10_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_13_10_1  (
            .in0(N__51045),
            .in1(N__51027),
            .in2(N__62653),
            .in3(N__51017),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_13_10_2  (
            .in0(N__50997),
            .in1(N__62558),
            .in2(N__50988),
            .in3(N__54533),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_13_10_3  (
            .in0(N__50967),
            .in1(N__50949),
            .in2(N__62654),
            .in3(N__74030),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.rudder_9_LC_13_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_13_10_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_13_10_4  (
            .in0(N__50937),
            .in1(N__50928),
            .in2(N__56951),
            .in3(N__62569),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.throttle_1_LC_13_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_13_10_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_13_10_5  (
            .in0(N__50910),
            .in1(N__50903),
            .in2(N__62655),
            .in3(N__59056),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.throttle_10_LC_13_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_13_10_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_13_10_6  (
            .in0(N__50877),
            .in1(N__50847),
            .in2(N__59867),
            .in3(N__62570),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83841),
            .ce(),
            .sr(N__77287));
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_c_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__59558),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__57185),
            .in2(N__60447),
            .in3(N__50841),
            .lcout(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_0 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__62879),
            .in2(_gnd_net_),
            .in3(N__51171),
            .lcout(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_1 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__59711),
            .in2(N__60448),
            .in3(N__51168),
            .lcout(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_2 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__57440),
            .in2(_gnd_net_),
            .in3(N__51165),
            .lcout(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_3 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__57413),
            .in2(_gnd_net_),
            .in3(N__51162),
            .lcout(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_4 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_11_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__51155),
            .in2(N__60449),
            .in3(N__51126),
            .lcout(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_5 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_11_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__51122),
            .in2(_gnd_net_),
            .in3(N__51087),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_12_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__54452),
            .in2(_gnd_net_),
            .in3(N__51084),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_12_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__51074),
            .in2(_gnd_net_),
            .in3(N__51048),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_12_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__57482),
            .in2(_gnd_net_),
            .in3(N__51357),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_12_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__51350),
            .in2(_gnd_net_),
            .in3(N__51324),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_12_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__54719),
            .in2(_gnd_net_),
            .in3(N__51321),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_12_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__57335),
            .in2(N__60520),
            .in3(N__51318),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51315),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83859),
            .ce(N__60726),
            .sr(N__77305));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_13_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_13_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__80504),
            .in2(_gnd_net_),
            .in3(N__83017),
            .lcout(xy_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_13_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_13_13_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_1_LC_13_13_1  (
            .in0(N__83018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73727),
            .lcout(xy_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_13_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_13_13_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_2_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__80249),
            .in2(_gnd_net_),
            .in3(N__83019),
            .lcout(xy_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_13_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_13_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_3_LC_13_13_3  (
            .in0(N__83020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79726),
            .lcout(xy_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_13_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_13_13_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__80106),
            .in2(_gnd_net_),
            .in3(N__83016),
            .lcout(xy_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_13_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_13_13_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_5_LC_13_13_5  (
            .in0(N__83021),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81081),
            .lcout(xy_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_13_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_13_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_6_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__79892),
            .in2(_gnd_net_),
            .in3(N__83022),
            .lcout(xy_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83869),
            .ce(N__51438),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_13_14_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_13_14_6 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_13_14_6  (
            .in0(N__51426),
            .in1(N__58304),
            .in2(N__51380),
            .in3(N__51417),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83879),
            .ce(),
            .sr(N__77321));
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_13_15_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_13_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_17_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67998),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_13_15_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_13_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_1_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68114),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_13_15_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_13_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_2_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75364),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_13_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_13_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_3_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60933),
            .lcout(\pid_side.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_13_15_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_13_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_4_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60825),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_15_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_13_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_5_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74996),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_6_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75076),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_13_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_12_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67932),
            .lcout(\pid_side.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83890),
            .ce(N__78352),
            .sr(N__77329));
    defparam \pid_front.error_d_reg_prev_esr_10_LC_13_16_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_10_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78831),
            .lcout(\pid_front.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83900),
            .ce(N__52559),
            .sr(N__52461));
    defparam \pid_front.error_d_reg_prev_esr_12_LC_13_16_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_13_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_12_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78765),
            .lcout(\pid_front.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83900),
            .ce(N__52559),
            .sr(N__52461));
    defparam \pid_front.error_d_reg_prev_esr_20_LC_13_16_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_20_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84399),
            .lcout(\pid_front.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83900),
            .ce(N__52559),
            .sr(N__52461));
    defparam \pid_front.error_d_reg_prev_esr_21_LC_13_16_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_13_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_21_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84351),
            .lcout(\pid_front.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83900),
            .ce(N__52559),
            .sr(N__52461));
    defparam \pid_front.error_d_reg_prev_esr_9_LC_13_16_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_13_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_9_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75790),
            .lcout(\pid_front.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83900),
            .ce(N__52559),
            .sr(N__52461));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_13_17_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_13_17_0 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_13_17_0  (
            .in0(N__75784),
            .in1(N__51766),
            .in2(N__78829),
            .in3(N__51787),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_13_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_13_17_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__51828),
            .in2(N__51537),
            .in3(N__51744),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_13_17_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_13_17_2 .LUT_INIT=16'b1111110111010000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_13_17_2  (
            .in0(N__51832),
            .in1(N__78828),
            .in2(N__51972),
            .in3(N__51843),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJ35VF_12_LC_13_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJ35VF_12_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJ35VF_12_LC_13_17_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJ35VF_12_LC_13_17_3  (
            .in0(N__51939),
            .in1(N__51969),
            .in2(N__51957),
            .in3(N__51927),
            .lcout(\pid_front.error_p_reg_esr_RNIJ35VFZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQT424_12_LC_13_17_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQT424_12_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQT424_12_LC_13_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQT424_12_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__51938),
            .in2(_gnd_net_),
            .in3(N__51926),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINH0UD_10_LC_13_17_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINH0UD_10_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINH0UD_10_LC_13_17_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINH0UD_10_LC_13_17_5  (
            .in0(N__51900),
            .in1(N__51807),
            .in2(N__51864),
            .in3(N__51861),
            .lcout(\pid_front.error_d_reg_prev_esr_RNINH0UDZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_13_17_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_13_17_6 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_13_17_6  (
            .in0(N__78821),
            .in1(N__51842),
            .in2(N__51834),
            .in3(N__51813),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_13_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_13_17_7 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_10_LC_13_17_7  (
            .in0(N__51786),
            .in1(N__78817),
            .in2(N__51770),
            .in3(N__75783),
            .lcout(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIE0RO1_0_LC_13_18_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIE0RO1_0_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIE0RO1_0_LC_13_18_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_front.state_RNIE0RO1_0_LC_13_18_0  (
            .in0(N__52196),
            .in1(N__52221),
            .in2(N__52209),
            .in3(N__67343),
            .lcout(),
            .ltout(\pid_front.N_196_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI4UFB2_0_LC_13_18_1 .C_ON=1'b0;
    defparam \pid_front.state_RNI4UFB2_0_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI4UFB2_0_LC_13_18_1 .LUT_INIT=16'b1111111101110010;
    LogicCell40 \pid_front.state_RNI4UFB2_0_LC_13_18_1  (
            .in0(N__52104),
            .in1(N__52197),
            .in2(N__51738),
            .in3(N__77591),
            .lcout(\pid_front.error_i_acumm_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_3_LC_13_18_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_3_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_3_LC_13_18_2 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \pid_front.error_i_acumm_3_LC_13_18_2  (
            .in0(N__51735),
            .in1(N__51714),
            .in2(N__55011),
            .in3(N__52105),
            .lcout(\pid_front.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83925),
            .ce(N__51640),
            .sr(_gnd_net_));
    defparam \pid_side.m153_e_5_LC_13_18_3 .C_ON=1'b0;
    defparam \pid_side.m153_e_5_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.m153_e_5_LC_13_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.m153_e_5_LC_13_18_3  (
            .in0(N__70359),
            .in1(N__73572),
            .in2(N__69602),
            .in3(N__71147),
            .lcout(pid_side_m153_e_5),
            .ltout(pid_side_m153_e_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIAHFQ1_0_LC_13_18_4 .C_ON=1'b0;
    defparam \pid_side.state_RNIAHFQ1_0_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIAHFQ1_0_LC_13_18_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_side.state_RNIAHFQ1_0_LC_13_18_4  (
            .in0(N__52205),
            .in1(N__67344),
            .in2(N__52215),
            .in3(N__67280),
            .lcout(),
            .ltout(\pid_side.N_196_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIOGDG2_0_LC_13_18_5 .C_ON=1'b0;
    defparam \pid_side.state_RNIOGDG2_0_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIOGDG2_0_LC_13_18_5 .LUT_INIT=16'b1111111101110100;
    LogicCell40 \pid_side.state_RNIOGDG2_0_LC_13_18_5  (
            .in0(N__67281),
            .in1(N__67139),
            .in2(N__52212),
            .in3(N__77592),
            .lcout(\pid_side.error_i_acumm_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m153_e_4_LC_13_18_6 .C_ON=1'b0;
    defparam \pid_side.m153_e_4_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.m153_e_4_LC_13_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.m153_e_4_LC_13_18_6  (
            .in0(N__57656),
            .in1(N__57680),
            .in2(N__57627),
            .in3(N__61637),
            .lcout(pid_side_m153_e_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIVIRQ_0_LC_13_18_7 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_LC_13_18_7 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_front.state_RNIVIRQ_0_LC_13_18_7  (
            .in0(N__67342),
            .in1(N__52195),
            .in2(N__52126),
            .in3(N__77590),
            .lcout(\pid_front.state_RNIVIRQZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_13_19_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_13_19_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_13_19_0  (
            .in0(N__52019),
            .in1(N__51998),
            .in2(_gnd_net_),
            .in3(N__84160),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_15_LC_13_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_13_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_15_LC_13_19_1  (
            .in0(N__84162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83938),
            .ce(N__52571),
            .sr(N__52447));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_13_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_13_19_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_15_LC_13_19_2  (
            .in0(N__52020),
            .in1(N__51999),
            .in2(_gnd_net_),
            .in3(N__84161),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_13_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_13_19_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_13_19_3  (
            .in0(N__52670),
            .in1(N__52649),
            .in2(_gnd_net_),
            .in3(N__84193),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_16_LC_13_19_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_13_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_16_LC_13_19_4  (
            .in0(N__84195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83938),
            .ce(N__52571),
            .sr(N__52447));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_13_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_13_19_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_16_LC_13_19_5  (
            .in0(N__52671),
            .in1(N__52650),
            .in2(_gnd_net_),
            .in3(N__84194),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_13_19_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_13_19_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_18_LC_13_19_6  (
            .in0(N__52626),
            .in1(N__52584),
            .in2(_gnd_net_),
            .in3(N__82229),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_18_LC_13_19_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_13_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_18_LC_13_19_7  (
            .in0(N__82230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83938),
            .ce(N__52571),
            .sr(N__52447));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_13_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79275),
            .lcout(side_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83952),
            .ce(N__65028),
            .sr(N__77357));
    defparam \pid_front.error_p_reg_esr_1_LC_13_21_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_1_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_1_LC_13_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_1_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52338),
            .lcout(\pid_front.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83966),
            .ce(N__83134),
            .sr(N__82858));
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_21_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIL1E8_1_LC_13_21_1  (
            .in0(N__52319),
            .in1(N__52297),
            .in2(_gnd_net_),
            .in3(N__53000),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_21_2 .LUT_INIT=16'b0000111111000011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_13_21_2  (
            .in0(N__52278),
            .in1(N__52947),
            .in2(N__52239),
            .in3(N__52902),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_1_LC_13_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_1_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_1_LC_13_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_1_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53025),
            .lcout(\pid_front.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83966),
            .ce(N__83134),
            .sr(N__82858));
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_13_21_4  (
            .in0(N__52977),
            .in1(N__52946),
            .in2(_gnd_net_),
            .in3(N__52901),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_0_LC_13_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_0_LC_13_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_0_LC_13_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_0_LC_13_21_7  (
            .in0(N__52914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83966),
            .ce(N__83134),
            .sr(N__82858));
    defparam \dron_frame_decoder_1.source_Altitude_15_LC_13_22_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_15_LC_13_22_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_15_LC_13_22_0 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_15_LC_13_22_0  (
            .in0(N__52839),
            .in1(N__65142),
            .in2(N__58518),
            .in3(N__52873),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83982),
            .ce(),
            .sr(N__77367));
    defparam \dron_frame_decoder_1.source_Altitude_7_LC_13_22_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_7_LC_13_22_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_7_LC_13_22_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_7_LC_13_22_1  (
            .in0(N__52757),
            .in1(N__52840),
            .in2(N__65148),
            .in3(N__58517),
            .lcout(drone_altitude_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83982),
            .ce(),
            .sr(N__77367));
    defparam \dron_frame_decoder_1.source_Altitude_RNIB343_7_LC_13_22_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_RNIB343_7_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_RNIB343_7_LC_13_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_RNIB343_7_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52756),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_15_LC_13_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_15_LC_13_22_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_15_LC_13_22_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_15_LC_13_22_3  (
            .in0(N__53304),
            .in1(N__65147),
            .in2(N__52727),
            .in3(N__53196),
            .lcout(drone_H_disp_front_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83982),
            .ce(),
            .sr(N__77367));
    defparam \dron_frame_decoder_1.source_H_disp_front_7_LC_13_22_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_7_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_7_LC_13_22_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_7_LC_13_22_4  (
            .in0(N__52707),
            .in1(N__53306),
            .in2(N__53209),
            .in3(N__65146),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83982),
            .ce(),
            .sr(N__77367));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIECVA_7_LC_13_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIECVA_7_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIECVA_7_LC_13_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIECVA_7_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52706),
            .lcout(drone_H_disp_front_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_10_LC_13_22_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_10_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_10_LC_13_22_6 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_10_LC_13_22_6  (
            .in0(N__53139),
            .in1(N__53305),
            .in2(N__53208),
            .in3(N__71838),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83982),
            .ce(),
            .sr(N__77367));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIO24A_10_LC_13_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIO24A_10_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIO24A_10_LC_13_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIO24A_10_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53138),
            .lcout(drone_H_disp_front_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIUOTV1_0_LC_13_23_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIUOTV1_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIUOTV1_0_LC_13_23_0 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \pid_front.error_cry_5_c_RNIUOTV1_0_LC_13_23_0  (
            .in0(N__72696),
            .in1(N__55788),
            .in2(N__72958),
            .in3(N__53802),
            .lcout(\pid_front.error_cry_5_c_RNIUOTV1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIUOTV1_LC_13_23_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIUOTV1_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIUOTV1_LC_13_23_1 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \pid_front.error_cry_5_c_RNIUOTV1_LC_13_23_1  (
            .in0(N__53803),
            .in1(N__72918),
            .in2(N__55805),
            .in3(N__72697),
            .lcout(),
            .ltout(\pid_front.error_cry_5_c_RNIUOTVZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIBO8P5_LC_13_23_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIBO8P5_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIBO8P5_LC_13_23_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_5_c_RNIBO8P5_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__53036),
            .in2(N__53121),
            .in3(N__53118),
            .lcout(\pid_front.N_49_0 ),
            .ltout(\pid_front.N_49_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_13_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_13_23_3 .LUT_INIT=16'b0001001110011011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_15_LC_13_23_3  (
            .in0(N__70469),
            .in1(N__66061),
            .in2(N__53088),
            .in3(N__55436),
            .lcout(),
            .ltout(\pid_front.m134_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_13_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_13_23_4 .LUT_INIT=16'b0000111000111110;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_15_LC_13_23_4  (
            .in0(N__53085),
            .in1(N__70470),
            .in2(N__53064),
            .in3(N__56473),
            .lcout(),
            .ltout(\pid_front.m19_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_15_LC_13_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_15_LC_13_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_15_LC_13_23_5 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_front.error_i_reg_esr_15_LC_13_23_5  (
            .in0(N__69695),
            .in1(N__69852),
            .in2(N__53061),
            .in3(N__55488),
            .lcout(\pid_front.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83999),
            .ce(N__59367),
            .sr(N__77374));
    defparam \pid_front.error_cry_4_c_RNIF6DP1_LC_13_23_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNIF6DP1_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNIF6DP1_LC_13_23_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_4_c_RNIF6DP1_LC_13_23_6  (
            .in0(N__72695),
            .in1(N__53566),
            .in2(_gnd_net_),
            .in3(N__53864),
            .lcout(\pid_front.N_48_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_13_LC_13_24_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_13_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_13_LC_13_24_0 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_13_LC_13_24_0  (
            .in0(N__53438),
            .in1(N__53307),
            .in2(N__53173),
            .in3(N__68638),
            .lcout(drone_H_disp_front_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84017),
            .ce(),
            .sr(N__77380));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIR54A_13_LC_13_24_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIR54A_13_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIR54A_13_LC_13_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIR54A_13_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53437),
            .lcout(drone_H_disp_front_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_5_LC_13_24_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_5_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_5_LC_13_24_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_5_LC_13_24_2  (
            .in0(N__53418),
            .in1(N__53308),
            .in2(N__53175),
            .in3(N__68639),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84017),
            .ce(),
            .sr(N__77380));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNICAVA_5_LC_13_24_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNICAVA_5_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNICAVA_5_LC_13_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNICAVA_5_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53417),
            .lcout(drone_H_disp_front_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_6_LC_13_24_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_6_LC_13_24_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_6_LC_13_24_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_6_LC_13_24_4  (
            .in0(N__53403),
            .in1(N__53309),
            .in2(N__53176),
            .in3(N__68562),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84017),
            .ce(),
            .sr(N__77380));
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIDBVA_6_LC_13_24_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIDBVA_6_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_RNIDBVA_6_LC_13_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_RNIDBVA_6_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53402),
            .lcout(drone_H_disp_front_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_14_LC_13_24_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_14_LC_13_24_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_14_LC_13_24_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_14_LC_13_24_6  (
            .in0(N__53303),
            .in1(N__68561),
            .in2(N__53174),
            .in3(N__53383),
            .lcout(drone_H_disp_front_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84017),
            .ce(),
            .sr(N__77380));
    defparam \dron_frame_decoder_1.state_RNI00RU_3_LC_13_24_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI00RU_3_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI00RU_3_LC_13_24_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI00RU_3_LC_13_24_7  (
            .in0(N__53367),
            .in1(N__53302),
            .in2(_gnd_net_),
            .in3(N__58350),
            .lcout(\dron_frame_decoder_1.N_122_mux_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_13_25_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_13_25_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_24_LC_13_25_0  (
            .in0(N__70459),
            .in1(N__58965),
            .in2(_gnd_net_),
            .in3(N__58949),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_1_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_24_LC_13_25_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_24_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_24_LC_13_25_1 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.error_i_reg_esr_24_LC_13_25_1  (
            .in0(N__69928),
            .in1(N__69696),
            .in2(N__53664),
            .in3(N__55920),
            .lcout(\pid_front.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84031),
            .ce(N__59403),
            .sr(N__77385));
    defparam \pid_front.error_cry_2_0_c_RNI198H2_0_LC_13_25_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI198H2_0_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI198H2_0_LC_13_25_2 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI198H2_0_LC_13_25_2  (
            .in0(N__71448),
            .in1(N__53503),
            .in2(N__72922),
            .in3(N__53558),
            .lcout(\pid_front.error_cry_2_0_c_RNI198H2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIU4PB5_LC_13_25_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNIU4PB5_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIU4PB5_LC_13_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_7_c_RNIU4PB5_LC_13_25_3  (
            .in0(N__53763),
            .in1(N__53646),
            .in2(_gnd_net_),
            .in3(N__53640),
            .lcout(\pid_front.N_22_0 ),
            .ltout(\pid_front.N_22_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI59S7C_LC_13_25_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI59S7C_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI59S7C_LC_13_25_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI59S7C_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__61639),
            .in2(N__53634),
            .in3(N__53612),
            .lcout(\pid_front.N_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI198H2_LC_13_25_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI198H2_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI198H2_LC_13_25_5 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI198H2_LC_13_25_5  (
            .in0(N__53559),
            .in1(N__72883),
            .in2(N__53515),
            .in3(N__71449),
            .lcout(),
            .ltout(\pid_front.error_cry_2_0_c_RNI198HZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIKP1K6_LC_13_25_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIKP1K6_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIKP1K6_LC_13_25_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIKP1K6_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__53631),
            .in2(N__53625),
            .in3(N__53622),
            .lcout(\pid_front.N_28_1 ),
            .ltout(\pid_front.N_28_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNID77CA_LC_13_25_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNID77CA_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNID77CA_LC_13_25_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNID77CA_LC_13_25_7  (
            .in0(N__61638),
            .in1(_gnd_net_),
            .in2(N__53601),
            .in3(N__58988),
            .lcout(\pid_front.N_60_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIUV922_LC_13_26_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIUV922_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIUV922_LC_13_26_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIUV922_LC_13_26_0  (
            .in0(N__71453),
            .in1(N__53572),
            .in2(_gnd_net_),
            .in3(N__53507),
            .lcout(\pid_front.N_25_0 ),
            .ltout(\pid_front.N_25_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI1C944_0_LC_13_26_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI1C944_0_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI1C944_0_LC_13_26_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI1C944_0_LC_13_26_1  (
            .in0(N__66040),
            .in1(N__72984),
            .in2(N__53448),
            .in3(N__53761),
            .lcout(\pid_front.error_cry_2_0_c_RNI1C944Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNISGUE1_LC_13_26_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNISGUE1_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNISGUE1_LC_13_26_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_4_c_RNISGUE1_LC_13_26_2  (
            .in0(N__71452),
            .in1(N__53872),
            .in2(_gnd_net_),
            .in3(N__53811),
            .lcout(\pid_front.N_21_1 ),
            .ltout(\pid_front.N_21_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIG4884_LC_13_26_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNIG4884_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIG4884_LC_13_26_3 .LUT_INIT=16'b0100010000111111;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIG4884_LC_13_26_3  (
            .in0(N__53747),
            .in1(N__61665),
            .in2(N__53766),
            .in3(N__72988),
            .lcout(\pid_front.m38_1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI1C944_LC_13_26_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI1C944_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI1C944_LC_13_26_4 .LUT_INIT=16'b1111111011001110;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI1C944_LC_13_26_4  (
            .in0(N__53762),
            .in1(N__66041),
            .in2(N__72998),
            .in3(N__53748),
            .lcout(\pid_front.error_cry_2_0_c_RNI1CZ0Z944 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIVMTQ7_LC_13_26_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNIVMTQ7_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIVMTQ7_LC_13_26_5 .LUT_INIT=16'b0011111000110010;
    LogicCell40 \pid_front.error_cry_7_c_RNIVMTQ7_LC_13_26_5  (
            .in0(N__55674),
            .in1(N__53739),
            .in2(N__61670),
            .in3(N__56033),
            .lcout(\pid_front.N_39_1 ),
            .ltout(\pid_front.N_39_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_18_LC_13_26_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_18_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_18_LC_13_26_6 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \pid_front.error_i_reg_esr_18_LC_13_26_6  (
            .in0(N__61910),
            .in1(_gnd_net_),
            .in2(N__53733),
            .in3(N__53730),
            .lcout(\pid_front.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84047),
            .ce(N__59363),
            .sr(N__77390));
    defparam \pid_front.error_i_reg_esr_26_LC_13_26_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_26_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_26_LC_13_26_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \pid_front.error_i_reg_esr_26_LC_13_26_7  (
            .in0(N__59224),
            .in1(N__53703),
            .in2(_gnd_net_),
            .in3(N__53696),
            .lcout(\pid_front.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84047),
            .ce(N__59363),
            .sr(N__77390));
    defparam \ppm_encoder_1.counter_0_LC_14_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_14_2_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_14_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(N__56607),
            .in2(N__55467),
            .in3(N__55466),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_2_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_1_LC_14_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_14_2_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_14_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(N__56625),
            .in2(_gnd_net_),
            .in3(N__53667),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_2_LC_14_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_14_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_14_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_14_2_2  (
            .in0(_gnd_net_),
            .in1(N__56187),
            .in2(_gnd_net_),
            .in3(N__53982),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_3_LC_14_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_14_2_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_14_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__56207),
            .in2(_gnd_net_),
            .in3(N__53979),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_4_LC_14_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_14_2_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_14_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__53975),
            .in2(_gnd_net_),
            .in3(N__53955),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_5_LC_14_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_14_2_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_14_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(N__53948),
            .in2(_gnd_net_),
            .in3(N__53928),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_6_LC_14_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_14_2_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_14_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(N__54026),
            .in2(_gnd_net_),
            .in3(N__53925),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_7_LC_14_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_14_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_14_2_7  (
            .in0(_gnd_net_),
            .in1(N__54004),
            .in2(_gnd_net_),
            .in3(N__53922),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__83815),
            .ce(),
            .sr(N__54053));
    defparam \ppm_encoder_1.counter_8_LC_14_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_14_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(N__54587),
            .in2(_gnd_net_),
            .in3(N__53919),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_3_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_9_LC_14_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_14_3_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_14_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(N__54631),
            .in2(_gnd_net_),
            .in3(N__53916),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_10_LC_14_3_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_14_3_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_14_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_14_3_2  (
            .in0(_gnd_net_),
            .in1(N__53912),
            .in2(_gnd_net_),
            .in3(N__53892),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_11_LC_14_3_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_14_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_14_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(N__54103),
            .in2(_gnd_net_),
            .in3(N__54081),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_12_LC_14_3_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_14_3_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_14_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_14_3_4  (
            .in0(_gnd_net_),
            .in1(N__54209),
            .in2(_gnd_net_),
            .in3(N__54078),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_13_LC_14_3_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_14_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_14_3_5  (
            .in0(_gnd_net_),
            .in1(N__54245),
            .in2(_gnd_net_),
            .in3(N__54075),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_14_LC_14_3_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_14_3_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_14_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(N__66308),
            .in2(_gnd_net_),
            .in3(N__54072),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_15_LC_14_3_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_14_3_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_14_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_14_3_7  (
            .in0(_gnd_net_),
            .in1(N__66347),
            .in2(_gnd_net_),
            .in3(N__54069),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__83816),
            .ce(),
            .sr(N__54041));
    defparam \ppm_encoder_1.counter_16_LC_14_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_14_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(N__62389),
            .in2(_gnd_net_),
            .in3(N__54066),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_4_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__83818),
            .ce(),
            .sr(N__54057));
    defparam \ppm_encoder_1.counter_17_LC_14_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_14_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(N__62366),
            .in2(_gnd_net_),
            .in3(N__54063),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__83818),
            .ce(),
            .sr(N__54057));
    defparam \ppm_encoder_1.counter_18_LC_14_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_14_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(N__56685),
            .in2(_gnd_net_),
            .in3(N__54060),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83818),
            .ce(),
            .sr(N__54057));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_5_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_5_0  (
            .in0(N__54027),
            .in1(N__54005),
            .in2(N__54255),
            .in3(N__54279),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_5_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_14_5_1  (
            .in0(N__54291),
            .in1(N__78204),
            .in2(_gnd_net_),
            .in3(N__66123),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83822),
            .ce(N__65865),
            .sr(N__77262));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_14_5_2  (
            .in0(N__78201),
            .in1(N__54273),
            .in2(_gnd_net_),
            .in3(N__54261),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83822),
            .ce(N__65865),
            .sr(N__77262));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_5_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_14_5_3  (
            .in0(N__57366),
            .in1(N__78203),
            .in2(_gnd_net_),
            .in3(N__56835),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83822),
            .ce(N__65865),
            .sr(N__77262));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_5_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_14_5_4  (
            .in0(N__54246),
            .in1(N__54225),
            .in2(N__54219),
            .in3(N__54210),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_14_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_14_5_6  (
            .in0(N__78202),
            .in1(N__54492),
            .in2(_gnd_net_),
            .in3(N__74010),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83822),
            .ce(N__65865),
            .sr(N__77262));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_6_0  (
            .in0(N__63446),
            .in1(N__54188),
            .in2(_gnd_net_),
            .in3(N__54161),
            .lcout(\ppm_encoder_1.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_6_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_6_1  (
            .in0(N__74852),
            .in1(N__66609),
            .in2(N__59984),
            .in3(N__74701),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_6_2  (
            .in0(N__74700),
            .in1(N__66690),
            .in2(_gnd_net_),
            .in3(N__54537),
            .lcout(),
            .ltout(\ppm_encoder_1.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_6_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_6_3  (
            .in0(N__74853),
            .in1(_gnd_net_),
            .in2(N__54117),
            .in3(N__56802),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIVDMN_3_LC_14_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIVDMN_3_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIVDMN_3_LC_14_6_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIVDMN_3_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__66481),
            .in2(_gnd_net_),
            .in3(N__78266),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_14_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_14_6_5 .LUT_INIT=16'b1111001110100011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_14_6_5  (
            .in0(N__76694),
            .in1(N__56803),
            .in2(N__54315),
            .in3(N__74702),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_14_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_14_6_6 .LUT_INIT=16'b1100110111101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_14_6_6  (
            .in0(N__66523),
            .in1(N__77654),
            .in2(N__76220),
            .in3(N__76461),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83825),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI78NT_LC_14_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI78NT_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI78NT_LC_14_7_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI78NT_LC_14_7_0  (
            .in0(N__78229),
            .in1(N__66515),
            .in2(N__66438),
            .in3(N__56242),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_14_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_14_7_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54312),
            .in3(N__56712),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_14_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_14_7_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_14_7_2 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_14_7_2  (
            .in0(N__63618),
            .in1(N__74571),
            .in2(N__54309),
            .in3(N__76017),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83830),
            .ce(),
            .sr(N__77275));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_14_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_14_7_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_1_LC_14_7_3  (
            .in0(N__76693),
            .in1(N__76159),
            .in2(_gnd_net_),
            .in3(N__76457),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_7_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_14_7_4  (
            .in0(N__54306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56244),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83830),
            .ce(),
            .sr(N__77275));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_7_5 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_14_7_5  (
            .in0(N__56243),
            .in1(N__54305),
            .in2(N__56302),
            .in3(N__56713),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83830),
            .ce(),
            .sr(N__77275));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_7_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__56292),
            .in2(_gnd_net_),
            .in3(N__56241),
            .lcout(\ppm_encoder_1.PPM_STATE_53_d ),
            .ltout(\ppm_encoder_1.PPM_STATE_53_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_LC_14_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_LC_14_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_LC_14_7_7  (
            .in0(N__66514),
            .in1(N__66433),
            .in2(N__54366),
            .in3(N__78228),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_14_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_14_8_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_14_8_0  (
            .in0(N__59082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54350),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_6 ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_14_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_14_8_1 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_14_8_1  (
            .in0(N__66470),
            .in1(N__66552),
            .in2(N__54363),
            .in3(N__76097),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_14_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_14_8_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54360),
            .in3(N__76407),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_14_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_14_8_3 .LUT_INIT=16'b0101010110000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_14_8_3  (
            .in0(N__74788),
            .in1(N__63502),
            .in2(N__63060),
            .in3(N__66468),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_14_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_14_8_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_14_8_4  (
            .in0(N__66469),
            .in1(N__77657),
            .in2(N__54357),
            .in3(N__76409),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83836),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_8_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_8_5  (
            .in0(N__76408),
            .in1(N__63059),
            .in2(N__54354),
            .in3(N__77663),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83836),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_14_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_14_8_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_14_8_6  (
            .in0(N__66553),
            .in1(N__78259),
            .in2(N__66480),
            .in3(N__76406),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIGU6S2_4_LC_14_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIGU6S2_4_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIGU6S2_4_LC_14_8_7 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIGU6S2_4_LC_14_8_7  (
            .in0(N__59159),
            .in1(N__54341),
            .in2(N__54318),
            .in3(N__63218),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_9_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNIEL7O2_8_LC_14_9_0  (
            .in0(N__54478),
            .in1(N__63156),
            .in2(N__54438),
            .in3(N__63361),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIB72M6_8_LC_14_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIB72M6_8_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIB72M6_8_LC_14_9_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIB72M6_8_LC_14_9_1  (
            .in0(N__74070),
            .in1(_gnd_net_),
            .in2(N__54504),
            .in3(N__54501),
            .lcout(\ppm_encoder_1.throttle_RNIB72M6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIF43T2_8_LC_14_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIF43T2_8_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIF43T2_8_LC_14_9_2 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \ppm_encoder_1.throttle_RNIF43T2_8_LC_14_9_2  (
            .in0(N__59933),
            .in1(N__74026),
            .in2(N__54381),
            .in3(N__63257),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_14_9_3  (
            .in0(N__63500),
            .in1(N__54379),
            .in2(_gnd_net_),
            .in3(N__54436),
            .lcout(),
            .ltout(\ppm_encoder_1.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_9_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_14_9_4  (
            .in0(N__54479),
            .in1(_gnd_net_),
            .in2(N__54495),
            .in3(N__63034),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_8_LC_14_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_14_9_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_14_9_5  (
            .in0(N__60062),
            .in1(N__60042),
            .in2(N__62749),
            .in3(N__54480),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83844),
            .ce(),
            .sr(N__77288));
    defparam \ppm_encoder_1.elevator_8_LC_14_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_14_9_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_14_9_6  (
            .in0(N__54437),
            .in1(N__62739),
            .in2(N__54468),
            .in3(N__54456),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83844),
            .ce(),
            .sr(N__77288));
    defparam \ppm_encoder_1.throttle_8_LC_14_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_14_9_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_14_9_7  (
            .in0(N__54423),
            .in1(N__54411),
            .in2(N__62750),
            .in3(N__54380),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83844),
            .ce(),
            .sr(N__77288));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_10_0 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_14_10_0  (
            .in0(N__73986),
            .in1(N__74787),
            .in2(N__74894),
            .in3(N__56944),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_14_10_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_14_10_1  (
            .in0(N__78200),
            .in1(_gnd_net_),
            .in2(N__54636),
            .in3(N__54564),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83853),
            .ce(N__65874),
            .sr(N__77296));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_10_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_14_10_2  (
            .in0(N__54632),
            .in1(N__54609),
            .in2(N__54597),
            .in3(N__54588),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_10_3  (
            .in0(N__63501),
            .in1(N__54553),
            .in2(_gnd_net_),
            .in3(N__56924),
            .lcout(),
            .ltout(\ppm_encoder_1.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_10_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_10_4  (
            .in0(N__57203),
            .in1(_gnd_net_),
            .in2(N__54567),
            .in3(N__63055),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_10_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_14_10_5  (
            .in0(N__74786),
            .in1(N__74879),
            .in2(_gnd_net_),
            .in3(N__73934),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_10_6 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNIGN7O2_9_LC_14_10_6  (
            .in0(N__57202),
            .in1(N__63155),
            .in2(N__54557),
            .in3(N__63360),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI552R2_12_LC_14_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI552R2_12_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI552R2_12_LC_14_11_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNI552R2_12_LC_14_11_0  (
            .in0(N__54529),
            .in1(N__59952),
            .in2(N__54654),
            .in3(N__63267),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI2ABA6_12_LC_14_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI2ABA6_12_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI2ABA6_12_LC_14_11_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI2ABA6_12_LC_14_11_1  (
            .in0(N__66714),
            .in1(_gnd_net_),
            .in2(N__54513),
            .in3(N__54510),
            .lcout(\ppm_encoder_1.elevator_RNI2ABA6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_11_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_11_2  (
            .in0(N__54745),
            .in1(N__63165),
            .in2(N__54705),
            .in3(N__63372),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_11_3  (
            .in0(N__63503),
            .in1(N__54652),
            .in2(_gnd_net_),
            .in3(N__54703),
            .lcout(),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_11_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_11_4  (
            .in0(N__54746),
            .in1(_gnd_net_),
            .in2(N__54762),
            .in3(N__63047),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_14_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_14_11_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_14_11_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_14_11_5  (
            .in0(N__60852),
            .in1(N__60768),
            .in2(N__62737),
            .in3(N__54747),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83862),
            .ce(),
            .sr(N__77306));
    defparam \ppm_encoder_1.elevator_12_LC_14_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_14_11_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_14_11_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_14_11_6  (
            .in0(N__54704),
            .in1(N__62720),
            .in2(N__54735),
            .in3(N__54726),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83862),
            .ce(),
            .sr(N__77306));
    defparam \ppm_encoder_1.throttle_12_LC_14_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_14_11_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_14_11_7  (
            .in0(N__54690),
            .in1(N__54666),
            .in2(N__62738),
            .in3(N__54653),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83862),
            .ce(),
            .sr(N__77306));
    defparam \pid_side.state_RNIH98N9_1_LC_14_12_1 .C_ON=1'b0;
    defparam \pid_side.state_RNIH98N9_1_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIH98N9_1_LC_14_12_1 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \pid_side.state_RNIH98N9_1_LC_14_12_1  (
            .in0(N__57510),
            .in1(N__57516),
            .in2(N__67116),
            .in3(N__54999),
            .lcout(\pid_side.un1_reset_0_i ),
            .ltout(\pid_side.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIA3KT9_1_LC_14_12_2 .C_ON=1'b0;
    defparam \pid_side.state_RNIA3KT9_1_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIA3KT9_1_LC_14_12_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.state_RNIA3KT9_1_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54639),
            .in3(N__67094),
            .lcout(\pid_side.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_4_LC_14_12_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_4_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_4_LC_14_12_5 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \pid_side.source_pid_1_esr_4_LC_14_12_5  (
            .in0(N__63870),
            .in1(N__67730),
            .in2(N__67656),
            .in3(N__66838),
            .lcout(side_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83872),
            .ce(N__67444),
            .sr(N__67425));
    defparam \pid_side.source_pid_1_esr_5_LC_14_12_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_5_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_5_LC_14_12_6 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \pid_side.source_pid_1_esr_5_LC_14_12_6  (
            .in0(N__67729),
            .in1(N__60876),
            .in2(N__64236),
            .in3(N__67655),
            .lcout(side_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83872),
            .ce(N__67444),
            .sr(N__67425));
    defparam \pid_side.source_pid_1_esr_0_LC_14_12_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_0_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_0_LC_14_12_7 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \pid_side.source_pid_1_esr_0_LC_14_12_7  (
            .in0(N__67651),
            .in1(N__67731),
            .in2(N__66846),
            .in3(N__63936),
            .lcout(side_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83872),
            .ce(N__67444),
            .sr(N__67425));
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_13_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_13_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_13_0  (
            .in0(N__67623),
            .in1(N__64896),
            .in2(_gnd_net_),
            .in3(N__64413),
            .lcout(\pid_side.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_14_13_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_14_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNII463_20_LC_14_13_2  (
            .in0(N__64593),
            .in1(N__64629),
            .in2(N__64563),
            .in3(N__64260),
            .lcout(\pid_side.un11lto30_i_a2_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_10_LC_14_13_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_10_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_10_LC_14_13_3 .LUT_INIT=16'b1010101110101011;
    LogicCell40 \pid_side.source_pid_1_esr_10_LC_14_13_3  (
            .in0(N__64101),
            .in1(N__67625),
            .in2(N__67758),
            .in3(_gnd_net_),
            .lcout(side_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83883),
            .ce(N__67445),
            .sr(N__67428));
    defparam \pid_side.source_pid_1_esr_11_LC_14_13_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_11_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_11_LC_14_13_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_11_LC_14_13_4  (
            .in0(N__67624),
            .in1(N__67742),
            .in2(_gnd_net_),
            .in3(N__64056),
            .lcout(side_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83883),
            .ce(N__67445),
            .sr(N__67428));
    defparam \pid_side.source_pid_1_esr_6_LC_14_13_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_6_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_6_LC_14_13_5 .LUT_INIT=16'b1010101110101011;
    LogicCell40 \pid_side.source_pid_1_esr_6_LC_14_13_5  (
            .in0(N__64188),
            .in1(N__67626),
            .in2(N__67759),
            .in3(_gnd_net_),
            .lcout(side_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83883),
            .ce(N__67445),
            .sr(N__67428));
    defparam \pid_side.source_pid_1_esr_7_LC_14_13_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_7_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_7_LC_14_13_6 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \pid_side.source_pid_1_esr_7_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__67741),
            .in2(N__67649),
            .in3(N__64167),
            .lcout(side_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83883),
            .ce(N__67445),
            .sr(N__67428));
    defparam \pid_side.source_pid_1_esr_8_LC_14_13_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_8_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_8_LC_14_13_7 .LUT_INIT=16'b1010101110101011;
    LogicCell40 \pid_side.source_pid_1_esr_8_LC_14_13_7  (
            .in0(N__64134),
            .in1(N__67627),
            .in2(N__67760),
            .in3(_gnd_net_),
            .lcout(side_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83883),
            .ce(N__67445),
            .sr(N__67428));
    defparam \pid_side.error_i_acumm_12_LC_14_14_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_12_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_12_LC_14_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_side.error_i_acumm_12_LC_14_14_0  (
            .in0(N__67035),
            .in1(N__55343),
            .in2(_gnd_net_),
            .in3(N__55140),
            .lcout(\pid_side.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83894),
            .ce(N__55091),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_7_LC_14_14_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_7_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_7_LC_14_14_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_acumm_7_LC_14_14_1  (
            .in0(N__55141),
            .in1(N__67036),
            .in2(_gnd_net_),
            .in3(N__55374),
            .lcout(\pid_side.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83894),
            .ce(N__55091),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_8_LC_14_14_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_8_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_8_LC_14_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_side.error_i_acumm_8_LC_14_14_2  (
            .in0(N__67037),
            .in1(N__55254),
            .in2(_gnd_net_),
            .in3(N__55142),
            .lcout(\pid_side.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83894),
            .ce(N__55091),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_9_LC_14_14_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_9_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_9_LC_14_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_acumm_9_LC_14_14_3  (
            .in0(N__55143),
            .in1(N__67038),
            .in2(_gnd_net_),
            .in3(N__55398),
            .lcout(\pid_side.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83894),
            .ce(N__55091),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_0_LC_14_14_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_0_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_0_LC_14_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_i_acumm_0_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__55230),
            .in2(_gnd_net_),
            .in3(N__55139),
            .lcout(\pid_side.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83894),
            .ce(N__55091),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_14_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_14_14_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_14_14_7  (
            .in0(N__73877),
            .in1(N__76224),
            .in2(_gnd_net_),
            .in3(N__76608),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_3_LC_14_15_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_3_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_3_LC_14_15_0 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \pid_side.error_i_acumm_3_LC_14_15_0  (
            .in0(N__55127),
            .in1(N__54791),
            .in2(N__67140),
            .in3(N__55007),
            .lcout(\pid_side.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83902),
            .ce(N__55092),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_1_LC_14_15_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_1_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_1_LC_14_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_i_acumm_1_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__54807),
            .in2(_gnd_net_),
            .in3(N__55125),
            .lcout(\pid_side.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83902),
            .ce(N__55092),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_2_LC_14_15_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_2_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_2_LC_14_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_i_acumm_2_LC_14_15_2  (
            .in0(N__55126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54777),
            .lcout(\pid_side.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83902),
            .ce(N__55092),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_14_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_14_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_14_15_3  (
            .in0(N__54868),
            .in1(N__54847),
            .in2(N__54830),
            .in3(N__54768),
            .lcout(\pid_side.error_i_acumm16lt9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_14_15_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_14_15_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_14_15_4  (
            .in0(N__54806),
            .in1(N__55226),
            .in2(N__54795),
            .in3(N__54776),
            .lcout(\pid_side.un10lt9_1 ),
            .ltout(\pid_side.un10lt9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_14_15_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_14_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_14_15_5  (
            .in0(N__54869),
            .in1(N__54826),
            .in2(N__55020),
            .in3(N__54848),
            .lcout(),
            .ltout(\pid_side.un10lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_14_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_14_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_14_15_6  (
            .in0(N__55373),
            .in1(N__55394),
            .in2(N__55017),
            .in3(N__55253),
            .lcout(),
            .ltout(\pid_side.un10lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_14_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_14_15_7 .LUT_INIT=16'b0101010011111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_14_15_7  (
            .in0(N__55342),
            .in1(N__55284),
            .in2(N__55014),
            .in3(N__68358),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_14_16_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_14_16_0 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_14_16_0  (
            .in0(N__55041),
            .in1(N__55311),
            .in2(N__67169),
            .in3(N__55003),
            .lcout(\pid_side.error_i_acumm_2_sqmuxa_1 ),
            .ltout(\pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_14_16_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_14_16_1 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_14_16_1  (
            .in0(N__67117),
            .in1(N__67165),
            .in2(N__54882),
            .in3(N__54879),
            .lcout(\pid_side.error_i_acumm_2_sqmuxa ),
            .ltout(\pid_side.error_i_acumm_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_11_LC_14_16_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_11_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_11_LC_14_16_2 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \pid_side.error_i_acumm_11_LC_14_16_2  (
            .in0(N__55275),
            .in1(N__67121),
            .in2(N__54873),
            .in3(N__55160),
            .lcout(\pid_side.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_4_LC_14_16_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_4_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_4_LC_14_16_3 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \pid_side.error_i_acumm_4_LC_14_16_3  (
            .in0(N__55162),
            .in1(N__54870),
            .in2(N__67138),
            .in3(N__55122),
            .lcout(\pid_side.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_5_LC_14_16_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_5_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_5_LC_14_16_4 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \pid_side.error_i_acumm_5_LC_14_16_4  (
            .in0(N__55123),
            .in1(N__55163),
            .in2(N__54855),
            .in3(N__67128),
            .lcout(\pid_side.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_13_LC_14_16_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_13_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_13_LC_14_16_5 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \pid_side.error_i_acumm_13_LC_14_16_5  (
            .in0(N__55161),
            .in1(N__55212),
            .in2(N__67137),
            .in3(N__55121),
            .lcout(\pid_side.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_6_LC_14_16_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_6_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_6_LC_14_16_6 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \pid_side.error_i_acumm_6_LC_14_16_6  (
            .in0(N__55124),
            .in1(N__55164),
            .in2(N__54834),
            .in3(N__67129),
            .lcout(\pid_side.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_10_LC_14_16_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_10_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_10_LC_14_16_7 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \pid_side.error_i_acumm_10_LC_14_16_7  (
            .in0(N__55159),
            .in1(N__55302),
            .in2(N__67136),
            .in3(N__55120),
            .lcout(\pid_side.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83915),
            .ce(N__55084),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_14_17_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_14_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_14_17_0  (
            .in0(N__68235),
            .in1(N__68390),
            .in2(N__68414),
            .in3(N__68673),
            .lcout(\pid_side.error_i_acumm16lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_14_17_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_14_17_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_14_17_1  (
            .in0(N__55208),
            .in1(_gnd_net_),
            .in2(N__55032),
            .in3(N__58065),
            .lcout(\pid_side.error_i_acumm16lto27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_14_17_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_14_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_14_17_2  (
            .in0(N__55182),
            .in1(N__58055),
            .in2(N__55194),
            .in3(N__55173),
            .lcout(\pid_side.error_i_acumm16lto27_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_14_17_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_14_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_14_17_3  (
            .in0(N__68193),
            .in1(N__68250),
            .in2(N__68342),
            .in3(N__68292),
            .lcout(),
            .ltout(\pid_side.error_i_acumm16lto27_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_14_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_14_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_14_17_4  (
            .in0(N__55062),
            .in1(N__55056),
            .in2(N__55050),
            .in3(N__55047),
            .lcout(\pid_side.error_i_acumm16lto27_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_14_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_14_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_14_17_5  (
            .in0(N__55172),
            .in1(N__55190),
            .in2(N__58056),
            .in3(N__55181),
            .lcout(),
            .ltout(\pid_side.un10lto27_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_14_17_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_14_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_14_17_6  (
            .in0(N__58064),
            .in1(N__55207),
            .in2(N__55035),
            .in3(N__55028),
            .lcout(\pid_side.un10lto27_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_17_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_14_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_26_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64865),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83928),
            .ce(N__78354),
            .sr(N__77347));
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_14_18_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_14_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_0_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__58659),
            .in2(_gnd_net_),
            .in3(N__57540),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_18_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_13_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78978),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_14_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_21_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61101),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_14_18_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_14_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_23_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61182),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_14_18_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_22_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61056),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_18_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_9_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75544),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_14_18_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_14_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_24_LC_14_18_6  (
            .in0(N__61037),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_14_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_14_18_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_16_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__60893),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83941),
            .ce(N__78356),
            .sr(N__77352));
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_19_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_7_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75247),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83955),
            .ce(N__78358),
            .sr(N__77358));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_19_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__55267),
            .in2(_gnd_net_),
            .in3(N__55297),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_19_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_19_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_19_2  (
            .in0(N__55387),
            .in1(N__55241),
            .in2(_gnd_net_),
            .in3(N__55366),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_19_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_19_3 .LUT_INIT=16'b0100010001001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_19_3  (
            .in0(N__55353),
            .in1(N__55347),
            .in2(N__55323),
            .in3(N__55320),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_19_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_10_LC_14_19_4  (
            .in0(N__75409),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83955),
            .ce(N__78358),
            .sr(N__77358));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_19_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_19_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__55268),
            .in2(_gnd_net_),
            .in3(N__55298),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_19_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_19_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_11_LC_14_19_6  (
            .in0(N__68151),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83955),
            .ce(N__78358),
            .sr(N__77358));
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_19_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_8_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75157),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83955),
            .ce(N__78358),
            .sr(N__77358));
    defparam \pid_side.error_i_reg_esr_13_LC_14_20_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_13_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_13_LC_14_20_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_13_LC_14_20_0  (
            .in0(N__62103),
            .in1(N__65280),
            .in2(_gnd_net_),
            .in3(N__61308),
            .lcout(\pid_side.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83968),
            .ce(N__69305),
            .sr(N__77364));
    defparam \pid_side.error_i_reg_esr_26_LC_14_20_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_26_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_26_LC_14_20_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_26_LC_14_20_1  (
            .in0(N__59244),
            .in1(N__61478),
            .in2(_gnd_net_),
            .in3(N__55626),
            .lcout(\pid_side.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83968),
            .ce(N__69305),
            .sr(N__77364));
    defparam \pid_side.error_i_reg_esr_7_LC_14_20_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_7_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_7_LC_14_20_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_side.error_i_reg_esr_7_LC_14_20_2  (
            .in0(N__65448),
            .in1(N__58698),
            .in2(_gnd_net_),
            .in3(N__55482),
            .lcout(\pid_side.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83968),
            .ce(N__69305),
            .sr(N__77364));
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_14_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_14_20_3 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_14_20_3  (
            .in0(N__73830),
            .in1(_gnd_net_),
            .in2(N__76609),
            .in3(N__76271),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_5  (
            .in0(N__76534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.N_2569_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_14_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_14_20_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__74176),
            .in3(N__76530),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_14_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_14_20_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_14_20_7  (
            .in0(N__76529),
            .in1(N__74164),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m64_e_LC_14_21_1 .C_ON=1'b0;
    defparam \pid_front.m64_e_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.m64_e_LC_14_21_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.m64_e_LC_14_21_1  (
            .in0(N__57657),
            .in1(N__57626),
            .in2(_gnd_net_),
            .in3(N__57684),
            .lcout(pid_front_N_331),
            .ltout(pid_front_N_331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m70_0_LC_14_21_2 .C_ON=1'b0;
    defparam \pid_front.m70_0_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.m70_0_LC_14_21_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_front.m70_0_LC_14_21_2  (
            .in0(N__69536),
            .in1(_gnd_net_),
            .in2(N__55446),
            .in3(N__70500),
            .lcout(pid_side_N_166_mux),
            .ltout(pid_side_N_166_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_3_LC_14_21_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_3_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_3_LC_14_21_3 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \pid_front.error_i_reg_esr_3_LC_14_21_3  (
            .in0(N__70706),
            .in1(N__55518),
            .in2(N__55443),
            .in3(N__55440),
            .lcout(\pid_front.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83984),
            .ce(N__59347),
            .sr(N__77368));
    defparam \pid_front.error_i_reg_9_sn_19_LC_14_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_9_sn_19_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_9_sn_19_LC_14_21_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \pid_front.error_i_reg_9_sn_19_LC_14_21_4  (
            .in0(N__69535),
            .in1(N__70499),
            .in2(_gnd_net_),
            .in3(N__69765),
            .lcout(pid_front_error_i_reg_9_sn_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIP9BO5_LC_14_21_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIP9BO5_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIP9BO5_LC_14_21_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_side.error_cry_2_c_RNIP9BO5_LC_14_21_5  (
            .in0(N__66045),
            .in1(N__58755),
            .in2(_gnd_net_),
            .in3(N__62024),
            .lcout(\pid_side.N_41_0 ),
            .ltout(\pid_side.N_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_14_21_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_14_21_6 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_26_LC_14_21_6  (
            .in0(N__69537),
            .in1(N__69766),
            .in2(N__55629),
            .in3(N__70079),
            .lcout(\pid_side.error_i_reg_9_rn_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI75LOB_LC_14_22_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI75LOB_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI75LOB_LC_14_22_0 .LUT_INIT=16'b0010000000101111;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI75LOB_LC_14_22_0  (
            .in0(N__61744),
            .in1(N__65742),
            .in2(N__70495),
            .in3(N__55857),
            .lcout(\pid_front.m8_2_03_3_i_0 ),
            .ltout(\pid_front.m8_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_4_LC_14_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_4_LC_14_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_4_LC_14_22_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \pid_front.error_i_reg_4_LC_14_22_1  (
            .in0(N__55616),
            .in1(N__65407),
            .in2(N__55620),
            .in3(N__55592),
            .lcout(\pid_front.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84002),
            .ce(),
            .sr(N__77375));
    defparam \pid_front.error_i_reg_11_LC_14_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_11_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_11_LC_14_22_2 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \pid_front.error_i_reg_11_LC_14_22_2  (
            .in0(N__65406),
            .in1(N__55532),
            .in2(N__55593),
            .in3(N__55554),
            .lcout(\pid_front.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84002),
            .ce(),
            .sr(N__77375));
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_14_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_14_22_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_15_LC_14_22_3  (
            .in0(N__65741),
            .in1(N__70408),
            .in2(_gnd_net_),
            .in3(N__55514),
            .lcout(\pid_front.m3_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_22_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_22_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_7_LC_14_22_4  (
            .in0(N__70407),
            .in1(N__65740),
            .in2(_gnd_net_),
            .in3(N__58678),
            .lcout(\pid_side.error_i_reg_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNI9UJ94_LC_14_22_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNI9UJ94_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNI9UJ94_LC_14_22_5 .LUT_INIT=16'b1010001010100111;
    LogicCell40 \pid_side.error_cry_6_c_RNI9UJ94_LC_14_22_5  (
            .in0(N__65508),
            .in1(N__71236),
            .in2(N__72276),
            .in3(N__71326),
            .lcout(\pid_side.N_49_0 ),
            .ltout(\pid_side.N_49_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_14_22_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_15_LC_14_22_6 .LUT_INIT=16'b0001001110011011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_15_LC_14_22_6  (
            .in0(N__70403),
            .in1(N__65739),
            .in2(N__55473),
            .in3(N__58865),
            .lcout(),
            .ltout(\pid_side.m134_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_22_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_22_7 .LUT_INIT=16'b0001111100011010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_15_LC_14_22_7  (
            .in0(N__70409),
            .in1(N__70083),
            .in2(N__55470),
            .in3(N__58200),
            .lcout(\pid_side.m19_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI9I2A2_LC_14_23_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI9I2A2_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI9I2A2_LC_14_23_0 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_side.error_cry_0_c_RNI9I2A2_LC_14_23_0  (
            .in0(N__73590),
            .in1(N__55661),
            .in2(N__65697),
            .in3(N__55649),
            .lcout(\pid_side.error_cry_0_c_RNI9I2AZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNIUIKS_LC_14_23_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNIUIKS_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNIUIKS_LC_14_23_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_side.error_cry_1_c_RNIUIKS_LC_14_23_1  (
            .in0(N__72677),
            .in1(N__73068),
            .in2(_gnd_net_),
            .in3(N__73160),
            .lcout(\pid_side.N_11_0 ),
            .ltout(\pid_side.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI3DQV1_LC_14_23_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI3DQV1_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI3DQV1_LC_14_23_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_0_c_RNI3DQV1_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__72253),
            .in2(N__55665),
            .in3(N__55660),
            .lcout(\pid_side.N_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI1D101_LC_14_23_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI1D101_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI1D101_LC_14_23_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_0_c_RNI1D101_LC_14_23_3  (
            .in0(N__71559),
            .in1(N__69156),
            .in2(_gnd_net_),
            .in3(N__71670),
            .lcout(\pid_side.N_14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_23_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_23_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_15_LC_14_23_4  (
            .in0(N__73591),
            .in1(N__55662),
            .in2(N__65698),
            .in3(N__55650),
            .lcout(),
            .ltout(\pid_side.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_14_23_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_14_23_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_15_LC_14_23_5  (
            .in0(N__70528),
            .in1(_gnd_net_),
            .in2(N__55641),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_15_LC_14_23_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_15_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_15_LC_14_23_6 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_side.error_i_reg_esr_15_LC_14_23_6  (
            .in0(N__69634),
            .in1(N__69865),
            .in2(N__55638),
            .in3(N__55635),
            .lcout(\pid_side.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84020),
            .ce(N__69323),
            .sr(N__77381));
    defparam \pid_side.error_cry_0_c_RNIUPMV_LC_14_23_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIUPMV_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIUPMV_LC_14_23_7 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_0_c_RNIUPMV_LC_14_23_7  (
            .in0(N__72678),
            .in1(N__71671),
            .in2(N__72271),
            .in3(N__73159),
            .lcout(\pid_side.g0_i_m4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_14_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_14_24_0 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_20_LC_14_24_0  (
            .in0(N__55887),
            .in1(N__70471),
            .in2(N__55908),
            .in3(N__55914),
            .lcout(),
            .ltout(\pid_front.m24_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_20_LC_14_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_20_LC_14_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_20_LC_14_24_1 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_front.error_i_reg_esr_20_LC_14_24_1  (
            .in0(N__69633),
            .in1(N__69847),
            .in2(N__55950),
            .in3(N__55947),
            .lcout(\pid_front.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84034),
            .ce(N__59425),
            .sr(N__77386));
    defparam \pid_front.error_cry_10_c_RNI6VKA3_LC_14_24_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNI6VKA3_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNI6VKA3_LC_14_24_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \pid_front.error_cry_10_c_RNI6VKA3_LC_14_24_2  (
            .in0(N__72971),
            .in1(N__56495),
            .in2(_gnd_net_),
            .in3(N__56029),
            .lcout(\pid_front.N_57_0 ),
            .ltout(\pid_front.N_57_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_14_24_3 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_24_LC_14_24_3  (
            .in0(N__56497),
            .in1(N__70656),
            .in2(N__55923),
            .in3(N__70468),
            .lcout(\pid_front.error_i_reg_esr_RNO_0_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_14_24_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_14_24_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_20_LC_14_24_4  (
            .in0(N__70467),
            .in1(N__65985),
            .in2(_gnd_net_),
            .in3(N__56496),
            .lcout(\pid_front.m138_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_14_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_14_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_12_LC_14_24_5  (
            .in0(N__65696),
            .in1(N__55903),
            .in2(_gnd_net_),
            .in3(N__55886),
            .lcout(),
            .ltout(\pid_front.N_129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .LUT_INIT=16'b0100110010001000;
    LogicCell40 \pid_front.error_i_reg_esr_12_LC_14_24_6  (
            .in0(N__61710),
            .in1(N__69866),
            .in2(N__55878),
            .in3(N__55839),
            .lcout(\pid_front.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84034),
            .ce(N__59425),
            .sr(N__77386));
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_14_24_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_14_24_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_12_LC_14_24_7  (
            .in0(N__69632),
            .in1(N__61709),
            .in2(_gnd_net_),
            .in3(N__55853),
            .lcout(\pid_front.error_i_reg_9_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIU0FF1_LC_14_25_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNIU0FF1_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIU0FF1_LC_14_25_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_7_c_RNIU0FF1_LC_14_25_0  (
            .in0(N__71450),
            .in1(N__55818),
            .in2(_gnd_net_),
            .in3(N__55740),
            .lcout(\pid_front.N_18_1 ),
            .ltout(\pid_front.N_18_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNI14OF3_LC_14_25_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_7_c_RNI14OF3_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNI14OF3_LC_14_25_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_7_c_RNI14OF3_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__73592),
            .in2(N__55668),
            .in3(N__56028),
            .lcout(\pid_front.N_37_1 ),
            .ltout(\pid_front.N_37_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_25_2 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_22_LC_14_25_2  (
            .in0(N__56519),
            .in1(N__70639),
            .in2(N__56166),
            .in3(N__70251),
            .lcout(\pid_front.m26_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIU65R1_LC_14_25_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_8_c_RNIU65R1_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIU65R1_LC_14_25_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_8_c_RNIU65R1_LC_14_25_3  (
            .in0(N__72663),
            .in1(N__56156),
            .in2(_gnd_net_),
            .in3(N__56082),
            .lcout(\pid_front.N_36_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_25_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_25_4 .LUT_INIT=16'b0000001111111010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_14_LC_14_25_4  (
            .in0(N__70773),
            .in1(N__70099),
            .in2(N__70514),
            .in3(N__58782),
            .lcout(),
            .ltout(\pid_side.m18_2_03_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_14_LC_14_25_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_14_LC_14_25_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_14_LC_14_25_5 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_14_LC_14_25_5  (
            .in0(N__69635),
            .in1(N__69953),
            .in2(N__56007),
            .in3(N__56004),
            .lcout(\pid_side.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84050),
            .ce(N__69316),
            .sr(N__77391));
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_25_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_25_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_14_LC_14_25_6  (
            .in0(N__70638),
            .in1(N__70250),
            .in2(_gnd_net_),
            .in3(N__58773),
            .lcout(\pid_side.m2_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNI6G8L2_LC_14_26_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI6G8L2_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI6G8L2_LC_14_26_0 .LUT_INIT=16'b0010000001110101;
    LogicCell40 \pid_front.error_cry_0_c_RNI6G8L2_LC_14_26_0  (
            .in0(N__72959),
            .in1(N__71578),
            .in2(N__61833),
            .in3(N__55998),
            .lcout(\pid_front.m2_0_03_3_i_0 ),
            .ltout(\pid_front.m2_0_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_1  (
            .in0(N__61634),
            .in1(_gnd_net_),
            .in2(N__55974),
            .in3(N__70457),
            .lcout(),
            .ltout(\pid_front.m2_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2  (
            .in0(N__69949),
            .in1(N__69565),
            .in2(N__55971),
            .in3(N__59021),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_14_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__62151),
            .in2(N__55968),
            .in3(N__56388),
            .lcout(\pid_front.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84067),
            .ce(N__59426),
            .sr(N__77394));
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_26_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_26_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_14_LC_14_26_4  (
            .in0(N__70702),
            .in1(N__56541),
            .in2(_gnd_net_),
            .in3(N__56520),
            .lcout(\pid_front.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNI15TSB_LC_14_26_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_0_c_RNI15TSB_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNI15TSB_LC_14_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_2_0_c_RNI15TSB_LC_14_26_5  (
            .in0(N__56378),
            .in1(N__56358),
            .in2(_gnd_net_),
            .in3(N__56352),
            .lcout(\pid_front.N_110 ),
            .ltout(\pid_front.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_6 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_6  (
            .in0(N__70458),
            .in1(N__61635),
            .in2(N__56346),
            .in3(N__59199),
            .lcout(),
            .ltout(\pid_front.m10_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_7 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_front.error_i_reg_esr_22_LC_14_26_7  (
            .in0(N__69566),
            .in1(N__69950),
            .in2(N__56343),
            .in3(N__56340),
            .lcout(\pid_front.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84067),
            .ce(N__59426),
            .sr(N__77394));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_14_27_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_14_27_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_14_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80493),
            .lcout(xy_ki_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84081),
            .ce(N__73413),
            .sr(N__77399));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_3_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_3_0  (
            .in0(N__56185),
            .in1(N__56623),
            .in2(N__56315),
            .in3(N__56203),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_3_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_3_1  (
            .in0(N__56624),
            .in1(N__56186),
            .in2(N__56208),
            .in3(N__56263),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_2  (
            .in0(N__56658),
            .in1(N__56202),
            .in2(N__56652),
            .in3(N__56184),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_15_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_15_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_15_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_15_3_3  (
            .in0(N__78198),
            .in1(N__62898),
            .in2(_gnd_net_),
            .in3(N__56817),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83819),
            .ce(N__65855),
            .sr(N__77255));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_15_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_15_3_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_15_3_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_15_3_4  (
            .in0(N__59577),
            .in1(N__78199),
            .in2(_gnd_net_),
            .in3(N__56829),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83819),
            .ce(N__65855),
            .sr(N__77255));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_3_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_15_3_5  (
            .in0(N__78196),
            .in1(N__56769),
            .in2(_gnd_net_),
            .in3(N__56643),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83819),
            .ce(N__65855),
            .sr(N__77255));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_3_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_3_6  (
            .in0(N__56631),
            .in1(N__56622),
            .in2(N__56577),
            .in3(N__56605),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_15_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_15_3_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_15_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_15_3_7  (
            .in0(N__78197),
            .in1(N__57078),
            .in2(_gnd_net_),
            .in3(N__56589),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83819),
            .ce(N__65855),
            .sr(N__77255));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_15_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__56568),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_15_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__56562),
            .in2(N__60598),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_4_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_15_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__56556),
            .in2(N__60593),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_4_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_15_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__56547),
            .in2(N__60595),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_4_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_15_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__56760),
            .in2(N__60594),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_4_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_15_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__56745),
            .in2(N__60596),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_4_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_15_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__60560),
            .in2(N__56733),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_4_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_15_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(N__66288),
            .in2(N__60597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_5_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_15_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__62346),
            .in2(N__60547),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_5_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_15_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(N__60494),
            .in2(N__56667),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56724),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(N__62307),
            .in2(_gnd_net_),
            .in3(N__56683),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(N__77616),
            .in2(_gnd_net_),
            .in3(N__76527),
            .lcout(\ppm_encoder_1.N_2569_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_5_5 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_5_5  (
            .in0(N__57060),
            .in1(N__74857),
            .in2(N__74743),
            .in3(N__74229),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_15_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_15_5_7 .LUT_INIT=16'b1101110111010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_15_5_7  (
            .in0(N__56807),
            .in1(N__74858),
            .in2(N__74744),
            .in3(N__76674),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_6_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_6_0  (
            .in0(N__74714),
            .in1(N__63433),
            .in2(N__62996),
            .in3(N__76147),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_6_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_6_1  (
            .in0(N__74732),
            .in1(N__77655),
            .in2(N__56820),
            .in3(N__76462),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83831),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_15_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_15_6_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_15_6_2  (
            .in0(N__56798),
            .in1(N__74854),
            .in2(N__74742),
            .in3(N__74109),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_6_3 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_6_3  (
            .in0(N__56882),
            .in1(N__56865),
            .in2(N__76528),
            .in3(N__77656),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83831),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_6_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_15_6_5  (
            .in0(N__63432),
            .in1(N__66482),
            .in2(_gnd_net_),
            .in3(N__66519),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_15_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_15_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_15_6_6  (
            .in0(N__63445),
            .in1(N__59492),
            .in2(_gnd_net_),
            .in3(N__59508),
            .lcout(),
            .ltout(\ppm_encoder_1.N_286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_15_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_15_6_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_15_6_7  (
            .in0(N__59469),
            .in1(_gnd_net_),
            .in2(N__56772),
            .in3(N__62956),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_7_0 .LUT_INIT=16'b1010101111101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_7_0  (
            .in0(N__77649),
            .in1(N__59084),
            .in2(N__76219),
            .in3(N__76401),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83837),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_7_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_15_7_1  (
            .in0(N__76400),
            .in1(N__56883),
            .in2(N__66563),
            .in3(N__77653),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83837),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_7_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_15_7_2  (
            .in0(N__56850),
            .in1(N__56871),
            .in2(N__77667),
            .in3(N__76402),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83837),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__56848),
            .in2(_gnd_net_),
            .in3(N__56864),
            .lcout(\ppm_encoder_1.N_221 ),
            .ltout(\ppm_encoder_1.N_221_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIMSNT_0_LC_15_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIMSNT_0_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIMSNT_0_LC_15_7_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIMSNT_0_LC_15_7_4  (
            .in0(N__66419),
            .in1(N__59083),
            .in2(N__56853),
            .in3(N__76399),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_15_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_15_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__66551),
            .in2(_gnd_net_),
            .in3(N__56849),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_0_LC_15_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_0_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_0_LC_15_7_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI7RM01_0_LC_15_7_6  (
            .in0(N__66418),
            .in1(N__78227),
            .in2(N__66524),
            .in3(N__76398),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_15_7_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI077O2_1_LC_15_7_7  (
            .in0(N__57155),
            .in1(N__57107),
            .in2(N__56838),
            .in3(N__63326),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_8_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNI6D7O2_4_LC_15_8_0  (
            .in0(N__57237),
            .in1(N__63117),
            .in2(N__59129),
            .in3(N__63329),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI0L5L6_4_LC_15_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI0L5L6_4_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI0L5L6_4_LC_15_8_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI0L5L6_4_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__66950),
            .in2(N__57024),
            .in3(N__57021),
            .lcout(\ppm_encoder_1.elevator_RNI0L5L6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNII07S2_5_LC_15_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNII07S2_5_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNII07S2_5_LC_15_8_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNII07S2_5_LC_15_8_2  (
            .in0(N__59936),
            .in1(N__66212),
            .in2(N__57006),
            .in3(N__63223),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI5Q5L6_5_LC_15_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5Q5L6_5_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5Q5L6_5_LC_15_8_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI5Q5L6_5_LC_15_8_3  (
            .in0(N__66251),
            .in1(_gnd_net_),
            .in2(N__57015),
            .in3(N__57012),
            .lcout(\ppm_encoder_1.elevator_RNI5Q5L6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_8_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI8F7O2_5_LC_15_8_4  (
            .in0(N__56962),
            .in1(N__63116),
            .in2(N__57390),
            .in3(N__63328),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_8_5  (
            .in0(N__63498),
            .in1(N__57005),
            .in2(_gnd_net_),
            .in3(N__57389),
            .lcout(),
            .ltout(\ppm_encoder_1.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_8_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_8_6  (
            .in0(N__56963),
            .in1(_gnd_net_),
            .in2(N__56979),
            .in3(N__62999),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_5_LC_15_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_5_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_5_LC_15_8_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_5_LC_15_8_7  (
            .in0(N__60183),
            .in1(N__60159),
            .in2(N__62751),
            .in3(N__56964),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83845),
            .ce(),
            .sr(N__77289));
    defparam \ppm_encoder_1.throttle_RNIH63T2_9_LC_15_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIH63T2_9_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIH63T2_9_LC_15_9_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIH63T2_9_LC_15_9_0  (
            .in0(N__56952),
            .in1(N__59946),
            .in2(N__56925),
            .in3(N__63258),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGC2M6_9_LC_15_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGC2M6_9_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGC2M6_9_LC_15_9_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIGC2M6_9_LC_15_9_1  (
            .in0(N__73958),
            .in1(_gnd_net_),
            .in2(N__56892),
            .in3(N__56889),
            .lcout(\ppm_encoder_1.throttle_RNIGC2M6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNIRV873_14_LC_15_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNIRV873_14_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNIRV873_14_LC_15_9_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNIRV873_14_LC_15_9_2  (
            .in0(N__74645),
            .in1(N__59947),
            .in2(N__57129),
            .in3(N__63259),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIG1J17_14_LC_15_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIG1J17_14_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIG1J17_14_LC_15_9_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIG1J17_14_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__74934),
            .in2(N__57132),
            .in3(N__59583),
            .lcout(\ppm_encoder_1.aileron_esr_RNIG1J17Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_15_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_15_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_15_9_4  (
            .in0(N__57128),
            .in1(N__63489),
            .in2(_gnd_net_),
            .in3(N__59603),
            .lcout(),
            .ltout(\ppm_encoder_1.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_15_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_15_9_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__63035),
            .in2(N__57111),
            .in3(N__60744),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_9_6  (
            .in0(N__63036),
            .in1(N__57066),
            .in2(_gnd_net_),
            .in3(N__57108),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_9_7  (
            .in0(N__63488),
            .in1(N__59064),
            .in2(_gnd_net_),
            .in3(N__57156),
            .lcout(\ppm_encoder_1.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI772R2_13_LC_15_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI772R2_13_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI772R2_13_LC_15_10_0 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \ppm_encoder_1.throttle_RNI772R2_13_LC_15_10_0  (
            .in0(N__59956),
            .in1(N__57059),
            .in2(N__57252),
            .in3(N__63263),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI7FBA6_13_LC_15_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI7FBA6_13_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI7FBA6_13_LC_15_10_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI7FBA6_13_LC_15_10_1  (
            .in0(N__66660),
            .in1(_gnd_net_),
            .in2(N__57033),
            .in3(N__57030),
            .lcout(\ppm_encoder_1.elevator_RNI7FBA6Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_15_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_15_10_2 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNI68LH2_13_LC_15_10_2  (
            .in0(N__57349),
            .in1(N__63160),
            .in2(N__57306),
            .in3(N__63363),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_10_3  (
            .in0(N__63491),
            .in1(N__57250),
            .in2(_gnd_net_),
            .in3(N__57304),
            .lcout(),
            .ltout(\ppm_encoder_1.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_10_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_10_4  (
            .in0(N__57350),
            .in1(_gnd_net_),
            .in2(N__57369),
            .in3(N__63037),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_15_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_15_10_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_15_10_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_15_10_5  (
            .in0(N__60756),
            .in1(N__57351),
            .in2(N__67485),
            .in3(N__62632),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83863),
            .ce(),
            .sr(N__77307));
    defparam \ppm_encoder_1.elevator_13_LC_15_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_15_10_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_15_10_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_15_10_6  (
            .in0(N__57305),
            .in1(N__57339),
            .in2(N__62694),
            .in3(N__57318),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83863),
            .ce(),
            .sr(N__77307));
    defparam \ppm_encoder_1.throttle_13_LC_15_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_15_10_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_15_10_7 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_15_10_7  (
            .in0(N__57291),
            .in1(N__57251),
            .in2(N__57267),
            .in3(N__62633),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83863),
            .ce(),
            .sr(N__77307));
    defparam \ppm_encoder_1.aileron_4_LC_15_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_4_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_4_LC_15_11_0 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_4_LC_15_11_0  (
            .in0(N__57236),
            .in1(N__60192),
            .in2(N__62707),
            .in3(N__60206),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_11_1  (
            .in0(N__63054),
            .in1(N__59097),
            .in2(_gnd_net_),
            .in3(N__57235),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_9_LC_15_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_15_11_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_15_11_2  (
            .in0(N__60027),
            .in1(N__67674),
            .in2(N__62708),
            .in3(N__57204),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \ppm_encoder_1.elevator_1_LC_15_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_1_LC_15_11_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_1_LC_15_11_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ppm_encoder_1.elevator_1_LC_15_11_3  (
            .in0(N__57154),
            .in1(N__62639),
            .in2(N__57189),
            .in3(N__57165),
            .lcout(\ppm_encoder_1.elevatorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \ppm_encoder_1.elevator_10_LC_15_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_15_11_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_15_11_4  (
            .in0(N__57486),
            .in1(N__57465),
            .in2(N__62709),
            .in3(N__59837),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \ppm_encoder_1.elevator_4_LC_15_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_4_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_4_LC_15_11_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_4_LC_15_11_5  (
            .in0(N__57453),
            .in1(N__57444),
            .in2(N__59128),
            .in3(N__62652),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \ppm_encoder_1.elevator_5_LC_15_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_5_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_5_LC_15_11_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_5_LC_15_11_6  (
            .in0(N__57423),
            .in1(N__57414),
            .in2(N__62710),
            .in3(N__57385),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83873),
            .ce(),
            .sr(N__77315));
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_12_0 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__60243),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\pid_side.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_12_1 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__60228),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2 ),
            .carryout(\pid_side.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_12_2 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__60858),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_0 ),
            .carryout(\pid_side.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_12_3 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__63780),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_1 ),
            .carryout(\pid_side.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_12_4 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_4_c_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__63771),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_2 ),
            .carryout(\pid_side.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_12_5 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_5_c_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__57556),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_3 ),
            .carryout(\pid_side.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_12_6 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_6_c_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__57594),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_4 ),
            .carryout(\pid_side.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_12_7 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__57577),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_5 ),
            .carryout(\pid_side.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_13_0 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_13_0 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_13_0  (
            .in0(N__67526),
            .in1(N__67632),
            .in2(N__64023),
            .in3(N__57525),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_o2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_15_13_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_15_13_1 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_15_13_1  (
            .in0(N__67546),
            .in1(N__66831),
            .in2(N__67650),
            .in3(N__57522),
            .lcout(\pid_side.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_13_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_13_2  (
            .in0(N__60872),
            .in1(N__60237),
            .in2(N__60252),
            .in3(N__67545),
            .lcout(\pid_side.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_15_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_15_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__57504),
            .in2(_gnd_net_),
            .in3(N__77618),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_15_13_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_15_13_4 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIRALN2_4_LC_15_13_4  (
            .in0(N__60871),
            .in1(N__67631),
            .in2(N__64235),
            .in3(N__63866),
            .lcout(\pid_side.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIVRQ8_20_LC_15_13_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIVRQ8_20_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIVRQ8_20_LC_15_13_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIVRQ8_20_LC_15_13_6  (
            .in0(N__57558),
            .in1(N__57579),
            .in2(_gnd_net_),
            .in3(N__57593),
            .lcout(),
            .ltout(\pid_side.pid_prereg_esr_RNIVRQ8Z0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_15_13_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_15_13_7 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIIATS_12_LC_15_13_7  (
            .in0(N__64022),
            .in1(N__63960),
            .in2(N__57489),
            .in3(N__67527),
            .lcout(\pid_side.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_15_14_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_15_14_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIV4S38_10_LC_15_14_0  (
            .in0(N__75432),
            .in1(N__75900),
            .in2(N__68175),
            .in3(N__75410),
            .lcout(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m101_e_LC_15_14_1 .C_ON=1'b0;
    defparam \pid_side.m101_e_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m101_e_LC_15_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.m101_e_LC_15_14_1  (
            .in0(N__57610),
            .in1(N__57643),
            .in2(N__69534),
            .in3(N__57673),
            .lcout(pid_side_N_166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_15_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_15_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_5_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80089),
            .lcout(xy_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83903),
            .ce(N__73383),
            .sr(N__77336));
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_15_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_15_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_15_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_6_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81093),
            .lcout(xy_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83903),
            .ce(N__73383),
            .sr(N__77336));
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_15_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_7_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79908),
            .lcout(xy_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83903),
            .ce(N__73383),
            .sr(N__77336));
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_15_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_15_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_4_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79284),
            .lcout(xy_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83903),
            .ce(N__73383),
            .sr(N__77336));
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_14_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_14_6  (
            .in0(N__64476),
            .in1(N__64500),
            .in2(N__64452),
            .in3(N__64530),
            .lcout(\pid_side.un11lto30_i_a2_5_and ),
            .ltout(\pid_side.un11lto30_i_a2_5_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_14_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_14_7  (
            .in0(N__57578),
            .in1(N__63959),
            .in2(N__57561),
            .in3(N__57557),
            .lcout(\pid_side.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_15_15_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_15_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIARAI_0_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__57536),
            .in2(N__58658),
            .in3(_gnd_net_),
            .lcout(\pid_side.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_15_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__57789),
            .in2(N__58635),
            .in3(N__57783),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_15_2 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__57780),
            .in2(N__58623),
            .in3(N__57774),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_15_15_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_15_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__57771),
            .in2(N__58845),
            .in3(N__57765),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_15_4 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__57762),
            .in2(N__61446),
            .in3(N__57756),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_15_5 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__57753),
            .in2(N__61503),
            .in3(N__57744),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_15_6 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__61410),
            .in2(N__57741),
            .in3(N__57732),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_15_15_7 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_15_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__57729),
            .in2(N__57717),
            .in3(N__57708),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_16_0 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIIDSN_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__57705),
            .in2(N__62205),
            .in3(N__57696),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNIIDSN ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_16_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNICNNJ_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__57693),
            .in2(N__65325),
            .in3(N__57888),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNICNNJ ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_16_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI6OOI_10_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__57885),
            .in2(N__61461),
            .in3(N__57879),
            .lcout(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_16_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIGRJR_11_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__57876),
            .in2(N__58179),
            .in3(N__57870),
            .lcout(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_16_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIJVKR_12_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__57867),
            .in2(N__62067),
            .in3(N__57855),
            .lcout(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_16_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM3MR_13_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__58102),
            .in2(N__57852),
            .in3(N__57837),
            .lcout(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_16_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO6NR_14_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__57834),
            .in2(N__58134),
            .in3(N__57819),
            .lcout(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_16_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__58106),
            .in2(N__57816),
            .in3(N__57798),
            .lcout(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_17_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISCPR_16_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__58107),
            .in2(N__61854),
            .in3(N__57795),
            .lcout(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_17_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUFQR_17_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__58830),
            .in2(N__58135),
            .in3(N__57792),
            .lcout(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_17_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI0JRR_18_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__58111),
            .in2(N__58593),
            .in3(N__57924),
            .lcout(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_17_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI2MSR_19_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__58602),
            .in2(N__58136),
            .in3(N__57921),
            .lcout(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_17_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIRGUR_20_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__58115),
            .in2(N__65535),
            .in3(N__57918),
            .lcout(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_17_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIK2OS_21_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__65571),
            .in2(N__58137),
            .in3(N__57915),
            .lcout(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_17_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM5PS_22_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__58119),
            .in2(N__69342),
            .in3(N__57912),
            .lcout(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_17_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO8QS_23_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__58806),
            .in2(N__58138),
            .in3(N__57909),
            .lcout(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_18_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQBRS_24_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__58794),
            .in2(N__58148),
            .in3(N__57906),
            .lcout(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_18_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISESS_25_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__58142),
            .in2(N__61527),
            .in3(N__57903),
            .lcout(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_18_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUHTS_26_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__57900),
            .in2(N__58149),
            .in3(N__57891),
            .lcout(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_18_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__58146),
            .in2(N__58167),
            .in3(N__58152),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_18_4 .C_ON=1'b0;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_15_18_4  (
            .in0(N__58147),
            .in1(N__58166),
            .in2(_gnd_net_),
            .in3(N__58068),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_18_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_15_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_28_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61380),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83956),
            .ce(N__78359),
            .sr(N__77359));
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_18_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_15_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_27_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61230),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83956),
            .ce(N__78359),
            .sr(N__77359));
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_15_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_15_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_25_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64832),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83956),
            .ce(N__78359),
            .sr(N__77359));
    defparam \dron_frame_decoder_1.source_H_disp_side_14_LC_15_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_14_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_14_LC_15_19_0 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_14_LC_15_19_0  (
            .in0(N__68563),
            .in1(N__71724),
            .in2(N__71970),
            .in3(N__68860),
            .lcout(drone_H_disp_side_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83969),
            .ce(),
            .sr(N__77365));
    defparam \dron_frame_decoder_1.state_RNI44RU_5_LC_15_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI44RU_5_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI44RU_5_LC_15_19_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI44RU_5_LC_15_19_1  (
            .in0(N__58044),
            .in1(N__71939),
            .in2(_gnd_net_),
            .in3(N__58346),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_1_0 ),
            .ltout(\dron_frame_decoder_1.un1_sink_data_valid_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_9_LC_15_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_9_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_9_LC_15_19_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_9_LC_15_19_2  (
            .in0(N__71946),
            .in1(N__58005),
            .in2(N__57927),
            .in3(N__61542),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83969),
            .ce(),
            .sr(N__77365));
    defparam \dron_frame_decoder_1.source_H_disp_side_4_LC_15_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_4_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_4_LC_15_19_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_4_LC_15_19_4  (
            .in0(N__58560),
            .in1(N__58349),
            .in2(N__71971),
            .in3(N__65221),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83969),
            .ce(),
            .sr(N__77365));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI7OL8_4_LC_15_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI7OL8_4_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI7OL8_4_LC_15_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNI7OL8_4_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58559),
            .lcout(drone_H_disp_side_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_19_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_15_19_6  (
            .in0(N__58347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77604),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_LC_15_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_15_19_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_15_19_7  (
            .in0(N__58513),
            .in1(N__58348),
            .in2(_gnd_net_),
            .in3(N__67312),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83969),
            .ce(),
            .sr(N__77365));
    defparam \pid_side.error_cry_7_c_RNIIEI03_LC_15_20_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIIEI03_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIIEI03_LC_15_20_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_side.error_cry_7_c_RNIIEI03_LC_15_20_0  (
            .in0(N__72272),
            .in1(N__70984),
            .in2(N__71148),
            .in3(N__70907),
            .lcout(),
            .ltout(\pid_side.m45_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNIVS265_LC_15_20_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNIVS265_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIVS265_LC_15_20_1 .LUT_INIT=16'b1101000011010011;
    LogicCell40 \pid_side.error_cry_9_c_RNIVS265_LC_15_20_1  (
            .in0(N__70041),
            .in1(N__73535),
            .in2(N__58206),
            .in3(N__70825),
            .lcout(\pid_side.N_46_1 ),
            .ltout(\pid_side.N_46_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_20_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_20_2 .LUT_INIT=16'b1000000011110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_23_LC_15_20_2  (
            .in0(N__70705),
            .in1(N__70497),
            .in2(N__58203),
            .in3(N__70042),
            .lcout(\pid_side.m27_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNIEOQK9_LC_15_20_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNIEOQK9_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIEOQK9_LC_15_20_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_cry_9_c_RNIEOQK9_LC_15_20_3  (
            .in0(N__70704),
            .in1(_gnd_net_),
            .in2(N__58683),
            .in3(N__58193),
            .lcout(\pid_side.N_50_1 ),
            .ltout(\pid_side.N_50_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_11_LC_15_20_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_11_LC_15_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_11_LC_15_20_4 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \pid_side.error_i_reg_esr_11_LC_15_20_4  (
            .in0(N__65449),
            .in1(N__70498),
            .in2(N__58182),
            .in3(N__58725),
            .lcout(\pid_side.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83985),
            .ce(N__69260),
            .sr(N__77369));
    defparam \pid_side.error_i_reg_esr_27_LC_15_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_27_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_27_LC_15_20_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_27_LC_15_20_5  (
            .in0(N__59239),
            .in1(N__58610),
            .in2(_gnd_net_),
            .in3(N__58713),
            .lcout(\pid_side.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83985),
            .ce(N__69260),
            .sr(N__77369));
    defparam \pid_side.error_i_reg_esr_19_LC_15_20_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_19_LC_15_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_19_LC_15_20_6 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \pid_side.error_i_reg_esr_19_LC_15_20_6  (
            .in0(N__58611),
            .in1(N__61892),
            .in2(_gnd_net_),
            .in3(N__58734),
            .lcout(\pid_side.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83985),
            .ce(N__69260),
            .sr(N__77369));
    defparam \pid_side.error_i_reg_esr_18_LC_15_21_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_18_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_18_LC_15_21_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_18_LC_15_21_0  (
            .in0(N__61891),
            .in1(N__61479),
            .in2(_gnd_net_),
            .in3(N__58572),
            .lcout(\pid_side.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84003),
            .ce(N__69304),
            .sr(N__77376));
    defparam \pid_side.error_cry_8_c_RNI9F7NB_LC_15_21_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNI9F7NB_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNI9F7NB_LC_15_21_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_cry_8_c_RNI9F7NB_LC_15_21_1  (
            .in0(N__70703),
            .in1(N__70769),
            .in2(_gnd_net_),
            .in3(N__61941),
            .lcout(\pid_side.N_39_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIQCIS_LC_15_21_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIQCIS_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIQCIS_LC_15_21_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_0_c_RNIQCIS_LC_15_21_2  (
            .in0(N__72679),
            .in1(N__71668),
            .in2(_gnd_net_),
            .in3(N__73161),
            .lcout(),
            .ltout(\pid_side.N_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI59GD1_LC_15_21_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI59GD1_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI59GD1_LC_15_21_3 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \pid_side.error_cry_0_c_RNI59GD1_LC_15_21_3  (
            .in0(N__72211),
            .in1(N__71076),
            .in2(N__58581),
            .in3(N__69165),
            .lcout(\pid_side.m2_0_03_3_i_0 ),
            .ltout(\pid_side.m2_0_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_15_21_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_15_21_4 .LUT_INIT=16'b0100000001010001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_18_LC_15_21_4  (
            .in0(N__70502),
            .in1(N__66029),
            .in2(N__58578),
            .in3(N__62025),
            .lcout(),
            .ltout(\pid_side.m6_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_15_21_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_15_21_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_18_LC_15_21_5  (
            .in0(N__70082),
            .in1(N__69786),
            .in2(N__58575),
            .in3(N__69550),
            .lcout(\pid_side.error_i_reg_9_rn_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIJGME2_LC_15_22_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNIJGME2_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIJGME2_LC_15_22_0 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIJGME2_LC_15_22_0  (
            .in0(N__71585),
            .in1(N__72786),
            .in2(N__73305),
            .in3(N__72581),
            .lcout(),
            .ltout(\pid_side.m51_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNICQ2H4_LC_15_22_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNICQ2H4_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNICQ2H4_LC_15_22_1 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_cry_2_0_c_RNICQ2H4_LC_15_22_1  (
            .in0(N__72210),
            .in1(N__72503),
            .in2(N__58566),
            .in3(N__72344),
            .lcout(\pid_side.N_39_0 ),
            .ltout(\pid_side.N_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_15_22_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_15_22_2 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_19_LC_15_22_2  (
            .in0(N__66027),
            .in1(N__70379),
            .in2(N__58563),
            .in3(N__58879),
            .lcout(\pid_side.m7_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_15_22_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_15_22_3 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_19_LC_15_22_3  (
            .in0(N__69682),
            .in1(N__70081),
            .in2(N__69867),
            .in3(N__58740),
            .lcout(\pid_side.error_i_reg_9_rn_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIJPVK6_LC_15_22_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIJPVK6_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIJPVK6_LC_15_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIJPVK6_LC_15_22_4  (
            .in0(N__66028),
            .in1(N__58880),
            .in2(_gnd_net_),
            .in3(N__58864),
            .lcout(\pid_side.N_53_0 ),
            .ltout(\pid_side.N_53_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_15_22_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_15_22_5 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_27_LC_15_22_5  (
            .in0(N__69681),
            .in1(N__69816),
            .in2(N__58716),
            .in3(N__70080),
            .lcout(\pid_side.error_i_reg_9_rn_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNI11I87_LC_15_22_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNI11I87_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNI11I87_LC_15_22_6 .LUT_INIT=16'b0011101000110000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNI11I87_LC_15_22_6  (
            .in0(N__65737),
            .in1(N__58704),
            .in2(N__70494),
            .in3(N__58863),
            .lcout(\pid_side.m104_ns_sx ),
            .ltout(\pid_side.m104_ns_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_22_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_22_7 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_23_LC_15_22_7  (
            .in0(N__70380),
            .in1(N__65738),
            .in2(N__58686),
            .in3(N__58679),
            .lcout(\pid_side.m11_2_03_3_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_0_LC_15_23_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_0_LC_15_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_0_LC_15_23_0 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_0_LC_15_23_0  (
            .in0(N__70643),
            .in1(N__61690),
            .in2(N__62137),
            .in3(N__62048),
            .lcout(\pid_side.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_1_LC_15_23_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_1_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_1_LC_15_23_1 .LUT_INIT=16'b1100000001010000;
    LogicCell40 \pid_side.error_i_reg_esr_1_LC_15_23_1  (
            .in0(N__65076),
            .in1(N__65781),
            .in2(N__62140),
            .in3(N__70644),
            .lcout(\pid_side.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_2_LC_15_23_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_2_LC_15_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_2_LC_15_23_2 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_2_LC_15_23_2  (
            .in0(N__70645),
            .in1(N__58772),
            .in2(N__62138),
            .in3(N__62022),
            .lcout(\pid_side.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_3_LC_15_23_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_3_LC_15_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_3_LC_15_23_3 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \pid_side.error_i_reg_esr_3_LC_15_23_3  (
            .in0(N__70660),
            .in1(N__58881),
            .in2(N__62139),
            .in3(N__58866),
            .lcout(\pid_side.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_23_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_23_4 .LUT_INIT=16'b0010000000100011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_17_LC_15_23_4  (
            .in0(N__65780),
            .in1(N__70527),
            .in2(N__70696),
            .in3(N__65075),
            .lcout(),
            .ltout(\pid_side.m5_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_17_LC_15_23_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_17_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_17_LC_15_23_5 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_side.error_i_reg_esr_17_LC_15_23_5  (
            .in0(N__69861),
            .in1(N__69501),
            .in2(N__58833),
            .in3(N__65493),
            .lcout(\pid_side.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_23_LC_15_23_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_23_LC_15_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_23_LC_15_23_6 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_side.error_i_reg_esr_23_LC_15_23_6  (
            .in0(N__69500),
            .in1(N__58821),
            .in2(N__69954),
            .in3(N__58812),
            .lcout(\pid_side.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_24_LC_15_23_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_24_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_24_LC_15_23_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \pid_side.error_i_reg_esr_24_LC_15_23_7  (
            .in0(N__69625),
            .in1(N__62235),
            .in2(N__69914),
            .in3(N__61977),
            .lcout(\pid_side.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84035),
            .ce(N__69306),
            .sr(N__77387));
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_15_24_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_15_24_0 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_14_LC_15_24_0  (
            .in0(N__61937),
            .in1(N__70434),
            .in2(N__62023),
            .in3(N__65679),
            .lcout(\pid_side.m136_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI13NVA_LC_15_24_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI13NVA_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI13NVA_LC_15_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_4_c_RNI13NVA_LC_15_24_1  (
            .in0(N__65678),
            .in1(N__62012),
            .in2(_gnd_net_),
            .in3(N__61936),
            .lcout(\pid_side.N_110 ),
            .ltout(\pid_side.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_15_24_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_15_24_2 .LUT_INIT=16'b0100011100000011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_22_LC_15_24_2  (
            .in0(N__66039),
            .in1(N__70433),
            .in2(N__58776),
            .in3(N__58768),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_24_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_24_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_6_LC_15_24_3  (
            .in0(N__58767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66038),
            .lcout(\pid_side.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_15_24_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_15_24_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_15_24_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_15_24_4  (
            .in0(N__80308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84051),
            .ce(N__73403),
            .sr(N__77392));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_15_24_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_15_24_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_15_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80307),
            .lcout(xy_ki_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84051),
            .ce(N__73403),
            .sr(N__77392));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_24_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_24_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_15_24_6  (
            .in0(N__80310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84051),
            .ce(N__73403),
            .sr(N__77392));
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_15_24_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_15_24_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_15_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_2_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80309),
            .lcout(xy_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84051),
            .ce(N__73403),
            .sr(N__77392));
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_15_25_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_15_25_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_12_LC_15_25_0  (
            .in0(N__61691),
            .in1(N__70427),
            .in2(_gnd_net_),
            .in3(N__65680),
            .lcout(\pid_side.m0_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_6_LC_15_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_6_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_6_LC_15_25_2 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_6_LC_15_25_2  (
            .in0(N__70358),
            .in1(N__59169),
            .in2(N__65460),
            .in3(N__59022),
            .lcout(\pid_front.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84068),
            .ce(N__59336),
            .sr(N__77395));
    defparam \pid_front.error_cry_0_c_RNI7N6N4_LC_15_25_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI7N6N4_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI7N6N4_LC_15_25_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \pid_front.error_cry_0_c_RNI7N6N4_LC_15_25_3  (
            .in0(N__61738),
            .in1(N__61591),
            .in2(_gnd_net_),
            .in3(N__58992),
            .lcout(\pid_front.N_32_0 ),
            .ltout(\pid_front.N_32_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_8_LC_15_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_8_LC_15_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_8_LC_15_25_4 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_front.error_i_reg_esr_8_LC_15_25_4  (
            .in0(N__65456),
            .in1(N__70432),
            .in2(N__58956),
            .in3(N__58953),
            .lcout(\pid_front.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84068),
            .ce(N__59336),
            .sr(N__77395));
    defparam \pid_front.error_i_reg_esr_RNO_0_5_LC_15_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_5_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_5_LC_15_25_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_5_LC_15_25_5  (
            .in0(N__65682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58920),
            .lcout(),
            .ltout(\pid_front.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_5_LC_15_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_5_LC_15_25_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_5_LC_15_25_6 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_front.error_i_reg_esr_5_LC_15_25_6  (
            .in0(N__65452),
            .in1(N__70431),
            .in2(N__58893),
            .in3(N__58890),
            .lcout(\pid_front.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84068),
            .ce(N__59336),
            .sr(N__77395));
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_15_25_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_15_25_7 .LUT_INIT=16'b0000100000001101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_16_LC_15_25_7  (
            .in0(N__65681),
            .in1(N__61692),
            .in2(N__70501),
            .in3(N__62049),
            .lcout(\pid_side.m4_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_9_sn_27_LC_15_26_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_9_sn_27_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_9_sn_27_LC_15_26_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \pid_side.error_i_reg_9_sn_27_LC_15_26_0  (
            .in0(N__69853),
            .in1(N__69480),
            .in2(_gnd_net_),
            .in3(N__70360),
            .lcout(pid_side_error_i_reg_9_sn_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_26_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_15_26_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_6_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__61636),
            .in2(_gnd_net_),
            .in3(N__59198),
            .lcout(\pid_front.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_16_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_16_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_16_6_0  (
            .in0(N__63419),
            .in1(N__59163),
            .in2(_gnd_net_),
            .in3(N__59130),
            .lcout(\ppm_encoder_1.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGA_0_LC_16_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGA_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGA_0_LC_16_6_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGA_0_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__66420),
            .in2(_gnd_net_),
            .in3(N__59085),
            .lcout(),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI2RGAZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIVG551_1_LC_16_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIVG551_1_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIVG551_1_LC_16_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIVG551_1_LC_16_6_2  (
            .in0(N__59063),
            .in1(N__78230),
            .in2(N__59034),
            .in3(N__76565),
            .lcout(),
            .ltout(\ppm_encoder_1.throttle_m_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIFL0A6_1_LC_16_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIFL0A6_1_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIFL0A6_1_LC_16_6_3 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIFL0A6_1_LC_16_6_3  (
            .in0(N__63641),
            .in1(N__59957),
            .in2(N__59031),
            .in3(N__59028),
            .lcout(\ppm_encoder_1.throttle_RNIFL0A6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_6_4 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_16_6_4  (
            .in0(N__77646),
            .in1(N__62952),
            .in2(N__66432),
            .in3(N__76568),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83838),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_6_5 .LUT_INIT=16'b1111111101010010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_6_5  (
            .in0(N__76566),
            .in1(N__76151),
            .in2(N__62995),
            .in3(N__77647),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83838),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_6_6  (
            .in0(N__59739),
            .in1(N__62948),
            .in2(_gnd_net_),
            .in3(N__59625),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_16_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_16_6_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_16_6_7  (
            .in0(N__76567),
            .in1(N__63420),
            .in2(N__62994),
            .in3(N__77648),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83838),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNI2Q3U4_0_LC_16_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNI2Q3U4_0_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNI2Q3U4_0_LC_16_7_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ppm_encoder_1.aileron_RNI2Q3U4_0_LC_16_7_0  (
            .in0(N__59466),
            .in1(N__63143),
            .in2(N__67866),
            .in3(N__59475),
            .lcout(\ppm_encoder_1.aileron_RNI2Q3U4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_0_LC_16_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_0_LC_16_7_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_0_LC_16_7_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.aileron_0_LC_16_7_1  (
            .in0(N__62582),
            .in1(N__59787),
            .in2(_gnd_net_),
            .in3(N__59468),
            .lcout(\ppm_encoder_1.aileronZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83846),
            .ce(),
            .sr(N__77290));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_7_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__62581),
            .in2(_gnd_net_),
            .in3(N__77617),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_0_LC_16_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_0_LC_16_7_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_0_LC_16_7_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.elevator_0_LC_16_7_3  (
            .in0(N__59507),
            .in1(N__62591),
            .in2(_gnd_net_),
            .in3(N__59565),
            .lcout(\ppm_encoder_1.elevatorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83846),
            .ce(),
            .sr(N__77290));
    defparam \ppm_encoder_1.throttle_0_LC_16_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_16_7_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_16_7_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_16_7_4  (
            .in0(N__62590),
            .in1(N__59541),
            .in2(_gnd_net_),
            .in3(N__59491),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83846),
            .ce(),
            .sr(N__77290));
    defparam \ppm_encoder_1.throttle_RNIPLIG2_0_LC_16_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIPLIG2_0_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIPLIG2_0_LC_16_7_5 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIPLIG2_0_LC_16_7_5  (
            .in0(N__59506),
            .in1(N__63342),
            .in2(N__59493),
            .in3(N__63217),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0 ),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_16_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_16_7_6 .LUT_INIT=16'b0110110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_16_7_6  (
            .in0(N__59467),
            .in1(N__67862),
            .in2(N__59451),
            .in3(N__63144),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_16_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_16_7_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_16_7_7 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_16_7_7  (
            .in0(N__73890),
            .in1(N__74550),
            .in2(N__59742),
            .in3(N__74378),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83846),
            .ce(),
            .sr(N__77290));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_16_8_0  (
            .in0(N__63462),
            .in1(N__59638),
            .in2(_gnd_net_),
            .in3(N__59693),
            .lcout(\ppm_encoder_1.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIVRIG2_3_LC_16_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIVRIG2_3_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIVRIG2_3_LC_16_8_1 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIVRIG2_3_LC_16_8_1  (
            .in0(N__59692),
            .in1(N__63369),
            .in2(N__59640),
            .in3(N__63222),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNIE64U4_3_LC_16_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNIE64U4_3_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNIE64U4_3_LC_16_8_2 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \ppm_encoder_1.aileron_RNIE64U4_3_LC_16_8_2  (
            .in0(N__59620),
            .in1(N__66984),
            .in2(N__59730),
            .in3(N__63142),
            .lcout(\ppm_encoder_1.aileron_RNIE64U4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_3_LC_16_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_3_LC_16_8_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_3_LC_16_8_4 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_3_LC_16_8_4  (
            .in0(N__59727),
            .in1(N__59715),
            .in2(N__62719),
            .in3(N__59694),
            .lcout(\ppm_encoder_1.elevatorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83854),
            .ce(),
            .sr(N__77297));
    defparam \ppm_encoder_1.throttle_3_LC_16_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_16_8_5 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_16_8_5  (
            .in0(N__59639),
            .in1(N__59682),
            .in2(N__59670),
            .in3(N__62693),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83854),
            .ce(),
            .sr(N__77297));
    defparam \ppm_encoder_1.aileron_3_LC_16_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_3_LC_16_8_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_3_LC_16_8_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.aileron_3_LC_16_8_6  (
            .in0(N__59621),
            .in1(N__60222),
            .in2(N__62718),
            .in3(N__66789),
            .lcout(\ppm_encoder_1.aileronZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83854),
            .ce(),
            .sr(N__77297));
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_16_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_16_8_7 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_16_8_7  (
            .in0(N__63141),
            .in1(N__60740),
            .in2(N__59607),
            .in3(N__63370),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI112R2_10_LC_16_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI112R2_10_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI112R2_10_LC_16_9_1 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNI112R2_10_LC_16_9_1  (
            .in0(N__59985),
            .in1(N__59958),
            .in2(N__59868),
            .in3(N__63264),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIOVAA6_10_LC_16_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIOVAA6_10_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIOVAA6_10_LC_16_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIOVAA6_10_LC_16_9_2  (
            .in0(N__66585),
            .in1(_gnd_net_),
            .in2(N__59877),
            .in3(N__59874),
            .lcout(\ppm_encoder_1.elevator_RNIOVAA6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_16_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_16_9_3 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNI02LH2_10_LC_16_9_3  (
            .in0(N__59797),
            .in1(N__63161),
            .in2(N__59838),
            .in3(N__63371),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_16_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_16_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_16_9_4  (
            .in0(N__63499),
            .in1(N__59866),
            .in2(_gnd_net_),
            .in3(N__59836),
            .lcout(),
            .ltout(\ppm_encoder_1.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_16_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_16_9_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_16_9_5  (
            .in0(N__59798),
            .in1(_gnd_net_),
            .in2(N__59814),
            .in3(N__62998),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_10_LC_16_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_16_9_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_16_9_6  (
            .in0(N__60018),
            .in1(N__59997),
            .in2(N__62717),
            .in3(N__59799),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83864),
            .ce(),
            .sr(N__77308));
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_16_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_16_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_c_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__59783),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_16_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_16_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__66905),
            .in2(N__60374),
            .in3(N__59748),
            .lcout(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_0 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_16_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_16_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__66869),
            .in2(_gnd_net_),
            .in3(N__59745),
            .lcout(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_1 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_16_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_16_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__66785),
            .in2(N__60375),
            .in3(N__60213),
            .lcout(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_2 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_16_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_16_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__60210),
            .in2(_gnd_net_),
            .in3(N__60186),
            .lcout(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_3 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_16_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_16_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__60182),
            .in2(_gnd_net_),
            .in3(N__60150),
            .lcout(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_4 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_16_10_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_16_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__60143),
            .in2(N__60376),
            .in3(N__60108),
            .lcout(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_5 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_10_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__60101),
            .in2(_gnd_net_),
            .in3(N__60066),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__60063),
            .in2(_gnd_net_),
            .in3(N__60030),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__67673),
            .in2(_gnd_net_),
            .in3(N__60021),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__60014),
            .in2(_gnd_net_),
            .in3(N__59988),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__60803),
            .in2(_gnd_net_),
            .in3(N__60771),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__60845),
            .in2(_gnd_net_),
            .in3(N__60759),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__67478),
            .in2(N__60373),
            .in3(N__60750),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60747),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83884),
            .ce(N__60723),
            .sr(N__77322));
    defparam CONSTANT_ONE_LUT4_LC_16_11_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_16_11_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_16_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_16_12_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_16_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_16_12_0  (
            .in0(N__66887),
            .in1(N__66805),
            .in2(N__64225),
            .in3(N__66926),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_12_1 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_RNO_LC_16_12_1  (
            .in0(N__66925),
            .in1(N__66886),
            .in2(N__66809),
            .in3(N__63928),
            .lcout(\pid_side.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_16_12_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_16_12_2 .LUT_INIT=16'b0001000000010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIQVTS_0_LC_16_12_2  (
            .in0(N__63929),
            .in1(N__64010),
            .in2(N__63865),
            .in3(_gnd_net_),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_16_12_3 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_16_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_RNO_LC_16_12_3  (
            .in0(N__64212),
            .in1(N__64183),
            .in2(N__64163),
            .in3(N__63855),
            .lcout(\pid_side.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_16_12_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_16_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKLMT_10_LC_16_12_4  (
            .in0(N__64184),
            .in1(N__64159),
            .in2(N__64055),
            .in3(N__64100),
            .lcout(),
            .ltout(\pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_16_12_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_16_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_16_12_5  (
            .in0(N__64127),
            .in1(N__67518),
            .in2(N__60879),
            .in3(N__67694),
            .lcout(\pid_side.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_16_12_6 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_16_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_RNO_LC_16_12_6  (
            .in0(N__67693),
            .in1(N__64099),
            .in2(N__64054),
            .in3(N__64126),
            .lcout(\pid_side.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_12_LC_16_12_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_12_LC_16_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_12_LC_16_12_7 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \pid_side.source_pid_1_esr_12_LC_16_12_7  (
            .in0(N__64011),
            .in1(N__67648),
            .in2(N__67559),
            .in3(N__67519),
            .lcout(side_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83895),
            .ce(N__67457),
            .sr(N__67426));
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_16_13_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_16_13_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_16_13_0  (
            .in0(N__79083),
            .in1(N__60834),
            .in2(N__74976),
            .in3(N__60824),
            .lcout(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_16_13_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_16_13_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_16_13_1  (
            .in0(N__79562),
            .in1(_gnd_net_),
            .in2(N__60951),
            .in3(N__74262),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ),
            .ltout(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_16_13_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_16_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_16_13_2  (
            .in0(N__79082),
            .in1(N__63884),
            .in2(N__60828),
            .in3(N__60823),
            .lcout(\pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_3_LC_16_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_16_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_3_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79563),
            .lcout(\pid_side.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83904),
            .ce(N__81257),
            .sr(N__81140));
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_16_13_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_16_13_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_16_13_5  (
            .in0(N__67878),
            .in1(N__60939),
            .in2(_gnd_net_),
            .in3(N__60932),
            .lcout(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_16_13_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_16_13_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_16_13_6  (
            .in0(N__74261),
            .in1(N__60947),
            .in2(_gnd_net_),
            .in3(N__79561),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ),
            .ltout(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_16_13_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_16_13_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI7U286_2_LC_16_13_7  (
            .in0(N__67877),
            .in1(N__60931),
            .in2(N__60912),
            .in3(N__75660),
            .lcout(\pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_16_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_16_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_16_14_0  (
            .in0(N__79043),
            .in1(N__79064),
            .in2(_gnd_net_),
            .in3(N__68693),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITHHEA_12_LC_16_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITHHEA_12_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITHHEA_12_LC_16_14_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITHHEA_12_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60909),
            .in3(N__60983),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITHHEAZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_16_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_16_14_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_16_14_2  (
            .in0(N__78999),
            .in1(N__79014),
            .in2(_gnd_net_),
            .in3(N__60900),
            .lcout(\pid_side.un1_pid_prereg_0_2 ),
            .ltout(\pid_side.un1_pid_prereg_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_16_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_16_14_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_16_14_3  (
            .in0(N__61014),
            .in1(N__60996),
            .in2(N__60906),
            .in3(N__67808),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_16_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_16_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_16_14_4  (
            .in0(N__79449),
            .in1(N__79470),
            .in2(_gnd_net_),
            .in3(N__67997),
            .lcout(\pid_side.un1_pid_prereg_0_3 ),
            .ltout(\pid_side.un1_pid_prereg_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_16_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_16_14_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60903),
            .in3(N__67826),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_16_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_16_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_16_14_6  (
            .in0(N__78998),
            .in1(N__79013),
            .in2(_gnd_net_),
            .in3(N__60899),
            .lcout(\pid_side.un1_pid_prereg_0_1 ),
            .ltout(\pid_side.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_16_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_16_14_7 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__61010),
            .in2(N__61017),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_16_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_16_15_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_16_15_0  (
            .in0(N__79047),
            .in1(N__79071),
            .in2(_gnd_net_),
            .in3(N__68692),
            .lcout(\pid_side.un1_pid_prereg_0_0 ),
            .ltout(\pid_side.un1_pid_prereg_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIJ1F8F_12_LC_16_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIJ1F8F_12_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIJ1F8F_12_LC_16_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIJ1F8F_12_LC_16_15_1  (
            .in0(N__60972),
            .in1(N__60984),
            .in2(N__60999),
            .in3(N__60995),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIJ1F8FZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMEJ18_12_LC_16_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMEJ18_12_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMEJ18_12_LC_16_15_2 .LUT_INIT=16'b1111101011101000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMEJ18_12_LC_16_15_2  (
            .in0(N__79323),
            .in1(N__79380),
            .in2(N__79353),
            .in3(N__61068),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIMEJ18Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINPDOK_12_LC_16_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINPDOK_12_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINPDOK_12_LC_16_15_3 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINPDOK_12_LC_16_15_3  (
            .in0(N__78918),
            .in1(N__60971),
            .in2(N__60960),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNINPDOKZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_16_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_16_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__61085),
            .in2(_gnd_net_),
            .in3(N__61274),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIG7B43_12_LC_16_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIG7B43_12_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIG7B43_12_LC_16_15_6 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIG7B43_12_LC_16_15_6  (
            .in0(N__81312),
            .in1(N__82644),
            .in2(_gnd_net_),
            .in3(N__78489),
            .lcout(),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIG7B43Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI83KO4_12_LC_16_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI83KO4_12_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI83KO4_12_LC_16_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI83KO4_12_LC_16_15_7  (
            .in0(N__78964),
            .in1(_gnd_net_),
            .in2(N__60957),
            .in3(N__79422),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI83KO4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_16_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_16_16_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_16_16_0  (
            .in0(N__80834),
            .in1(N__81574),
            .in2(N__64734),
            .in3(N__64828),
            .lcout(\pid_side.un1_pid_prereg_0_19 ),
            .ltout(\pid_side.un1_pid_prereg_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_16_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_16_16_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60954),
            .in3(N__64778),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISG2C3_13_LC_16_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISG2C3_13_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISG2C3_13_LC_16_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISG2C3_13_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__79415),
            .in2(_gnd_net_),
            .in3(N__78485),
            .lcout(\pid_side.un1_pid_prereg_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_16_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_16_16_3 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_16_16_3  (
            .in0(N__81573),
            .in1(N__80833),
            .in2(N__64733),
            .in3(N__61038),
            .lcout(\pid_side.un1_pid_prereg_0_18 ),
            .ltout(\pid_side.un1_pid_prereg_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_16_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_16_16_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_16_16_4  (
            .in0(N__61134),
            .in1(N__61119),
            .in2(N__61062),
            .in3(N__64790),
            .lcout(\pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_16_5  (
            .in0(N__61395),
            .in1(N__65040),
            .in2(_gnd_net_),
            .in3(N__61055),
            .lcout(\pid_side.un1_pid_prereg_0_14 ),
            .ltout(\pid_side.un1_pid_prereg_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_16_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_16_6  (
            .in0(N__61151),
            .in1(N__61275),
            .in2(N__61059),
            .in3(N__61086),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__61150),
            .in2(_gnd_net_),
            .in3(N__61166),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_16_17_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_16_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_16_17_0  (
            .in0(N__61394),
            .in1(N__65039),
            .in2(_gnd_net_),
            .in3(N__61054),
            .lcout(\pid_side.un1_pid_prereg_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_17_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_17_1 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_17_1  (
            .in0(N__81591),
            .in1(N__80830),
            .in2(N__64730),
            .in3(N__61180),
            .lcout(\pid_side.un1_pid_prereg_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_16_17_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_16_17_2 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_16_17_2  (
            .in0(N__80832),
            .in1(N__81593),
            .in2(N__64732),
            .in3(N__61033),
            .lcout(\pid_side.un1_pid_prereg_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_17_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_17_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_16_17_3  (
            .in0(N__81966),
            .in1(N__82161),
            .in2(_gnd_net_),
            .in3(N__68212),
            .lcout(\pid_side.un1_pid_prereg_0_10 ),
            .ltout(\pid_side.un1_pid_prereg_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_16_17_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_16_17_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_16_17_4  (
            .in0(N__68478),
            .in1(N__61298),
            .in2(N__61185),
            .in3(N__68025),
            .lcout(\pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_16_17_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_16_17_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_16_17_5  (
            .in0(N__81592),
            .in1(N__80831),
            .in2(N__64731),
            .in3(N__61181),
            .lcout(\pid_side.un1_pid_prereg_0_16 ),
            .ltout(\pid_side.un1_pid_prereg_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_16_17_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_16_17_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_16_17_6  (
            .in0(N__61167),
            .in1(N__61155),
            .in2(N__61137),
            .in3(N__61132),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_16_17_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_16_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_16_17_7  (
            .in0(N__61133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61115),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_18_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_18_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_18_0  (
            .in0(N__61335),
            .in1(N__61360),
            .in2(N__61253),
            .in3(N__61359),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_16_18_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_16_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_16_18_1  (
            .in0(N__64649),
            .in1(N__67187),
            .in2(_gnd_net_),
            .in3(N__61099),
            .lcout(\pid_side.un1_pid_prereg_0_11 ),
            .ltout(\pid_side.un1_pid_prereg_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_16_18_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_16_18_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61104),
            .in3(N__61286),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_16_18_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_16_18_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_16_18_3  (
            .in0(N__64650),
            .in1(N__67188),
            .in2(_gnd_net_),
            .in3(N__61100),
            .lcout(\pid_side.un1_pid_prereg_0_12 ),
            .ltout(\pid_side.un1_pid_prereg_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_16_18_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_16_18_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_16_18_4  (
            .in0(N__61299),
            .in1(N__61287),
            .in2(N__61278),
            .in3(N__61267),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_18_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_18_5 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_side.pid_prereg_esr_RNO_0_30_LC_16_18_5  (
            .in0(N__61249),
            .in1(N__61361),
            .in2(N__61254),
            .in3(N__61362),
            .lcout(\pid_side.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_16_18_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_16_18_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_16_18_6  (
            .in0(N__61199),
            .in1(N__64806),
            .in2(N__64764),
            .in3(N__61213),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_18_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_18_7 .LUT_INIT=16'b1111101100100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_18_7  (
            .in0(N__80835),
            .in1(N__64729),
            .in2(N__81594),
            .in3(N__61378),
            .lcout(\pid_side.un1_pid_prereg_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_16_19_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_16_19_0 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_16_19_0  (
            .in0(N__80812),
            .in1(N__64727),
            .in2(N__81571),
            .in3(N__61228),
            .lcout(\pid_side.un1_pid_prereg_0_23 ),
            .ltout(\pid_side.un1_pid_prereg_0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_16_19_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_16_19_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61233),
            .in3(N__61214),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_16_19_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_16_19_2 .LUT_INIT=16'b1111101100100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_16_19_2  (
            .in0(N__80811),
            .in1(N__64726),
            .in2(N__81570),
            .in3(N__64861),
            .lcout(\pid_side.un1_pid_prereg_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_16_19_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_16_19_3 .LUT_INIT=16'b1010111010001010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_16_19_3  (
            .in0(N__61229),
            .in1(N__81543),
            .in2(N__64737),
            .in3(N__80813),
            .lcout(\pid_side.un1_pid_prereg_0_24 ),
            .ltout(\pid_side.un1_pid_prereg_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_16_19_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_16_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_16_19_4  (
            .in0(N__61215),
            .in1(N__61200),
            .in2(N__61188),
            .in3(N__61358),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_19_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_19_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_19_5  (
            .in0(N__64722),
            .in1(N__81542),
            .in2(_gnd_net_),
            .in3(N__80810),
            .lcout(\pid_side.un1_pid_prereg_370_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_16_19_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_16_19_6 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_16_19_6  (
            .in0(N__80814),
            .in1(N__64728),
            .in2(N__81572),
            .in3(N__61379),
            .lcout(\pid_side.un1_pid_prereg_0_25 ),
            .ltout(\pid_side.un1_pid_prereg_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_16_19_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_16_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__61338),
            .in3(N__61334),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIJGL43_LC_16_20_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNIJGL43_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIJGL43_LC_16_20_0 .LUT_INIT=16'b1010000110101011;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIJGL43_LC_16_20_0  (
            .in0(N__61323),
            .in1(N__72787),
            .in2(N__72269),
            .in3(N__72582),
            .lcout(\pid_side.N_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNIH0S81_LC_16_20_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNIH0S81_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNIH0S81_LC_16_20_1 .LUT_INIT=16'b0001001111010011;
    LogicCell40 \pid_side.error_cry_1_c_RNIH0S81_LC_16_20_1  (
            .in0(N__73054),
            .in1(N__71582),
            .in2(N__73299),
            .in3(N__73166),
            .lcout(\pid_side.m11_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIAA9L2_LC_16_20_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIAA9L2_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIAA9L2_LC_16_20_2 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIAA9L2_LC_16_20_2  (
            .in0(N__71583),
            .in1(N__72502),
            .in2(N__73303),
            .in3(N__72337),
            .lcout(),
            .ltout(\pid_side.m88_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNI0PMD4_LC_16_20_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI0PMD4_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI0PMD4_LC_16_20_3 .LUT_INIT=16'b1011000010110101;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI0PMD4_LC_16_20_3  (
            .in0(N__72246),
            .in1(N__69032),
            .in2(N__61317),
            .in3(N__72425),
            .lcout(\pid_side.N_89_0 ),
            .ltout(\pid_side.N_89_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIOVKQ7_LC_16_20_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIOVKQ7_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIOVKQ7_LC_16_20_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIOVKQ7_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__65746),
            .in2(N__61314),
            .in3(N__65066),
            .lcout(\pid_side.N_116_0 ),
            .ltout(\pid_side.N_116_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_16_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_16_20_5 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_13_LC_16_20_5  (
            .in0(N__69599),
            .in1(N__69868),
            .in2(N__61311),
            .in3(N__65601),
            .lcout(\pid_side.error_i_reg_9_rn_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNICTL8_9_LC_16_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNICTL8_9_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNICTL8_9_LC_16_20_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNICTL8_9_LC_16_20_7  (
            .in0(N__61541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_21_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_21_0 .LUT_INIT=16'b1000000011011111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_25_LC_16_21_0  (
            .in0(N__70411),
            .in1(N__65292),
            .in2(N__70732),
            .in3(N__70092),
            .lcout(),
            .ltout(\pid_side.m29_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_25_LC_16_21_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_25_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_25_LC_16_21_1 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_side.error_i_reg_esr_25_LC_16_21_1  (
            .in0(N__69851),
            .in1(N__69587),
            .in2(N__61530),
            .in3(N__65466),
            .lcout(\pid_side.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84021),
            .ce(N__69303),
            .sr(N__77382));
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_16_21_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_16_21_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_21_LC_16_21_2  (
            .in0(N__69586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70091),
            .lcout(\pid_side.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_16_21_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_16_21_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_5_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__65779),
            .in2(_gnd_net_),
            .in3(N__70698),
            .lcout(),
            .ltout(\pid_side.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_5_LC_16_21_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_5_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_5_LC_16_21_4 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \pid_side.error_i_reg_esr_5_LC_16_21_4  (
            .in0(N__65430),
            .in1(N__70512),
            .in2(N__61515),
            .in3(N__61512),
            .lcout(\pid_side.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84021),
            .ce(N__69303),
            .sr(N__77382));
    defparam \pid_side.error_i_reg_esr_10_LC_16_21_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_10_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_10_LC_16_21_5 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_10_LC_16_21_5  (
            .in0(N__70510),
            .in1(N__61488),
            .in2(N__65450),
            .in3(N__61477),
            .lcout(\pid_side.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84021),
            .ce(N__69303),
            .sr(N__77382));
    defparam \pid_side.error_i_reg_esr_4_LC_16_21_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_4_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_4_LC_16_21_6 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \pid_side.error_i_reg_esr_4_LC_16_21_6  (
            .in0(N__65429),
            .in1(N__63795),
            .in2(N__70496),
            .in3(N__62187),
            .lcout(\pid_side.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84021),
            .ce(N__69303),
            .sr(N__77382));
    defparam \pid_side.error_i_reg_esr_6_LC_16_21_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_6_LC_16_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_6_LC_16_21_7 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_6_LC_16_21_7  (
            .in0(N__70511),
            .in1(N__61431),
            .in2(N__65451),
            .in3(N__61422),
            .lcout(\pid_side.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84021),
            .ce(N__69303),
            .sr(N__77382));
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_16_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_16_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_0_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80514),
            .lcout(xy_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84036),
            .ce(N__73404),
            .sr(N__77388));
    defparam \pid_front.m12_1_LC_16_22_1 .C_ON=1'b0;
    defparam \pid_front.m12_1_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.m12_1_LC_16_22_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.m12_1_LC_16_22_1  (
            .in0(N__61805),
            .in1(N__71060),
            .in2(_gnd_net_),
            .in3(N__72992),
            .lcout(\pid_front.m0_0_03 ),
            .ltout(\pid_front.m0_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un4_error_i_reg_22_ns_1_LC_16_22_2 .C_ON=1'b0;
    defparam \pid_front.un4_error_i_reg_22_ns_1_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un4_error_i_reg_22_ns_1_LC_16_22_2 .LUT_INIT=16'b0001000100110001;
    LogicCell40 \pid_front.un4_error_i_reg_22_ns_1_LC_16_22_2  (
            .in0(N__69576),
            .in1(N__70295),
            .in2(N__61713),
            .in3(N__66030),
            .lcout(\pid_front.un4_error_i_reg_22_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_16_22_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_16_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73750),
            .lcout(xy_ki_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84036),
            .ce(N__73404),
            .sr(N__77388));
    defparam \pid_side.m12_1_LC_16_22_4 .C_ON=1'b0;
    defparam \pid_side.m12_1_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.m12_1_LC_16_22_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.m12_1_LC_16_22_4  (
            .in0(N__71059),
            .in1(N__72180),
            .in2(_gnd_net_),
            .in3(N__69142),
            .lcout(\pid_side.m0_0_03 ),
            .ltout(\pid_side.m0_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI6NL53_LC_16_22_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNI6NL53_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI6NL53_LC_16_22_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \pid_side.error_cry_2_c_RNI6NL53_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__61605),
            .in2(N__61548),
            .in3(N__62044),
            .lcout(\pid_side.N_32_0 ),
            .ltout(\pid_side.N_32_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_16_22_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_24_LC_16_22_6 .LUT_INIT=16'b1101000111110011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_24_LC_16_22_6  (
            .in0(N__70646),
            .in1(N__70296),
            .in2(N__61545),
            .in3(N__61963),
            .lcout(\pid_side.error_i_reg_esr_RNO_2Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_16_22_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_24_LC_16_22_7 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_24_LC_16_22_7  (
            .in0(N__61964),
            .in1(N__70647),
            .in2(N__70410),
            .in3(N__62216),
            .lcout(\pid_side.error_i_reg_esr_RNO_3Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNI4SA4A_LC_16_23_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNI4SA4A_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNI4SA4A_LC_16_23_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_cry_6_c_RNI4SA4A_LC_16_23_0  (
            .in0(N__65812),
            .in1(N__70615),
            .in2(_gnd_net_),
            .in3(N__61965),
            .lcout(\pid_side.N_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI8GMC2_LC_16_23_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNI8GMC2_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI8GMC2_LC_16_23_1 .LUT_INIT=16'b1111001100000101;
    LogicCell40 \pid_side.error_cry_2_c_RNI8GMC2_LC_16_23_1  (
            .in0(N__73053),
            .in1(N__72785),
            .in2(N__72219),
            .in3(N__65799),
            .lcout(\pid_side.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIIKRK2_LC_16_23_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNIIKRK2_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIIKRK2_LC_16_23_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIIKRK2_LC_16_23_2  (
            .in0(N__71558),
            .in1(N__72580),
            .in2(_gnd_net_),
            .in3(N__72501),
            .lcout(\pid_side.N_27_1 ),
            .ltout(\pid_side.N_27_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIGEO64_LC_16_23_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIGEO64_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIGEO64_LC_16_23_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_side.error_cry_2_c_RNIGEO64_LC_16_23_3  (
            .in0(N__72179),
            .in1(_gnd_net_),
            .in2(N__62028),
            .in3(N__65787),
            .lcout(\pid_side.N_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_16_23_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_16_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_24_LC_16_23_4  (
            .in0(N__65813),
            .in1(N__61989),
            .in2(_gnd_net_),
            .in3(N__61983),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIKEKT4_LC_16_23_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIKEKT4_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIKEKT4_LC_16_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIKEKT4_LC_16_23_5  (
            .in0(N__72178),
            .in1(N__61971),
            .in2(_gnd_net_),
            .in3(N__61950),
            .lcout(\pid_side.N_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIUCK52_LC_16_23_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIUCK52_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIUCK52_LC_16_23_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIUCK52_LC_16_23_6  (
            .in0(N__71557),
            .in1(N__72335),
            .in2(_gnd_net_),
            .in3(N__72411),
            .lcout(\pid_side.N_25_0 ),
            .ltout(\pid_side.N_25_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNICULG6_LC_16_23_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNICULG6_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNICULG6_LC_16_23_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \pid_side.error_cry_4_c_RNICULG6_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__65793),
            .in2(N__61944),
            .in3(N__65271),
            .lcout(\pid_side.N_38_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_24_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_16_24_0 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_16_LC_16_24_0  (
            .in0(N__69636),
            .in1(N__62253),
            .in2(N__69951),
            .in3(N__61923),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_16_LC_16_24_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_16_LC_16_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_16_LC_16_24_1 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \pid_side.error_i_reg_esr_16_LC_16_24_1  (
            .in0(N__62229),
            .in1(_gnd_net_),
            .in2(N__61917),
            .in3(N__61911),
            .lcout(\pid_side.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84069),
            .ce(N__69322),
            .sr(N__77396));
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_24_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_24_2 .LUT_INIT=16'b1011001100010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_16_LC_16_24_2  (
            .in0(N__73595),
            .in1(N__70089),
            .in2(N__66063),
            .in3(N__62247),
            .lcout(\pid_side.N_58_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIVV702_LC_16_24_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNIVV702_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIVV702_LC_16_24_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_8_c_RNIVV702_LC_16_24_3  (
            .in0(N__71116),
            .in1(N__70915),
            .in2(_gnd_net_),
            .in3(N__70823),
            .lcout(\pid_side.N_36_0 ),
            .ltout(\pid_side.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNITP583_LC_16_24_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNITP583_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNITP583_LC_16_24_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \pid_side.error_cry_10_c_RNITP583_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__73544),
            .in2(N__62241),
            .in3(N__70087),
            .lcout(\pid_side.N_57_0 ),
            .ltout(\pid_side.N_57_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_16_24_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_16_24_5 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_24_LC_16_24_5  (
            .in0(N__70090),
            .in1(N__70614),
            .in2(N__62238),
            .in3(N__70245),
            .lcout(\pid_side.error_i_reg_esr_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_16_24_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_16_24_6 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_21_LC_16_24_6  (
            .in0(N__70824),
            .in1(N__71117),
            .in2(N__73602),
            .in3(N__70088),
            .lcout(\pid_side.N_126_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_8_LC_16_24_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_8_LC_16_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_8_LC_16_24_7 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \pid_side.error_i_reg_esr_8_LC_16_24_7  (
            .in0(N__62228),
            .in1(N__70246),
            .in2(N__65457),
            .in3(N__62220),
            .lcout(\pid_side.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84069),
            .ce(N__69322),
            .sr(N__77396));
    defparam \pid_side.error_cry_2_c_RNIHL8M6_LC_16_25_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIHL8M6_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIHL8M6_LC_16_25_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_2_c_RNIHL8M6_LC_16_25_2  (
            .in0(N__65999),
            .in1(N__66075),
            .in2(_gnd_net_),
            .in3(N__72102),
            .lcout(\pid_side.N_60_0 ),
            .ltout(\pid_side.N_60_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_25_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_25_3 .LUT_INIT=16'b1000100000001010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_12_LC_16_25_3  (
            .in0(N__69886),
            .in1(N__62175),
            .in2(N__62169),
            .in3(N__69654),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_12_LC_16_25_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_12_LC_16_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_12_LC_16_25_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_side.error_i_reg_esr_12_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(N__62141),
            .in2(N__62070),
            .in3(N__62397),
            .lcout(\pid_side.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84082),
            .ce(N__69317),
            .sr(N__77400));
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_25_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_12_LC_16_25_5  (
            .in0(N__70616),
            .in1(N__65817),
            .in2(_gnd_net_),
            .in3(N__62403),
            .lcout(\pid_side.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_4_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_4_0  (
            .in0(N__62390),
            .in1(N__62318),
            .in2(N__62291),
            .in3(N__62367),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIL5IF_0_LC_17_4_4 .C_ON=1'b0;
    defparam \pid_side.state_RNIL5IF_0_LC_17_4_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIL5IF_0_LC_17_4_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIL5IF_0_LC_17_4_4  (
            .in0(_gnd_net_),
            .in1(N__67273),
            .in2(_gnd_net_),
            .in3(N__77586),
            .lcout(\pid_side.state_RNIL5IFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_17_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_17_4_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_17_4_6  (
            .in0(N__74602),
            .in1(_gnd_net_),
            .in2(N__76641),
            .in3(N__76270),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_17_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_17_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_17_4_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_17_4_7  (
            .in0(N__76269),
            .in1(N__76634),
            .in2(_gnd_net_),
            .in3(N__74603),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_17_LC_17_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_17_5_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_17_5_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_17_5_0  (
            .in0(N__74307),
            .in1(N__62319),
            .in2(N__66390),
            .in3(N__76640),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83839),
            .ce(),
            .sr(N__77280));
    defparam \ppm_encoder_1.pulses2count_18_LC_17_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_17_5_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_17_5_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_17_5_1  (
            .in0(N__76639),
            .in1(N__66389),
            .in2(N__77949),
            .in3(N__62306),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83839),
            .ce(),
            .sr(N__77280));
    defparam \ppm_encoder_1.pulses2count_16_LC_17_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_17_5_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_17_5_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_17_5_7  (
            .in0(N__76638),
            .in1(N__74604),
            .in2(N__62292),
            .in3(N__66385),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83839),
            .ce(),
            .sr(N__77280));
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_17_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_17_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_17_6_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_1_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__73726),
            .in2(_gnd_net_),
            .in3(N__83027),
            .lcout(xy_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83847),
            .ce(N__80912),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_17_7_0  (
            .in0(N__63463),
            .in1(N__62788),
            .in2(_gnd_net_),
            .in3(N__62846),
            .lcout(\ppm_encoder_1.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITPIG2_2_LC_17_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITPIG2_2_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITPIG2_2_LC_17_7_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNITPIG2_2_LC_17_7_1  (
            .in0(N__62845),
            .in1(N__63368),
            .in2(N__62790),
            .in3(N__63249),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_RNIA24U4_2_LC_17_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNIA24U4_2_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNIA24U4_2_LC_17_7_2 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \ppm_encoder_1.aileron_RNIA24U4_2_LC_17_7_2  (
            .in0(N__67010),
            .in1(N__62764),
            .in2(N__63168),
            .in3(N__63162),
            .lcout(\ppm_encoder_1.aileron_RNIA24U4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_17_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_17_7_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_17_7_3  (
            .in0(N__62765),
            .in1(N__63066),
            .in2(N__62997),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_2_LC_17_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_2_LC_17_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_2_LC_17_7_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_2_LC_17_7_4  (
            .in0(N__62886),
            .in1(N__62862),
            .in2(N__62850),
            .in3(N__62597),
            .lcout(\ppm_encoder_1.elevatorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83855),
            .ce(),
            .sr(N__77298));
    defparam \ppm_encoder_1.throttle_2_LC_17_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_17_7_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_17_7_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_17_7_5  (
            .in0(N__62789),
            .in1(N__62832),
            .in2(N__62673),
            .in3(N__62817),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83855),
            .ce(),
            .sr(N__77298));
    defparam \ppm_encoder_1.aileron_2_LC_17_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_2_LC_17_7_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_2_LC_17_7_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_2_LC_17_7_6  (
            .in0(N__62766),
            .in1(N__62593),
            .in2(N__66873),
            .in3(N__62775),
            .lcout(\ppm_encoder_1.aileronZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83855),
            .ce(),
            .sr(N__77298));
    defparam \ppm_encoder_1.rudder_6_LC_17_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_17_7_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_17_7_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_17_7_7  (
            .in0(N__62592),
            .in1(N__62424),
            .in2(_gnd_net_),
            .in3(N__66142),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83855),
            .ce(),
            .sr(N__77298));
    defparam \ppm_encoder_1.aileron_RNI8VQU5_0_LC_17_8_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.aileron_RNI8VQU5_0_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNI8VQU5_0_LC_17_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.aileron_RNI8VQU5_0_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__63657),
            .in2(N__67861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_8_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__63651),
            .in2(N__63642),
            .in3(N__63606),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_8_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__63603),
            .in2(N__67011),
            .in3(N__63597),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_8_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__63594),
            .in2(N__66983),
            .in3(N__63588),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_8_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__63585),
            .in2(N__66951),
            .in3(N__63576),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_8_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__63573),
            .in2(N__66252),
            .in3(N__63564),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_8_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__63561),
            .in2(N__66167),
            .in3(N__63549),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_8_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__63546),
            .in2(N__63533),
            .in3(N__63507),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__63762),
            .in2(N__74069),
            .in3(N__63753),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__63750),
            .in2(N__73959),
            .in3(N__63741),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__63738),
            .in2(N__66581),
            .in3(N__63732),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__63729),
            .in2(N__66761),
            .in3(N__63720),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__63717),
            .in2(N__66710),
            .in3(N__63705),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__63702),
            .in2(N__66656),
            .in3(N__63690),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__74933),
            .in2(N__63687),
            .in3(N__63675),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__73800),
            .in2(N__63831),
            .in3(N__63672),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__63669),
            .in2(_gnd_net_),
            .in3(N__63660),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__63822),
            .in2(_gnd_net_),
            .in3(N__63837),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__73842),
            .in2(_gnd_net_),
            .in3(N__63834),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__76287),
            .in2(_gnd_net_),
            .in3(N__76563),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_17_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_17_10_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_17_10_7  (
            .in0(N__76564),
            .in1(_gnd_net_),
            .in2(N__76293),
            .in3(N__74299),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIIIOO_0_LC_17_11_4 .C_ON=1'b0;
    defparam \pid_side.state_RNIIIOO_0_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIIIOO_0_LC_17_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.state_RNIIIOO_0_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__83001),
            .in2(_gnd_net_),
            .in3(N__78368),
            .lcout(\pid_side.state_RNIIIOOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_17_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_4_LC_17_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_4_LC_17_11_6  (
            .in0(N__73594),
            .in1(N__71166),
            .in2(N__70755),
            .in3(N__69164),
            .lcout(\pid_side.N_61_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_14_LC_17_12_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_14_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_14_LC_17_12_0 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_side.pid_prereg_14_LC_17_12_0  (
            .in0(N__63977),
            .in1(N__78462),
            .in2(N__67272),
            .in3(N__64395),
            .lcout(\pid_side.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83905),
            .ce(),
            .sr(N__77337));
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_17_12_1 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_17_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_RNO_LC_17_12_1  (
            .in0(N__67517),
            .in1(N__63976),
            .in2(N__64018),
            .in3(N__64376),
            .lcout(\pid_side.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_4_c_RNO_LC_17_12_2 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_4_c_RNO_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_4_c_RNO_LC_17_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_4_c_RNO_LC_17_12_2  (
            .in0(N__64292),
            .in1(N__64316),
            .in2(N__64278),
            .in3(N__64346),
            .lcout(\pid_side.un11lto30_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIE1A2_17_LC_17_12_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIE1A2_17_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIE1A2_17_LC_17_12_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIE1A2_17_LC_17_12_3  (
            .in0(N__64317),
            .in1(N__64277),
            .in2(_gnd_net_),
            .in3(N__64293),
            .lcout(),
            .ltout(\pid_side.pid_prereg_esr_RNIE1A2Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_17_12_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_17_12_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIAEHI_15_LC_17_12_4  (
            .in0(N__64377),
            .in1(N__63978),
            .in2(N__63963),
            .in3(N__64347),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_0_LC_17_12_7 .C_ON=1'b0;
    defparam \pid_side.state_0_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_0_LC_17_12_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.state_0_LC_17_12_7  (
            .in0(N__67370),
            .in1(N__67076),
            .in2(_gnd_net_),
            .in3(N__67260),
            .lcout(\pid_side.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83905),
            .ce(),
            .sr(N__77337));
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_13_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__81734),
            .in2(N__81741),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_0_LC_17_13_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_0_LC_17_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_0_LC_17_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_0_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__68427),
            .in2(N__68450),
            .in3(N__63915),
            .lcout(\pid_side.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_1_LC_17_13_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_1_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_1_LC_17_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_1_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__68113),
            .in2(N__68079),
            .in3(N__63912),
            .lcout(\pid_side.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_1 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_2_LC_17_13_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_2_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_2_LC_17_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_2_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__75330),
            .in2(N__75368),
            .in3(N__63909),
            .lcout(\pid_side.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_2 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_3_LC_17_13_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_3_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_3_LC_17_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_3_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__75659),
            .in2(N__63906),
            .in3(N__63894),
            .lcout(\pid_side.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_3 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_4_LC_17_13_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_4_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_4_LC_17_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_4_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__63891),
            .in2(N__63885),
            .in3(N__63840),
            .lcout(\pid_side.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_4 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_5_LC_17_13_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_5_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_5_LC_17_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_5_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__74972),
            .in2(N__64245),
            .in3(N__64191),
            .lcout(\pid_side.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_5 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_6_LC_17_13_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_6_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_6_LC_17_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_6_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__75033),
            .in2(N__75105),
            .in3(N__64170),
            .lcout(\pid_side.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_6 ),
            .clk(N__83916),
            .ce(N__78353),
            .sr(N__77342));
    defparam \pid_side.pid_prereg_esr_7_LC_17_14_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_7_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_7_LC_17_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_7_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__67017),
            .in2(N__75219),
            .in3(N__64137),
            .lcout(\pid_side.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_7 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_8_LC_17_14_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_8_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_8_LC_17_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_8_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__75126),
            .in2(N__75180),
            .in3(N__64107),
            .lcout(\pid_side.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_8 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_9_LC_17_14_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_9_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_9_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_9_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__75558),
            .in2(N__75578),
            .in3(N__64104),
            .lcout(\pid_side.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_9 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_10_LC_17_14_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_10_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_10_LC_17_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_10_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__75384),
            .in2(N__75516),
            .in3(N__64074),
            .lcout(\pid_side.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_10 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_11_LC_17_14_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_11_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_11_LC_17_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_11_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__68165),
            .in2(N__64071),
            .in3(N__64026),
            .lcout(\pid_side.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_11 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_12_LC_17_14_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_12_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_12_LC_17_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_12_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__68121),
            .in2(N__67905),
            .in3(N__63981),
            .lcout(\pid_side.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_12 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.pid_prereg_esr_13_LC_17_14_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_13_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_13_LC_17_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_13_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__67952),
            .in2(N__67941),
            .in3(N__64398),
            .lcout(\pid_side.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_13 ),
            .clk(N__83929),
            .ce(N__78355),
            .sr(N__77348));
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_14_7 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__78458),
            .in2(_gnd_net_),
            .in3(N__64386),
            .lcout(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_15_LC_17_15_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_15_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_15_LC_17_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_15_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__64383),
            .in2(N__78917),
            .in3(N__64365),
            .lcout(\pid_side.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_15 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_16_LC_17_15_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_16_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_16_LC_17_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_16_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__64362),
            .in2(N__64356),
            .in3(N__64335),
            .lcout(\pid_side.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_16 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_17_LC_17_15_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_17_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_17_LC_17_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_17_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__64332),
            .in2(N__64326),
            .in3(N__64305),
            .lcout(\pid_side.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_17 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_18_LC_17_15_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_18_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_18_LC_17_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_18_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__67797),
            .in2(N__64302),
            .in3(N__64281),
            .lcout(\pid_side.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_18 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_19_LC_17_15_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_19_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_19_LC_17_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_19_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__67767),
            .in2(N__67788),
            .in3(N__64263),
            .lcout(\pid_side.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_19 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_20_LC_17_15_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_20_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_20_LC_17_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_20_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__68004),
            .in2(N__68034),
            .in3(N__64248),
            .lcout(\pid_side.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_20 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_21_LC_17_15_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_21_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_21_LC_17_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_21_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__64641),
            .in2(N__68460),
            .in3(N__64617),
            .lcout(\pid_side.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_21 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_22_LC_17_15_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_22_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_22_LC_17_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_22_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__64614),
            .in2(N__64605),
            .in3(N__64581),
            .lcout(\pid_side.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_22 ),
            .clk(N__83942),
            .ce(N__78357),
            .sr(N__77353));
    defparam \pid_side.pid_prereg_esr_23_LC_17_16_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_23_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_23_LC_17_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_23_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__64578),
            .in2(N__64572),
            .in3(N__64548),
            .lcout(\pid_side.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_23 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_24_LC_17_16_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_24_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_24_LC_17_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_24_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__64545),
            .in2(N__64539),
            .in3(N__64518),
            .lcout(\pid_side.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_24 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_25_LC_17_16_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_25_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_25_LC_17_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_25_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__64515),
            .in2(N__64509),
            .in3(N__64488),
            .lcout(\pid_side.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_25 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_26_LC_17_16_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_26_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_26_LC_17_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_26_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__64743),
            .in2(N__64485),
            .in3(N__64464),
            .lcout(\pid_side.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_26 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_27_LC_17_16_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_27_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_27_LC_17_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_27_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__64461),
            .in2(N__64842),
            .in3(N__64437),
            .lcout(\pid_side.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_27 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_28_LC_17_16_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_28_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_28_LC_17_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_28_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__64434),
            .in2(N__64425),
            .in3(N__64401),
            .lcout(\pid_side.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_28 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_29_LC_17_16_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_29_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_29_LC_17_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_29_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__64920),
            .in2(N__64911),
            .in3(N__64884),
            .lcout(\pid_side.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_29 ),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.pid_prereg_esr_30_LC_17_16_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_30_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_30_LC_17_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.pid_prereg_esr_30_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__64881),
            .in2(_gnd_net_),
            .in3(N__64872),
            .lcout(\pid_side.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83957),
            .ce(N__78360),
            .sr(N__77360));
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_17_17_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_17_17_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_17_17_0  (
            .in0(N__81586),
            .in1(N__80809),
            .in2(N__64736),
            .in3(N__64869),
            .lcout(\pid_side.un1_pid_prereg_0_21 ),
            .ltout(\pid_side.un1_pid_prereg_0_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_17_17_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_17_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__64845),
            .in3(N__64802),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_17_17_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_17_17_2 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_17_17_2  (
            .in0(N__81585),
            .in1(N__80808),
            .in2(N__64735),
            .in3(N__64833),
            .lcout(\pid_side.un1_pid_prereg_0_20 ),
            .ltout(\pid_side.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_17_17_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_17_17_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_17_17_3  (
            .in0(N__64791),
            .in1(N__64779),
            .in2(N__64767),
            .in3(N__64754),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_22_LC_17_17_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_22_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_22_LC_17_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_22_LC_17_17_4  (
            .in0(N__81587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83970),
            .ce(N__81258),
            .sr(N__81138));
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_17_17_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_17_17_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_17_17_5  (
            .in0(N__80806),
            .in1(N__65048),
            .in2(_gnd_net_),
            .in3(N__82513),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_21_LC_17_17_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_17_17_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_21_LC_17_17_6  (
            .in0(N__82515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83970),
            .ce(N__81258),
            .sr(N__81138));
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_17_17_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_17_17_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_17_17_7  (
            .in0(N__80807),
            .in1(N__65049),
            .in2(_gnd_net_),
            .in3(N__82514),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_17_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_17_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80471),
            .lcout(side_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_17_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_17_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_17_18_1  (
            .in0(N__73725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(side_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_17_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_17_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80295),
            .lcout(side_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_17_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_17_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79716),
            .lcout(side_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_17_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_17_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80081),
            .lcout(side_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_17_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_17_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81102),
            .lcout(side_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_17_18_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_17_18_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_17_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79889),
            .lcout(side_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83986),
            .ce(N__65027),
            .sr(N__77370));
    defparam \dron_frame_decoder_1.source_H_disp_side_11_LC_17_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_11_LC_17_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_11_LC_17_19_0 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_11_LC_17_19_0  (
            .in0(N__65259),
            .in1(N__71972),
            .in2(N__71751),
            .in3(N__64996),
            .lcout(drone_H_disp_side_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84004),
            .ce(),
            .sr(N__77377));
    defparam \pid_side.error_axb_7_LC_17_19_1 .C_ON=1'b0;
    defparam \pid_side.error_axb_7_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_7_LC_17_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_axb_7_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__65243),
            .in2(_gnd_net_),
            .in3(N__65257),
            .lcout(\pid_side.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_8_l_ofx_LC_17_19_2 .C_ON=1'b0;
    defparam \pid_side.error_axb_8_l_ofx_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_8_l_ofx_LC_17_19_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_side.error_axb_8_l_ofx_LC_17_19_2  (
            .in0(N__65258),
            .in1(_gnd_net_),
            .in2(N__65247),
            .in3(N__68942),
            .lcout(\pid_side.error_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_12_LC_17_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_12_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_12_LC_17_19_3 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_12_LC_17_19_3  (
            .in0(N__68941),
            .in1(N__71728),
            .in2(N__71984),
            .in3(N__65231),
            .lcout(drone_H_disp_side_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84004),
            .ce(),
            .sr(N__77377));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIMF9E_12_LC_17_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIMF9E_12_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIMF9E_12_LC_17_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNIMF9E_12_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68940),
            .lcout(drone_H_disp_side_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_15_LC_17_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_15_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_15_LC_17_19_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_15_LC_17_19_5  (
            .in0(N__71976),
            .in1(N__65124),
            .in2(N__68880),
            .in3(N__71729),
            .lcout(drone_H_disp_side_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84004),
            .ce(),
            .sr(N__77377));
    defparam \dron_frame_decoder_1.source_H_disp_side_7_LC_17_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_7_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_7_LC_17_19_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_7_LC_17_19_6  (
            .in0(N__65085),
            .in1(N__71977),
            .in2(N__71752),
            .in3(N__65125),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84004),
            .ce(),
            .sr(N__77377));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIARL8_7_LC_17_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIARL8_7_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIARL8_7_LC_17_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNIARL8_7_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65084),
            .lcout(drone_H_disp_side_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNI5MBC4_LC_17_20_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNI5MBC4_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNI5MBC4_LC_17_20_0 .LUT_INIT=16'b0111001101000011;
    LogicCell40 \pid_side.error_cry_0_0_c_RNI5MBC4_LC_17_20_0  (
            .in0(N__65778),
            .in1(N__65744),
            .in2(N__70415),
            .in3(N__65065),
            .lcout(\pid_side.m93_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNIGQK82_LC_17_20_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNIGQK82_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIGQK82_LC_17_20_1 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \pid_side.error_cry_9_c_RNIGQK82_LC_17_20_1  (
            .in0(N__72244),
            .in1(N__70012),
            .in2(N__71150),
            .in3(N__70808),
            .lcout(\pid_side.N_126 ),
            .ltout(\pid_side.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_17_20_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_17_20_2 .LUT_INIT=16'b0000001111101110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_17_LC_17_20_2  (
            .in0(N__70013),
            .in1(N__70312),
            .in2(N__65499),
            .in3(N__65745),
            .lcout(),
            .ltout(\pid_side.m131_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_17_20_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_17_20_3 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_17_LC_17_20_3  (
            .in0(N__65304),
            .in1(N__70308),
            .in2(N__65496),
            .in3(N__65481),
            .lcout(\pid_side.m21_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIDGRBE_LC_17_20_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIDGRBE_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIDGRBE_LC_17_20_4 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \pid_side.error_cry_7_c_RNIDGRBE_LC_17_20_4  (
            .in0(N__65480),
            .in1(N__65303),
            .in2(N__70416),
            .in3(N__65472),
            .lcout(\pid_side.m13_2_03_4_i_0 ),
            .ltout(\pid_side.m13_2_03_4_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_9_LC_17_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_9_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_9_LC_17_20_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \pid_side.error_i_reg_9_LC_17_20_5  (
            .in0(N__65384),
            .in1(N__67217),
            .in2(N__65328),
            .in3(N__65318),
            .lcout(\pid_side.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84022),
            .ce(),
            .sr(N__77383));
    defparam \pid_side.error_cry_7_c_RNI13LC5_LC_17_20_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNI13LC5_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNI13LC5_LC_17_20_6 .LUT_INIT=16'b1010101000011011;
    LogicCell40 \pid_side.error_cry_7_c_RNI13LC5_LC_17_20_6  (
            .in0(N__71337),
            .in1(N__70966),
            .in2(N__70914),
            .in3(N__72245),
            .lcout(\pid_side.N_88_0 ),
            .ltout(\pid_side.N_88_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_20_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_20_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_13_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__70742),
            .in2(N__65295),
            .in3(N__65291),
            .lcout(\pid_side.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNINOG52_1_LC_17_21_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNINOG52_1_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNINOG52_1_LC_17_21_0 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_side.error_cry_4_c_RNINOG52_1_LC_17_21_0  (
            .in0(N__71541),
            .in1(N__69016),
            .in2(N__72220),
            .in3(N__71302),
            .lcout(\pid_side.error_cry_4_c_RNINOG52Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_8_20_LC_17_21_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_8_20_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_8_20_LC_17_21_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_8_20_LC_17_21_1  (
            .in0(N__71089),
            .in1(N__70894),
            .in2(_gnd_net_),
            .in3(N__70807),
            .lcout(),
            .ltout(\pid_side.N_36_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_17_21_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_17_21_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_20_LC_17_21_2  (
            .in0(N__73505),
            .in1(_gnd_net_),
            .in2(N__65262),
            .in3(N__70038),
            .lcout(\pid_side.N_57_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_17_21_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_17_21_3 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_7_20_LC_17_21_3  (
            .in0(N__71303),
            .in1(N__73506),
            .in2(N__69036),
            .in3(N__71127),
            .lcout(),
            .ltout(\pid_side.g0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_17_21_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_17_21_4 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_20_LC_17_21_4  (
            .in0(N__73507),
            .in1(N__71212),
            .in2(N__65550),
            .in3(N__70967),
            .lcout(),
            .ltout(\pid_side.N_22_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_17_21_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_17_21_5 .LUT_INIT=16'b1100111011011111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_20_LC_17_21_5  (
            .in0(N__70731),
            .in1(N__69601),
            .in2(N__65547),
            .in3(N__65544),
            .lcout(),
            .ltout(\pid_side.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_20_LC_17_21_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_20_LC_17_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_20_LC_17_21_6 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_side.error_i_reg_esr_20_LC_17_21_6  (
            .in0(N__65517),
            .in1(N__69952),
            .in2(N__65538),
            .in3(N__65895),
            .lcout(\pid_side.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84037),
            .ce(N__69299),
            .sr(N__77389));
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_17_21_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_17_21_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_20_LC_17_21_7  (
            .in0(N__70039),
            .in1(N__69600),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_17_22_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_17_22_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_12_21_LC_17_22_0  (
            .in0(N__73254),
            .in1(N__72488),
            .in2(N__72708),
            .in3(N__72336),
            .lcout(),
            .ltout(\pid_side.m88_0_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_17_22_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_17_22_1 .LUT_INIT=16'b1111000001010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_9_21_LC_17_22_1  (
            .in0(N__69040),
            .in1(N__72421),
            .in2(N__65511),
            .in3(N__72983),
            .lcout(\pid_side.N_89_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNI7FAB2_LC_17_22_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI7FAB2_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI7FAB2_LC_17_22_2 .LUT_INIT=16'b0001101101010101;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI7FAB2_LC_17_22_2  (
            .in0(N__71526),
            .in1(N__69037),
            .in2(N__72430),
            .in3(N__73206),
            .lcout(\pid_side.m48_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNINOG52_0_LC_17_22_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNINOG52_0_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNINOG52_0_LC_17_22_3 .LUT_INIT=16'b0100001101001111;
    LogicCell40 \pid_side.error_cry_4_c_RNINOG52_0_LC_17_22_3  (
            .in0(N__69039),
            .in1(N__72187),
            .in2(N__71577),
            .in3(N__71310),
            .lcout(),
            .ltout(\pid_side.m21_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIAGI15_LC_17_22_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNIAGI15_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIAGI15_LC_17_22_4 .LUT_INIT=16'b1100000111110001;
    LogicCell40 \pid_side.error_cry_6_c_RNIAGI15_LC_17_22_4  (
            .in0(N__71223),
            .in1(N__72218),
            .in2(N__65820),
            .in3(N__70977),
            .lcout(\pid_side.N_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIDQP81_LC_17_22_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIDQP81_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIDQP81_LC_17_22_5 .LUT_INIT=16'b0001100100111011;
    LogicCell40 \pid_side.error_cry_0_c_RNIDQP81_LC_17_22_5  (
            .in0(N__73205),
            .in1(N__71525),
            .in2(N__71669),
            .in3(N__73136),
            .lcout(\pid_side.m30_1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNINOG52_LC_17_22_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNINOG52_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNINOG52_LC_17_22_6 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pid_side.error_cry_4_c_RNINOG52_LC_17_22_6  (
            .in0(N__71309),
            .in1(N__71553),
            .in2(N__72221),
            .in3(N__69038),
            .lcout(\pid_side.error_cry_4_c_RNINOGZ0Z52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIQCOE1_LC_17_22_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIQCOE1_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIQCOE1_LC_17_22_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_2_c_RNIQCOE1_LC_17_22_7  (
            .in0(N__71552),
            .in1(N__73055),
            .in2(_gnd_net_),
            .in3(N__72769),
            .lcout(\pid_side.N_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI6H9Q_LC_17_23_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI6H9Q_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI6H9Q_LC_17_23_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \pid_side.error_cry_0_c_RNI6H9Q_LC_17_23_0  (
            .in0(N__72209),
            .in1(N__71660),
            .in2(N__71109),
            .in3(N__69157),
            .lcout(\pid_side.m1_0_03 ),
            .ltout(\pid_side.m1_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_23_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_17_23_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_13_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__70252),
            .in2(N__65754),
            .in3(N__65736),
            .lcout(\pid_side.m1_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_17_23_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_17_23_2 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_21_LC_17_23_2  (
            .in0(N__71250),
            .in1(N__69653),
            .in2(N__70746),
            .in3(N__65589),
            .lcout(),
            .ltout(\pid_side.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_21_LC_17_23_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_21_LC_17_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_21_LC_17_23_3 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_side.error_i_reg_esr_21_LC_17_23_3  (
            .in0(N__65583),
            .in1(N__69929),
            .in2(N__65574),
            .in3(N__66102),
            .lcout(\pid_side.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84070),
            .ce(N__69321),
            .sr(N__77397));
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_17_23_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_17_23_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_21_LC_17_23_4  (
            .in0(N__65556),
            .in1(N__66044),
            .in2(_gnd_net_),
            .in3(N__71592),
            .lcout(),
            .ltout(\pid_side.N_116_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_17_23_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_17_23_5 .LUT_INIT=16'b0011000110111001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_21_LC_17_23_5  (
            .in0(N__69652),
            .in1(N__70253),
            .in2(N__66105),
            .in3(N__66093),
            .lcout(\pid_side.un4_error_i_reg_31_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_17_23_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_17_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_10_21_LC_17_23_6  (
            .in0(N__71064),
            .in1(N__71661),
            .in2(_gnd_net_),
            .in3(N__69158),
            .lcout(),
            .ltout(\pid_side.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_17_23_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_17_23_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_21_LC_17_23_7  (
            .in0(N__66043),
            .in1(_gnd_net_),
            .in2(N__66096),
            .in3(N__73488),
            .lcout(\pid_side.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIPFJ32_LC_17_24_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIPFJ32_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIPFJ32_LC_17_24_0 .LUT_INIT=16'b1010000110101011;
    LogicCell40 \pid_side.error_cry_2_c_RNIPFJ32_LC_17_24_0  (
            .in0(N__66087),
            .in1(N__73069),
            .in2(N__72270),
            .in3(N__72790),
            .lcout(\pid_side.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_17_24_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_17_24_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_20_LC_17_24_2  (
            .in0(N__69146),
            .in1(N__73487),
            .in2(N__66062),
            .in3(N__71149),
            .lcout(\pid_side.N_61_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_17_24_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_17_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_20_LC_17_24_4  (
            .in0(N__66034),
            .in1(N__72714),
            .in2(_gnd_net_),
            .in3(N__73314),
            .lcout(),
            .ltout(\pid_side.N_60_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_17_24_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_17_24_5 .LUT_INIT=16'b0111010000110011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_20_LC_17_24_5  (
            .in0(N__65904),
            .in1(N__70244),
            .in2(N__65898),
            .in3(N__69651),
            .lcout(\pid_side.un4_error_i_reg_30_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_17_25_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_17_25_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_17_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_3_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79734),
            .lcout(xy_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84091),
            .ce(N__73412),
            .sr(N__77402));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_6_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_18_6_5  (
            .in0(N__65886),
            .in1(N__78178),
            .in2(_gnd_net_),
            .in3(N__74625),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83856),
            .ce(N__65873),
            .sr(N__77299));
    defparam \ppm_encoder_1.init_pulses_5_LC_18_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_18_7_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_18_7_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_18_7_0  (
            .in0(N__74410),
            .in1(N__77823),
            .in2(N__74505),
            .in3(N__66258),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83865),
            .ce(),
            .sr(N__77309));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_18_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_18_7_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_18_7_1  (
            .in0(N__76491),
            .in1(_gnd_net_),
            .in2(N__76225),
            .in3(N__66227),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_7_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_7_2  (
            .in0(N__66226),
            .in1(N__76170),
            .in2(_gnd_net_),
            .in3(N__76492),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_7_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_7_3  (
            .in0(N__74898),
            .in1(N__66228),
            .in2(N__74785),
            .in3(N__66216),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_6_LC_18_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_18_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_18_7_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_18_7_4  (
            .in0(N__74411),
            .in1(N__77784),
            .in2(N__74506),
            .in3(N__66174),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83865),
            .ce(),
            .sr(N__77309));
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_18_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_18_7_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICBN01_6_LC_18_7_5  (
            .in0(N__76493),
            .in1(_gnd_net_),
            .in2(N__76226),
            .in3(N__74191),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_18_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_18_7_6 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_18_7_6  (
            .in0(N__74192),
            .in1(N__74899),
            .in2(N__66150),
            .in3(N__74770),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_18_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_18_7_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_18_7_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_18_7_7  (
            .in0(N__74507),
            .in1(N__74412),
            .in2(N__77763),
            .in3(N__66111),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83865),
            .ce(),
            .sr(N__77309));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_18_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_18_8_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_18_8_0  (
            .in0(N__76625),
            .in1(_gnd_net_),
            .in2(N__76284),
            .in3(N__66605),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_18_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_18_8_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_18_8_1  (
            .in0(N__66377),
            .in1(N__74154),
            .in2(_gnd_net_),
            .in3(N__76627),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_18_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_18_8_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_18_8_2  (
            .in0(N__74413),
            .in1(N__77703),
            .in2(N__66618),
            .in3(N__66615),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83874),
            .ce(),
            .sr(N__77316));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_18_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_18_8_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_10_LC_18_8_3  (
            .in0(N__66604),
            .in1(N__76254),
            .in2(_gnd_net_),
            .in3(N__76626),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_18_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_18_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_18_8_4  (
            .in0(N__66564),
            .in1(N__66528),
            .in2(N__66486),
            .in3(N__66437),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_153_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_15_LC_18_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_18_8_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_18_8_5  (
            .in0(N__73823),
            .in1(N__66326),
            .in2(N__66366),
            .in3(N__76628),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83874),
            .ce(),
            .sr(N__77316));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_18_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_18_8_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_18_8_6  (
            .in0(N__66363),
            .in1(N__66354),
            .in2(N__66327),
            .in3(N__66315),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_18_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_18_8_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_18_8_7  (
            .in0(N__74469),
            .in1(N__78009),
            .in2(N__66273),
            .in3(N__74414),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83874),
            .ce(),
            .sr(N__77316));
    defparam \ppm_encoder_1.init_pulses_11_LC_18_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_18_9_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_18_9_0 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_18_9_0  (
            .in0(N__77679),
            .in1(N__74385),
            .in2(N__74503),
            .in3(N__66264),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83885),
            .ce(),
            .sr(N__77323));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_18_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_18_9_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_18_9_1  (
            .in0(N__66733),
            .in1(N__76263),
            .in2(_gnd_net_),
            .in3(N__76633),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_9_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_18_9_2  (
            .in0(N__76630),
            .in1(_gnd_net_),
            .in2(N__76285),
            .in3(N__66734),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_12_LC_18_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_18_9_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_18_9_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_18_9_3  (
            .in0(N__74384),
            .in1(N__78096),
            .in2(N__74504),
            .in3(N__66720),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83885),
            .ce(),
            .sr(N__77323));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_18_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_18_9_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_18_9_4  (
            .in0(N__76631),
            .in1(_gnd_net_),
            .in2(N__76286),
            .in3(N__66679),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_18_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_18_9_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_18_9_5  (
            .in0(N__66680),
            .in1(N__76255),
            .in2(_gnd_net_),
            .in3(N__76629),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_18_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_18_9_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_18_9_6 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_18_9_6  (
            .in0(N__74473),
            .in1(N__78054),
            .in2(N__74421),
            .in3(N__66666),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83885),
            .ce(),
            .sr(N__77323));
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_18_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_18_9_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_18_9_7  (
            .in0(N__74212),
            .in1(N__76262),
            .in2(_gnd_net_),
            .in3(N__76632),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_18_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_18_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_18_10_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_18_10_0  (
            .in0(N__66633),
            .in1(N__74417),
            .in2(N__74562),
            .in3(N__77874),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83896),
            .ce(),
            .sr(N__77330));
    defparam \ppm_encoder_1.init_pulses_2_LC_18_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_18_10_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_18_10_1 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_18_10_1  (
            .in0(N__74415),
            .in1(N__75984),
            .in2(N__74563),
            .in3(N__66627),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83896),
            .ce(),
            .sr(N__77330));
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_18_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_18_10_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI87N01_2_LC_18_10_2  (
            .in0(N__74095),
            .in1(N__76246),
            .in2(_gnd_net_),
            .in3(N__76622),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_18_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_18_10_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_18_10_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_18_10_3  (
            .in0(N__74416),
            .in1(N__75963),
            .in2(N__74564),
            .in3(N__66993),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83896),
            .ce(),
            .sr(N__77330));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_18_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_18_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_3_LC_18_10_4  (
            .in0(N__76657),
            .in1(N__76250),
            .in2(_gnd_net_),
            .in3(N__76624),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_18_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_18_10_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_18_10_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_18_10_6  (
            .in0(N__74540),
            .in1(N__66960),
            .in2(N__77853),
            .in3(N__74418),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83896),
            .ce(),
            .sr(N__77330));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_18_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_18_10_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_18_10_7  (
            .in0(N__76623),
            .in1(_gnd_net_),
            .in2(N__76283),
            .in3(N__76306),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_1_LC_18_11_0 .C_ON=1'b0;
    defparam \pid_side.state_1_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_1_LC_18_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.state_1_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67261),
            .lcout(\pid_side.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83906),
            .ce(),
            .sr(N__77338));
    defparam \pid_side.source_pid_1_esr_1_LC_18_12_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_1_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_1_LC_18_12_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \pid_side.source_pid_1_esr_1_LC_18_12_0  (
            .in0(N__67644),
            .in1(N__66848),
            .in2(N__66930),
            .in3(N__67756),
            .lcout(side_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83917),
            .ce(N__67461),
            .sr(N__67427));
    defparam \pid_side.source_pid_1_esr_2_LC_18_12_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_2_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_2_LC_18_12_1 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \pid_side.source_pid_1_esr_2_LC_18_12_1  (
            .in0(N__66847),
            .in1(N__67647),
            .in2(N__67761),
            .in3(N__66888),
            .lcout(side_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83917),
            .ce(N__67461),
            .sr(N__67427));
    defparam \pid_side.source_pid_1_esr_3_LC_18_12_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_3_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_3_LC_18_12_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \pid_side.source_pid_1_esr_3_LC_18_12_2  (
            .in0(N__67645),
            .in1(N__66849),
            .in2(N__66810),
            .in3(N__67757),
            .lcout(side_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83917),
            .ce(N__67461),
            .sr(N__67427));
    defparam \pid_side.source_pid_1_esr_9_LC_18_12_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_9_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_9_LC_18_12_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_9_LC_18_12_3  (
            .in0(N__67752),
            .in1(N__67646),
            .in2(_gnd_net_),
            .in3(N__67698),
            .lcout(side_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83917),
            .ce(N__67461),
            .sr(N__67427));
    defparam \pid_side.source_pid_1_esr_13_LC_18_12_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_13_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_13_LC_18_12_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_13_LC_18_12_4  (
            .in0(N__67643),
            .in1(N__67560),
            .in2(_gnd_net_),
            .in3(N__67525),
            .lcout(side_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83917),
            .ce(N__67461),
            .sr(N__67427));
    defparam \pid_side.state_RNINK4U_0_LC_18_12_5 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_LC_18_12_5 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \pid_side.state_RNINK4U_0_LC_18_12_5  (
            .in0(N__67059),
            .in1(N__67369),
            .in2(N__67279),
            .in3(N__77605),
            .lcout(),
            .ltout(\pid_side.state_RNINK4UZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIK1B71_0_LC_18_12_6 .C_ON=1'b0;
    defparam \pid_side.state_RNIK1B71_0_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIK1B71_0_LC_18_12_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.state_RNIK1B71_0_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67392),
            .in3(N__83004),
            .lcout(\pid_side.N_513_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIQ7UK_0_LC_18_12_7 .C_ON=1'b0;
    defparam \pid_side.state_RNIQ7UK_0_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIQ7UK_0_LC_18_12_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.state_RNIQ7UK_0_LC_18_12_7  (
            .in0(N__67058),
            .in1(N__67368),
            .in2(_gnd_net_),
            .in3(N__67268),
            .lcout(\pid_side.state_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_18_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_18_13_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_18_13_0  (
            .in0(N__82011),
            .in1(N__81980),
            .in2(_gnd_net_),
            .in3(N__82487),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_20_LC_18_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_18_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_18_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_20_LC_18_13_1  (
            .in0(N__82488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83930),
            .ce(N__81243),
            .sr(N__81143));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_13_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_13_2  (
            .in0(N__67170),
            .in1(N__67077),
            .in2(_gnd_net_),
            .in3(N__77607),
            .lcout(\pid_side.error_i_acumm_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_13_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_13_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_13_3  (
            .in0(N__75093),
            .in1(N__75051),
            .in2(_gnd_net_),
            .in3(N__75080),
            .lcout(\pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_18_13_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_18_13_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5SNH3_7_LC_18_13_4  (
            .in0(N__75930),
            .in1(N__75192),
            .in2(_gnd_net_),
            .in3(N__75159),
            .lcout(\pid_side.error_p_reg_esr_RNI5SNH3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_18_13_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_18_13_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_2_LC_18_13_5  (
            .in0(N__75312),
            .in1(N__75287),
            .in2(_gnd_net_),
            .in3(N__78656),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_2_LC_18_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_18_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_18_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_2_LC_18_13_6  (
            .in0(N__78657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83930),
            .ce(N__81243),
            .sr(N__81143));
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_18_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_18_13_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI65N01_0_LC_18_13_7  (
            .in0(N__73935),
            .in1(N__76245),
            .in2(_gnd_net_),
            .in3(N__76621),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_18_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_18_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_18_14_0  (
            .in0(N__67830),
            .in1(N__67778),
            .in2(N__67815),
            .in3(N__67966),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_18_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_18_14_1  (
            .in0(N__79490),
            .in1(N__79121),
            .in2(_gnd_net_),
            .in3(N__68315),
            .lcout(\pid_side.un1_pid_prereg_0_5 ),
            .ltout(\pid_side.un1_pid_prereg_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_18_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_18_14_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__67791),
            .in3(N__67967),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_18_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_18_14_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_18_14_3  (
            .in0(N__79491),
            .in1(N__79122),
            .in2(_gnd_net_),
            .in3(N__68316),
            .lcout(\pid_side.un1_pid_prereg_0_6 ),
            .ltout(\pid_side.un1_pid_prereg_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_18_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_18_14_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_18_14_4  (
            .in0(N__68063),
            .in1(N__67779),
            .in2(N__67770),
            .in3(N__67968),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_18_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_18_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_18_14_5  (
            .in0(N__80615),
            .in1(N__80636),
            .in2(_gnd_net_),
            .in3(N__68269),
            .lcout(\pid_side.un1_pid_prereg_0_7 ),
            .ltout(\pid_side.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_18_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_18_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__68007),
            .in3(N__68048),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_18_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_18_14_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_18_14_7  (
            .in0(N__79445),
            .in1(N__79466),
            .in2(_gnd_net_),
            .in3(N__67996),
            .lcout(\pid_side.un1_pid_prereg_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI3AMCB_10_LC_18_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI3AMCB_10_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI3AMCB_10_LC_18_15_0 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI3AMCB_10_LC_18_15_0  (
            .in0(N__67931),
            .in1(N__67956),
            .in2(N__80571),
            .in3(N__67893),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI3AMCBZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIE3IM2_12_LC_18_15_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIE3IM2_12_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIE3IM2_12_LC_18_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIE3IM2_12_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__80567),
            .in2(_gnd_net_),
            .in3(N__67930),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIO56DB_10_LC_18_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIO56DB_10_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIO56DB_10_LC_18_15_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIO56DB_10_LC_18_15_2  (
            .in0(N__68130),
            .in1(N__68154),
            .in2(N__67908),
            .in3(N__67892),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIO56DBZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_18_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_18_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_18_15_3  (
            .in0(N__75469),
            .in1(N__75117),
            .in2(_gnd_net_),
            .in3(N__75483),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_18_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_18_15_4 .LUT_INIT=16'b1111101010110010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_18_15_4  (
            .in0(N__82112),
            .in1(N__75473),
            .in2(N__67896),
            .in3(N__78515),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_18_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_18_15_5 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_18_15_5  (
            .in0(N__78516),
            .in1(N__82113),
            .in2(N__75474),
            .in3(N__67884),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__68178),
            .in3(N__68152),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_18_15_7  (
            .in0(N__68153),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68129),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_1_LC_18_16_0  (
            .in0(N__81899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83971),
            .ce(N__81256),
            .sr(N__81139));
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_16_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI98EQ_1_LC_18_16_1  (
            .in0(N__78555),
            .in1(N__75621),
            .in2(_gnd_net_),
            .in3(N__81898),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_16_2 .LUT_INIT=16'b0101101000001111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_16_2  (
            .in0(N__81936),
            .in1(N__68115),
            .in2(N__68082),
            .in3(N__75642),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_16_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_16_3  (
            .in0(N__80619),
            .in1(N__80643),
            .in2(_gnd_net_),
            .in3(N__68276),
            .lcout(\pid_side.un1_pid_prereg_0_8 ),
            .ltout(\pid_side.un1_pid_prereg_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_16_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_16_4  (
            .in0(N__68067),
            .in1(N__68052),
            .in2(N__68037),
            .in3(N__68018),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_16_5  (
            .in0(N__81962),
            .in1(N__82157),
            .in2(_gnd_net_),
            .in3(N__68220),
            .lcout(\pid_side.un1_pid_prereg_0_9 ),
            .ltout(\pid_side.un1_pid_prereg_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_16_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__68481),
            .in3(N__68471),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_16_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_16_7  (
            .in0(N__75641),
            .in1(N__68451),
            .in2(_gnd_net_),
            .in3(N__81935),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_18_17_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_18_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_18_17_0  (
            .in0(N__68415),
            .in1(N__68666),
            .in2(N__68394),
            .in3(N__68231),
            .lcout(),
            .ltout(\pid_side.un10lto27_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_18_17_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_18_17_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__68322),
            .in2(N__68370),
            .in3(N__68367),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_18_17_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_18_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_18_17_2  (
            .in0(N__68189),
            .in1(N__68246),
            .in2(N__68346),
            .in3(N__68288),
            .lcout(\pid_side.un10lto27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_18_17_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_18_17_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_18_LC_18_17_3  (
            .in0(N__68314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83987),
            .ce(N__78361),
            .sr(N__77371));
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_18_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_18_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_19_LC_18_17_4  (
            .in0(N__68277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83987),
            .ce(N__78361),
            .sr(N__77371));
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_18_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_18_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_18_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_14_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78951),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83987),
            .ce(N__78361),
            .sr(N__77371));
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_18_17_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_18_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_18_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_20_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68219),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83987),
            .ce(N__78361),
            .sr(N__77371));
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_18_17_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_18_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_18_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_15_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68697),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83987),
            .ce(N__78361),
            .sr(N__77371));
    defparam \dron_frame_decoder_1.source_H_disp_side_13_LC_18_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_13_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_13_LC_18_18_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_13_LC_18_18_0  (
            .in0(N__68909),
            .in1(N__71957),
            .in2(N__68654),
            .in3(N__71753),
            .lcout(drone_H_disp_side_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84005),
            .ce(),
            .sr(N__77378));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNING9E_13_LC_18_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNING9E_13_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNING9E_13_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNING9E_13_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68908),
            .lcout(drone_H_disp_side_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_5_LC_18_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_5_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_5_LC_18_18_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_5_LC_18_18_2  (
            .in0(N__68592),
            .in1(N__71959),
            .in2(N__68655),
            .in3(N__71755),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84005),
            .ce(),
            .sr(N__77378));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI8PL8_5_LC_18_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI8PL8_5_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI8PL8_5_LC_18_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNI8PL8_5_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68591),
            .lcout(drone_H_disp_side_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_2_LC_18_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_2_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_2_LC_18_18_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_2_LC_18_18_4  (
            .in0(N__68583),
            .in1(N__71958),
            .in2(N__71844),
            .in3(N__71754),
            .lcout(drone_H_disp_side_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84005),
            .ce(),
            .sr(N__77378));
    defparam \pid_side.error_axb_2_LC_18_18_5 .C_ON=1'b0;
    defparam \pid_side.error_axb_2_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_2_LC_18_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_2_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68582),
            .lcout(\pid_side.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_6_LC_18_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_6_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_6_LC_18_18_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_6_LC_18_18_6  (
            .in0(N__68490),
            .in1(N__71960),
            .in2(N__68564),
            .in3(N__71756),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84005),
            .ce(),
            .sr(N__77378));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI9QL8_6_LC_18_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI9QL8_6_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNI9QL8_6_LC_18_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNI9QL8_6_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68489),
            .lcout(drone_H_disp_side_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_inv_LC_18_19_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_inv_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_inv_LC_18_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_cry_0_c_inv_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__68838),
            .in3(N__72000),
            .lcout(\pid_side.error_axb_0 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\pid_side.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIRKB9_LC_18_19_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_RNIRKB9_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIRKB9_LC_18_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_cry_0_c_RNIRKB9_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__68829),
            .in3(N__68808),
            .lcout(\pid_side.error_1 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0 ),
            .carryout(\pid_side.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNITNC9_LC_18_19_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_c_RNITNC9_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNITNC9_LC_18_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_1_c_RNITNC9_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__68805),
            .in2(_gnd_net_),
            .in3(N__68799),
            .lcout(\pid_side.error_2 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1 ),
            .carryout(\pid_side.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIVQD9_LC_18_19_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_c_RNIVQD9_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIVQD9_LC_18_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_2_c_RNIVQD9_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__68796),
            .in2(_gnd_net_),
            .in3(N__68775),
            .lcout(\pid_side.error_3 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2 ),
            .carryout(\pid_side.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIODAN_LC_18_19_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_c_RNIODAN_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIODAN_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_c_RNIODAN_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__68772),
            .in2(N__68766),
            .in3(N__68754),
            .lcout(\pid_side.error_4 ),
            .ltout(),
            .carryin(\pid_side.error_cry_3 ),
            .carryout(\pid_side.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNI6LA11_LC_18_19_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_0_c_RNI6LA11_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNI6LA11_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_0_0_c_RNI6LA11_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__68751),
            .in2(N__68745),
            .in3(N__68736),
            .lcout(\pid_side.error_5 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0_0 ),
            .carryout(\pid_side.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNI9RG51_LC_18_19_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_0_c_RNI9RG51_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNI9RG51_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNI9RG51_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__68733),
            .in2(N__68727),
            .in3(N__68718),
            .lcout(\pid_side.error_6 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1_0 ),
            .carryout(\pid_side.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIC1NP_LC_18_19_7 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_0_c_RNIC1NP_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIC1NP_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIC1NP_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__68715),
            .in2(N__68709),
            .in3(N__68700),
            .lcout(\pid_side.error_7 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2_0 ),
            .carryout(\pid_side.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIF7TT_LC_18_20_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_0_c_RNIF7TT_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIF7TT_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIF7TT_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__72081),
            .in2(N__69078),
            .in3(N__69066),
            .lcout(\pid_side.error_8 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\pid_side.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI3QBN_LC_18_20_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_4_c_RNI3QBN_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI3QBN_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_4_c_RNI3QBN_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__69063),
            .in2(N__69054),
            .in3(N__68979),
            .lcout(\pid_side.error_9 ),
            .ltout(),
            .carryin(\pid_side.error_cry_4 ),
            .carryout(\pid_side.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIDD0T_LC_18_20_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_5_c_RNIDD0T_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIDD0T_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_5_c_RNIDD0T_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__71685),
            .in2(N__68976),
            .in3(N__68964),
            .lcout(\pid_side.error_10 ),
            .ltout(),
            .carryin(\pid_side.error_cry_5 ),
            .carryout(\pid_side.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIHK4U_LC_18_20_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_6_c_RNIHK4U_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIHK4U_LC_18_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_6_c_RNIHK4U_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__68961),
            .in2(_gnd_net_),
            .in3(N__68955),
            .lcout(\pid_side.error_11 ),
            .ltout(),
            .carryin(\pid_side.error_cry_6 ),
            .carryout(\pid_side.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIULOQ1_LC_18_20_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_7_c_RNIULOQ1_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIULOQ1_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_7_c_RNIULOQ1_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__68952),
            .in2(N__68946),
            .in3(N__68925),
            .lcout(\pid_side.error_12 ),
            .ltout(),
            .carryin(\pid_side.error_cry_7 ),
            .carryout(\pid_side.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNICGHT_LC_18_20_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_8_c_RNICGHT_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNICGHT_LC_18_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_8_c_RNICGHT_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__68922),
            .in2(N__68916),
            .in3(N__68895),
            .lcout(\pid_side.error_13 ),
            .ltout(),
            .carryin(\pid_side.error_cry_8 ),
            .carryout(\pid_side.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNIFKIT_LC_18_20_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_9_c_RNIFKIT_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIFKIT_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_9_c_RNIFKIT_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__68892),
            .in2(N__68865),
            .in3(N__68883),
            .lcout(\pid_side.error_14 ),
            .ltout(),
            .carryin(\pid_side.error_cry_9 ),
            .carryout(\pid_side.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNIPTP21_LC_18_20_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIPTP21_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIPTP21_LC_18_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_cry_10_c_RNIPTP21_LC_18_20_7  (
            .in0(N__68876),
            .in1(N__68864),
            .in2(_gnd_net_),
            .in3(N__68841),
            .lcout(\pid_side.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIJF6H2_LC_18_21_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNIJF6H2_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIJF6H2_LC_18_21_0 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_side.error_cry_6_c_RNIJF6H2_LC_18_21_0  (
            .in0(N__71542),
            .in1(N__71198),
            .in2(N__73304),
            .in3(N__71304),
            .lcout(\pid_side.m87_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_18_21_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_18_21_1 .LUT_INIT=16'b0010011101010101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_7_21_LC_18_21_1  (
            .in0(N__71146),
            .in1(N__71308),
            .in2(N__71216),
            .in3(N__72275),
            .lcout(),
            .ltout(\pid_side.m87_0_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_18_21_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_18_21_2 .LUT_INIT=16'b1100000111110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_21_LC_18_21_2  (
            .in0(N__70962),
            .in1(N__73504),
            .in2(N__71253),
            .in3(N__70893),
            .lcout(\pid_side.N_88_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNINI513_LC_18_21_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_6_c_RNINI513_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNINI513_LC_18_21_3 .LUT_INIT=16'b0100001101001111;
    LogicCell40 \pid_side.error_cry_6_c_RNINI513_LC_18_21_3  (
            .in0(N__71199),
            .in1(N__72274),
            .in2(N__71161),
            .in3(N__70961),
            .lcout(),
            .ltout(\pid_side.m36_1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNINJD15_LC_18_21_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNINJD15_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNINJD15_LC_18_21_4 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_cry_8_c_RNINJD15_LC_18_21_4  (
            .in0(N__73503),
            .in1(N__70892),
            .in2(N__70842),
            .in3(N__70809),
            .lcout(\pid_side.N_37_1 ),
            .ltout(\pid_side.N_37_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_18_21_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_18_21_5 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_22_LC_18_21_5  (
            .in0(N__70697),
            .in1(N__70509),
            .in2(N__70110),
            .in3(N__70040),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_22_LC_18_21_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_22_LC_18_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_22_LC_18_21_6 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \pid_side.error_i_reg_esr_22_LC_18_21_6  (
            .in0(N__69873),
            .in1(N__69626),
            .in2(N__69357),
            .in3(N__69354),
            .lcout(\pid_side.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84052),
            .ce(N__69324),
            .sr(N__77393));
    defparam \dron_frame_decoder_1.source_H_disp_side_0_LC_18_22_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_0_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_0_LC_18_22_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_0_LC_18_22_1  (
            .in0(N__71978),
            .in1(N__72054),
            .in2(N__71765),
            .in3(N__69133),
            .lcout(drone_H_disp_side_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84071),
            .ce(),
            .sr(N__77398));
    defparam \dron_frame_decoder_1.source_H_disp_side_8_LC_18_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_8_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_8_LC_18_22_3 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_8_LC_18_22_3  (
            .in0(N__71761),
            .in1(N__72055),
            .in2(N__71985),
            .in3(N__72093),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84071),
            .ce(),
            .sr(N__77398));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIBSL8_8_LC_18_22_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIBSL8_8_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIBSL8_8_LC_18_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNIBSL8_8_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72092),
            .lcout(drone_H_disp_side_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_0_LC_18_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_0_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_0_LC_18_22_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_fast_0_LC_18_22_5  (
            .in0(N__71983),
            .in1(N__72056),
            .in2(N__71766),
            .in3(N__71999),
            .lcout(dron_frame_decoder_1_source_H_disp_side_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84071),
            .ce(),
            .sr(N__77398));
    defparam \dron_frame_decoder_1.source_H_disp_side_10_LC_18_22_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_10_LC_18_22_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_10_LC_18_22_6 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_10_LC_18_22_6  (
            .in0(N__71694),
            .in1(N__71979),
            .in2(N__71843),
            .in3(N__71760),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84071),
            .ce(),
            .sr(N__77398));
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIKD9E_10_LC_18_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIKD9E_10_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_RNIKD9E_10_LC_18_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_RNIKD9E_10_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71693),
            .lcout(drone_H_disp_side_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_11_20_LC_18_23_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_11_20_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_11_20_LC_18_23_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_11_20_LC_18_23_0  (
            .in0(N__73227),
            .in1(N__71659),
            .in2(N__72707),
            .in3(N__73154),
            .lcout(\pid_side.m30_1_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_23_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_23_3 .LUT_INIT=16'b1010000110101011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_8_21_LC_18_23_3  (
            .in0(N__73080),
            .in1(N__72788),
            .in2(N__72999),
            .in3(N__72573),
            .lcout(\pid_side.N_12_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80510),
            .lcout(xy_ki_0_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84083),
            .ce(N__73411),
            .sr(N__77401));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_23_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_23_5  (
            .in0(N__80509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84083),
            .ce(N__73411),
            .sr(N__77401));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_23_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_23_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73769),
            .lcout(xy_ki_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84083),
            .ce(N__73411),
            .sr(N__77401));
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_18_23_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_18_23_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_18_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_1_LC_18_23_7  (
            .in0(N__73770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84083),
            .ce(N__73411),
            .sr(N__77401));
    defparam \pid_side.error_i_reg_esr_RNO_12_20_LC_18_24_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_12_20_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_12_20_LC_18_24_3 .LUT_INIT=16'b0100001101001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_12_20_LC_18_24_3  (
            .in0(N__72569),
            .in1(N__72989),
            .in2(N__72699),
            .in3(N__72504),
            .lcout(),
            .ltout(\pid_side.g0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_10_20_LC_18_24_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_10_20_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_10_20_LC_18_24_4 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_10_20_LC_18_24_4  (
            .in0(N__72990),
            .in1(N__72345),
            .in2(N__73317),
            .in3(N__72426),
            .lcout(\pid_side.N_28_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_18_24_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_18_24_5 .LUT_INIT=16'b0000011110100111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_11_21_LC_18_24_5  (
            .in0(N__73228),
            .in1(N__73051),
            .in2(N__72698),
            .in3(N__73158),
            .lcout(\pid_side.m11_0_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_9_20_LC_18_24_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_9_20_LC_18_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_9_20_LC_18_24_6 .LUT_INIT=16'b1100000111110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_9_20_LC_18_24_6  (
            .in0(N__73052),
            .in1(N__72991),
            .in2(N__72810),
            .in3(N__72789),
            .lcout(\pid_side.N_15_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNILTPJ2_LC_18_25_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNILTPJ2_LC_18_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNILTPJ2_LC_18_25_6 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_0_0_c_RNILTPJ2_LC_18_25_6  (
            .in0(N__72703),
            .in1(N__72583),
            .in2(N__72273),
            .in3(N__72505),
            .lcout(),
            .ltout(\pid_side.g0_i_m4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNIKJIE4_LC_18_25_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_0_c_RNIKJIE4_LC_18_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNIKJIE4_LC_18_25_7 .LUT_INIT=16'b1111000001010011;
    LogicCell40 \pid_side.error_cry_2_0_c_RNIKJIE4_LC_18_25_7  (
            .in0(N__72410),
            .in1(N__72346),
            .in2(N__72279),
            .in3(N__72260),
            .lcout(\pid_side.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_20_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_20_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_20_7_1  (
            .in0(_gnd_net_),
            .in1(N__76475),
            .in2(_gnd_net_),
            .in3(N__76155),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_20_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_20_7_2 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILVE13_0_LC_20_7_2  (
            .in0(N__76480),
            .in1(N__73923),
            .in2(N__73938),
            .in3(N__74178),
            .lcout(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_20_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_20_7_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_20_7_3  (
            .in0(N__74303),
            .in1(N__76477),
            .in2(_gnd_net_),
            .in3(N__76157),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_20_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_20_7_4 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_20_7_4  (
            .in0(N__76479),
            .in1(N__77906),
            .in2(N__73933),
            .in3(N__74177),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_20_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_20_7_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_20_7_5  (
            .in0(N__73870),
            .in1(N__76476),
            .in2(_gnd_net_),
            .in3(N__76156),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_20_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_20_7_7 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_20_7_7  (
            .in0(N__77905),
            .in1(N__76478),
            .in2(N__77948),
            .in3(N__76158),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_20_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_20_8_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_20_8_0  (
            .in0(N__77904),
            .in1(N__76612),
            .in2(N__76292),
            .in3(N__73822),
            .lcout(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_20_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_20_8_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_20_8_2  (
            .in0(N__73976),
            .in1(N__76277),
            .in2(_gnd_net_),
            .in3(N__76611),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_20_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_20_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_20_8_3  (
            .in0(N__76610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74150),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_20_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_20_8_4 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_20_8_4  (
            .in0(N__77903),
            .in1(N__74225),
            .in2(N__74168),
            .in3(N__76613),
            .lcout(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_20_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_20_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_20_8_5  (
            .in0(N__76615),
            .in1(N__77902),
            .in2(N__74175),
            .in3(N__74199),
            .lcout(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_20_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_20_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_20_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_20_8_7  (
            .in0(N__76614),
            .in1(N__77901),
            .in2(N__74174),
            .in3(N__74108),
            .lcout(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_20_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_20_9_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_20_9_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_20_9_0  (
            .in0(N__74419),
            .in1(N__77739),
            .in2(N__74568),
            .in3(N__74079),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83908),
            .ce(),
            .sr(N__77339));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_20_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_20_9_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_20_9_1  (
            .in0(N__74044),
            .in1(N__76616),
            .in2(_gnd_net_),
            .in3(N__76272),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_20_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_20_9_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_20_9_2  (
            .in0(N__76617),
            .in1(_gnd_net_),
            .in2(N__76291),
            .in3(N__74045),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_20_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_20_9_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_20_9_3  (
            .in0(N__74046),
            .in1(N__74903),
            .in2(N__74789),
            .in3(N__74034),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_20_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_20_9_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_20_9_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_20_9_4  (
            .in0(N__74420),
            .in1(N__77724),
            .in2(N__74569),
            .in3(N__73995),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83908),
            .ce(),
            .sr(N__77339));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_20_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_20_9_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_20_9_5  (
            .in0(N__73975),
            .in1(N__76618),
            .in2(_gnd_net_),
            .in3(N__76276),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_20_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_20_10_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_20_10_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_20_10_0  (
            .in0(N__74422),
            .in1(N__78036),
            .in2(N__74570),
            .in3(N__74946),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83919),
            .ce(),
            .sr(N__77344));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_20_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_20_10_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_20_10_1  (
            .in0(N__76619),
            .in1(N__74803),
            .in2(_gnd_net_),
            .in3(N__76278),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_20_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_20_10_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_20_10_2  (
            .in0(N__76279),
            .in1(_gnd_net_),
            .in2(N__74808),
            .in3(N__76620),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_20_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_20_10_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_20_10_3  (
            .in0(N__74904),
            .in1(N__74807),
            .in2(N__74793),
            .in3(N__74652),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_20_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_20_10_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_20_10_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_20_10_4  (
            .in0(N__74613),
            .in1(N__74560),
            .in2(N__74427),
            .in3(N__77979),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83919),
            .ce(),
            .sr(N__77344));
    defparam \ppm_encoder_1.init_pulses_17_LC_20_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_20_10_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_20_10_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_20_10_5  (
            .in0(N__74561),
            .in1(N__74426),
            .in2(N__77961),
            .in3(N__74316),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83919),
            .ce(),
            .sr(N__77344));
    defparam \pid_side.error_p_reg_esr_3_LC_20_11_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_3_LC_20_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_3_LC_20_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_3_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74277),
            .lcout(\pid_side.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83932),
            .ce(N__82451),
            .sr(N__82866));
    defparam \pid_side.error_p_reg_esr_2_LC_20_12_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_2_LC_20_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_2_LC_20_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_2_LC_20_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74244),
            .lcout(\pid_side.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83944),
            .ce(N__82414),
            .sr(N__82862));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_13_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_13_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_13_0  (
            .in0(N__79094),
            .in1(N__79106),
            .in2(_gnd_net_),
            .in3(N__79526),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_13_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_13_1 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_13_1  (
            .in0(N__78311),
            .in1(N__81362),
            .in2(N__75108),
            .in3(N__78290),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_13_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_13_2  (
            .in0(N__75005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75017),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_13_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_13_3 .LUT_INIT=16'b0110100100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_13_3  (
            .in0(N__78313),
            .in1(N__74955),
            .in2(N__81774),
            .in3(N__78288),
            .lcout(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_13_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_13_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__75084),
            .in3(N__75081),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_13_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_13_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_13_5  (
            .in0(N__75018),
            .in1(N__75047),
            .in2(N__75036),
            .in3(N__75006),
            .lcout(\pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_13_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_13_6  (
            .in0(N__78289),
            .in1(N__78312),
            .in2(N__81363),
            .in3(N__75024),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ),
            .ltout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_13_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_13_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__75009),
            .in3(N__75004),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_20_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_20_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_20_14_0  (
            .in0(_gnd_net_),
            .in1(N__75202),
            .in2(_gnd_net_),
            .in3(N__78414),
            .lcout(\pid_side.N_1869_i ),
            .ltout(\pid_side.N_1869_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_20_14_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_20_14_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_20_14_1  (
            .in0(N__78314),
            .in1(N__78291),
            .in2(N__74949),
            .in3(N__81773),
            .lcout(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_20_14_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_20_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_20_14_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIODMH3_6_LC_20_14_2  (
            .in0(_gnd_net_),
            .in1(N__75264),
            .in2(N__75267),
            .in3(N__75249),
            .lcout(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_20_14_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_20_14_3 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_20_14_3  (
            .in0(N__78415),
            .in1(N__81335),
            .in2(N__75207),
            .in3(N__78401),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_20_14_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_20_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_20_14_4  (
            .in0(_gnd_net_),
            .in1(N__75258),
            .in2(N__75252),
            .in3(N__75248),
            .lcout(\pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_6_LC_20_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_20_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_6_LC_20_14_5  (
            .in0(N__78417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83973),
            .ce(N__81190),
            .sr(N__81145));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_20_14_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_20_14_6 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_7_LC_20_14_6  (
            .in0(N__78402),
            .in1(N__75206),
            .in2(N__81339),
            .in3(N__78416),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIT9E37_7_LC_20_14_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIT9E37_7_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIT9E37_7_LC_20_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIT9E37_7_LC_20_14_7  (
            .in0(N__75176),
            .in1(N__75926),
            .in2(N__75162),
            .in3(N__75158),
            .lcout(\pid_side.error_p_reg_esr_RNIT9E37Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_15_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_15_0 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_15_0  (
            .in0(N__75448),
            .in1(N__78507),
            .in2(N__81810),
            .in3(N__78585),
            .lcout(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_9_LC_20_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_20_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_20_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_9_LC_20_15_1  (
            .in0(N__78588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83989),
            .ce(N__81199),
            .sr(N__81144));
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_15_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_15_2 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_15_2  (
            .in0(N__75447),
            .in1(N__78506),
            .in2(N__81809),
            .in3(N__78584),
            .lcout(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_20_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_20_15_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_20_15_3  (
            .in0(N__78586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75449),
            .lcout(\pid_side.N_1887_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_10_LC_20_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_20_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_20_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_10_LC_20_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78509),
            .lcout(\pid_side.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83989),
            .ce(N__81199),
            .sr(N__81144));
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_20_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_20_15_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_20_15_5  (
            .in0(N__78508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75468),
            .lcout(),
            .ltout(\pid_side.N_1893_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_20_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_20_15_6 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_20_15_6  (
            .in0(N__75450),
            .in1(N__81808),
            .in2(N__75435),
            .in3(N__78587),
            .lcout(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ),
            .ltout(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_20_15_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_20_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIBMBO6_10_LC_20_15_7  (
            .in0(N__75893),
            .in1(N__75512),
            .in2(N__75417),
            .in3(N__75414),
            .lcout(\pid_side.error_p_reg_esr_RNIBMBO6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_20_16_0  (
            .in0(N__75273),
            .in1(N__75318),
            .in2(N__75372),
            .in3(N__75590),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_20_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_20_16_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_20_16_1  (
            .in0(N__81889),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75618),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_16_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_16_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_20_16_2  (
            .in0(N__78647),
            .in1(N__75308),
            .in2(_gnd_net_),
            .in3(N__75291),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ),
            .ltout(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_16_3 .LUT_INIT=16'b1110100011111010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_20_16_3  (
            .in0(N__75591),
            .in1(N__81900),
            .in2(N__75663),
            .in3(N__75620),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_16_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_16_4 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_1_LC_20_16_4  (
            .in0(N__75634),
            .in1(N__81887),
            .in2(N__78550),
            .in3(N__81927),
            .lcout(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_20_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_0_LC_20_16_5  (
            .in0(N__81929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84007),
            .ce(N__81248),
            .sr(N__81142));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_16_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_16_6 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_20_16_6  (
            .in0(N__75635),
            .in1(N__81888),
            .in2(N__78551),
            .in3(N__81928),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_16_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_20_16_7  (
            .in0(_gnd_net_),
            .in1(N__75619),
            .in2(N__75600),
            .in3(N__75597),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_20_17_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_20_17_0 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_8_LC_20_17_0  (
            .in0(N__78621),
            .in1(N__80670),
            .in2(N__78393),
            .in3(N__75939),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ),
            .ltout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_20_17_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_20_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIECBV6_8_LC_20_17_1  (
            .in0(N__75582),
            .in1(N__75491),
            .in2(N__75561),
            .in3(N__75545),
            .lcout(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_20_17_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_20_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI9GJD3_8_LC_20_17_2  (
            .in0(N__75546),
            .in1(_gnd_net_),
            .in2(N__75495),
            .in3(N__75522),
            .lcout(\pid_side.error_p_reg_esr_RNI9GJD3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_20_17_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_20_17_3 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_20_17_3  (
            .in0(N__78880),
            .in1(N__81434),
            .in2(N__78863),
            .in3(N__75911),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_20_17_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_20_17_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(N__78856),
            .in2(_gnd_net_),
            .in3(N__78879),
            .lcout(\pid_side.N_1881_i ),
            .ltout(\pid_side.N_1881_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_20_17_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_20_17_5 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_20_17_5  (
            .in0(N__80669),
            .in1(N__78389),
            .in2(N__75933),
            .in3(N__78620),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_20_17_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_20_17_7 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_20_17_7  (
            .in0(N__78881),
            .in1(N__81435),
            .in2(N__78864),
            .in3(N__75912),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_4_LC_20_18_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_4_LC_20_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_4_LC_20_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_4_LC_20_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75876),
            .lcout(\pid_front.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84039),
            .ce(N__83182),
            .sr(N__82854));
    defparam \pid_front.error_d_reg_esr_2_LC_20_18_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_2_LC_20_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_2_LC_20_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_2_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75843),
            .lcout(\pid_front.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84039),
            .ce(N__83182),
            .sr(N__82854));
    defparam \pid_front.error_d_reg_esr_9_LC_20_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_9_LC_20_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_9_LC_20_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_9_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75807),
            .lcout(\pid_front.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84054),
            .ce(N__83156),
            .sr(N__82852));
    defparam \pid_front.error_d_reg_esr_11_LC_20_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_11_LC_20_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_11_LC_20_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_11_LC_20_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75747),
            .lcout(\pid_front.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84073),
            .ce(N__83183),
            .sr(N__82850));
    defparam \pid_front.error_d_reg_esr_3_LC_20_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_3_LC_20_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_3_LC_20_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_3_LC_20_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75702),
            .lcout(\pid_front.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84092),
            .ce(N__83184),
            .sr(N__82849));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_29_7.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_29_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_29_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_29_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77587),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_21_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_21_7_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_21_7_0  (
            .in0(N__76698),
            .in1(N__76166),
            .in2(_gnd_net_),
            .in3(N__76488),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_21_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_21_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_21_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_21_7_1  (
            .in0(N__76490),
            .in1(N__76670),
            .in2(_gnd_net_),
            .in3(N__76175),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_21_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_21_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_21_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_21_7_5  (
            .in0(N__76489),
            .in1(N__76319),
            .in2(_gnd_net_),
            .in3(N__76174),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_21_8_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_21_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_21_8_0  (
            .in0(_gnd_net_),
            .in1(N__76044),
            .in2(N__76032),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_8_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_21_8_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_21_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_21_8_1  (
            .in0(_gnd_net_),
            .in1(N__76023),
            .in2(_gnd_net_),
            .in3(N__76002),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_21_8_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_21_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_21_8_2  (
            .in0(_gnd_net_),
            .in1(N__75999),
            .in2(N__75993),
            .in3(N__75972),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_21_8_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_21_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_21_8_3  (
            .in0(_gnd_net_),
            .in1(N__75969),
            .in2(_gnd_net_),
            .in3(N__75951),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_21_8_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_21_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_21_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_21_8_4  (
            .in0(_gnd_net_),
            .in1(N__75948),
            .in2(_gnd_net_),
            .in3(N__77838),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_21_8_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_21_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_21_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_21_8_5  (
            .in0(_gnd_net_),
            .in1(N__77835),
            .in2(_gnd_net_),
            .in3(N__77811),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_21_8_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_21_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_21_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_21_8_6  (
            .in0(_gnd_net_),
            .in1(N__77808),
            .in2(N__77793),
            .in3(N__77772),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_21_8_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_21_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_21_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_21_8_7  (
            .in0(_gnd_net_),
            .in1(N__77769),
            .in2(_gnd_net_),
            .in3(N__77748),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_21_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_21_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_21_9_0  (
            .in0(_gnd_net_),
            .in1(N__77745),
            .in2(_gnd_net_),
            .in3(N__77733),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_21_9_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_21_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_21_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_21_9_1  (
            .in0(_gnd_net_),
            .in1(N__77730),
            .in2(_gnd_net_),
            .in3(N__77718),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_21_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_21_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_21_9_2  (
            .in0(_gnd_net_),
            .in1(N__77715),
            .in2(_gnd_net_),
            .in3(N__77691),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_21_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_21_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_21_9_3  (
            .in0(_gnd_net_),
            .in1(N__77688),
            .in2(_gnd_net_),
            .in3(N__77670),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_21_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_21_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_21_9_4  (
            .in0(_gnd_net_),
            .in1(N__78105),
            .in2(_gnd_net_),
            .in3(N__78087),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_21_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_21_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(N__78084),
            .in2(N__78063),
            .in3(N__78045),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_21_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_21_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_21_9_6  (
            .in0(_gnd_net_),
            .in1(N__78042),
            .in2(_gnd_net_),
            .in3(N__78030),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_21_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_21_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_21_9_7  (
            .in0(_gnd_net_),
            .in1(N__78027),
            .in2(_gnd_net_),
            .in3(N__77997),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_21_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_21_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_21_10_0  (
            .in0(_gnd_net_),
            .in1(N__77994),
            .in2(_gnd_net_),
            .in3(N__77973),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_21_10_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_21_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_21_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(N__77970),
            .in2(_gnd_net_),
            .in3(N__77952),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_21_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_21_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_21_10_2  (
            .in0(N__77941),
            .in1(N__77913),
            .in2(_gnd_net_),
            .in3(N__77877),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_4_LC_21_12_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_4_LC_21_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_4_LC_21_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_4_LC_21_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77865),
            .lcout(\pid_side.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83959),
            .ce(N__82415),
            .sr(N__82867));
    defparam \pid_side.error_d_reg_esr_5_LC_21_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_5_LC_21_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_5_LC_21_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_5_LC_21_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78441),
            .lcout(\pid_side.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83974),
            .ce(N__82431),
            .sr(N__82863));
    defparam \pid_side.error_d_reg_esr_6_LC_21_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_6_LC_21_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_6_LC_21_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_6_LC_21_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78429),
            .lcout(\pid_side.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83974),
            .ce(N__82431),
            .sr(N__82863));
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_21_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_21_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_21_14_0  (
            .in0(_gnd_net_),
            .in1(N__78380),
            .in2(_gnd_net_),
            .in3(N__78613),
            .lcout(\pid_side.N_1875_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_7_LC_21_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_21_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_21_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_7_LC_21_14_1  (
            .in0(N__78614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83990),
            .ce(N__81189),
            .sr(N__81146));
    defparam \pid_side.state_RNI7OA81_0_LC_21_14_2 .C_ON=1'b0;
    defparam \pid_side.state_RNI7OA81_0_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI7OA81_0_LC_21_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNI7OA81_0_LC_21_14_2  (
            .in0(_gnd_net_),
            .in1(N__78369),
            .in2(_gnd_net_),
            .in3(N__81153),
            .lcout(\pid_side.N_478_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_4_LC_21_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_21_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_21_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_4_LC_21_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79530),
            .lcout(\pid_side.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83990),
            .ce(N__81189),
            .sr(N__81146));
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_21_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_13_LC_21_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82583),
            .lcout(\pid_side.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83990),
            .ce(N__81189),
            .sr(N__81146));
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_21_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_5_LC_21_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78315),
            .lcout(\pid_side.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83990),
            .ce(N__81189),
            .sr(N__81146));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_21_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_21_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_21_14_7  (
            .in0(_gnd_net_),
            .in1(N__78273),
            .in2(_gnd_net_),
            .in3(N__78243),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_2_LC_21_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_2_LC_21_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_2_LC_21_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_2_LC_21_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78666),
            .lcout(\pid_side.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84008),
            .ce(N__82432),
            .sr(N__82860));
    defparam \pid_side.error_d_reg_esr_7_LC_21_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_7_LC_21_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_7_LC_21_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_7_LC_21_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78636),
            .lcout(\pid_side.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84008),
            .ce(N__82432),
            .sr(N__82860));
    defparam \pid_side.error_d_reg_esr_9_LC_21_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_9_LC_21_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_9_LC_21_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_9_LC_21_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78600),
            .lcout(\pid_side.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84008),
            .ce(N__82432),
            .sr(N__82860));
    defparam \pid_side.error_p_reg_esr_1_LC_21_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_1_LC_21_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_1_LC_21_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_1_LC_21_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78570),
            .lcout(\pid_side.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84008),
            .ce(N__82432),
            .sr(N__82860));
    defparam \pid_side.error_d_reg_esr_10_LC_21_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_10_LC_21_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_10_LC_21_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_10_LC_21_15_7  (
            .in0(N__78528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84008),
            .ce(N__82432),
            .sr(N__82860));
    defparam \pid_side.error_p_reg_esr_RNIQOFJ2_12_LC_21_16_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIQOFJ2_12_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIQOFJ2_12_LC_21_16_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIQOFJ2_12_LC_21_16_0  (
            .in0(N__81321),
            .in1(N__82069),
            .in2(_gnd_net_),
            .in3(N__80526),
            .lcout(\pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12 ),
            .ltout(\pid_side.error_p_reg_esr_RNIQOFJ2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIVTS3_12_LC_21_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIVTS3_12_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIVTS3_12_LC_21_16_1 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIVTS3_12_LC_21_16_1  (
            .in0(N__82633),
            .in1(N__81308),
            .in2(N__78468),
            .in3(N__79411),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIIVTS3Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_0_12_LC_21_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_0_12_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_0_12_LC_21_16_2 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ7S9A_0_12_LC_21_16_2  (
            .in0(N__78973),
            .in1(N__78949),
            .in2(N__78465),
            .in3(N__78984),
            .lcout(\pid_side.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_16_4 .LUT_INIT=16'b0011100110011100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7J5H1_13_LC_21_16_4  (
            .in0(N__79371),
            .in1(N__79316),
            .in2(N__82582),
            .in3(N__80738),
            .lcout(),
            .ltout(\pid_side.error_d_reg_prev_esr_RNI7J5H1Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_5 .LUT_INIT=16'b0010110110110100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_5  (
            .in0(N__79302),
            .in1(N__79410),
            .in2(N__78987),
            .in3(N__79296),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_12_LC_21_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_12_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ7S9A_12_LC_21_16_6 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ7S9A_12_LC_21_16_6  (
            .in0(N__78974),
            .in1(N__78950),
            .in2(N__78927),
            .in3(N__78924),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQ7S9AZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_21_16_7  (
            .in0(N__80737),
            .in1(N__79370),
            .in2(_gnd_net_),
            .in3(N__82572),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2OIO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_8_LC_21_17_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_8_LC_21_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_8_LC_21_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_8_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78894),
            .lcout(\pid_side.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84040),
            .ce(N__82456),
            .sr(N__82859));
    defparam \pid_side.error_d_reg_prev_esr_8_LC_21_18_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_21_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_21_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_8_LC_21_18_3  (
            .in0(N__78882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84055),
            .ce(N__81249),
            .sr(N__81141));
    defparam \pid_front.error_d_reg_esr_10_LC_21_19_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_10_LC_21_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_10_LC_21_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_10_LC_21_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78846),
            .lcout(\pid_front.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84074),
            .ce(N__83188),
            .sr(N__82855));
    defparam \pid_front.error_d_reg_esr_12_LC_21_19_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_12_LC_21_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_12_LC_21_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_12_LC_21_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78786),
            .lcout(\pid_front.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84074),
            .ce(N__83188),
            .sr(N__82855));
    defparam \pid_front.error_d_reg_esr_13_LC_21_19_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_13_LC_21_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_13_LC_21_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_13_LC_21_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78711),
            .lcout(\pid_front.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84074),
            .ce(N__83188),
            .sr(N__82855));
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_21_22_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_21_22_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_21_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_4_LC_21_22_4  (
            .in0(_gnd_net_),
            .in1(N__79290),
            .in2(_gnd_net_),
            .in3(N__83006),
            .lcout(xy_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84099),
            .ce(N__80918),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_22_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_22_13_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_22_13_0  (
            .in0(N__81408),
            .in1(N__79503),
            .in2(_gnd_net_),
            .in3(N__81705),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_13_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_22_13_3  (
            .in0(N__79107),
            .in1(N__79095),
            .in2(_gnd_net_),
            .in3(N__79522),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_14_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_22_14_0  (
            .in0(N__80696),
            .in1(N__79337),
            .in2(_gnd_net_),
            .in3(N__82541),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_14_LC_22_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_22_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_22_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_14_LC_22_14_1  (
            .in0(N__82542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84009),
            .ce(N__81191),
            .sr(N__81148));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_22_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_22_14_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_22_14_2  (
            .in0(N__81464),
            .in1(N__79022),
            .in2(_gnd_net_),
            .in3(N__81619),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_22_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_15_LC_22_14_3  (
            .in0(N__81621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84009),
            .ce(N__81191),
            .sr(N__81148));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_22_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_22_14_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_22_14_4  (
            .in0(N__81465),
            .in1(N__79023),
            .in2(_gnd_net_),
            .in3(N__81620),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_22_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_22_14_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_22_14_5  (
            .in0(N__81488),
            .in1(N__79478),
            .in2(_gnd_net_),
            .in3(N__81643),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_16_LC_22_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_22_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_22_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_16_LC_22_14_6  (
            .in0(N__81645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84009),
            .ce(N__81191),
            .sr(N__81148));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_22_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_22_14_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_22_14_7  (
            .in0(N__81489),
            .in1(N__79479),
            .in2(_gnd_net_),
            .in3(N__81644),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_22_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_22_15_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_22_15_0  (
            .in0(N__81407),
            .in1(N__79502),
            .in2(_gnd_net_),
            .in3(N__81704),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_1_12_LC_22_15_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_1_12_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_1_12_LC_22_15_4 .LUT_INIT=16'b0010001000101011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR3TQ1_1_12_LC_22_15_4  (
            .in0(N__80585),
            .in1(N__81851),
            .in2(N__82071),
            .in3(N__80545),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_167_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIJAB43_12_LC_22_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIJAB43_12_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIJAB43_12_LC_22_15_5 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIJAB43_12_LC_22_15_5  (
            .in0(N__79406),
            .in1(N__81296),
            .in2(N__79383),
            .in3(N__82640),
            .lcout(\pid_side.un1_pid_prereg_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_22_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_22_15_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_22_15_6  (
            .in0(N__80739),
            .in1(N__79369),
            .in2(_gnd_net_),
            .in3(N__82584),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2OIOZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_22_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_22_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_22_16_1  (
            .in0(N__79338),
            .in1(N__80697),
            .in2(_gnd_net_),
            .in3(N__82535),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_22_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_22_16_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_22_16_2  (
            .in0(_gnd_net_),
            .in1(N__81295),
            .in2(_gnd_net_),
            .in3(N__82632),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMERG_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_22_17_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_22_17_6 .LUT_INIT=16'b1101110111010100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_22_17_6  (
            .in0(N__80586),
            .in1(N__81852),
            .in2(N__80550),
            .in3(N__82070),
            .lcout(\pid_side.error_p_reg_esr_RNIR3TQ1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_22_19_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_0_LC_22_19_0  (
            .in0(_gnd_net_),
            .in1(N__80516),
            .in2(_gnd_net_),
            .in3(N__83008),
            .lcout(xy_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84085),
            .ce(N__80913),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_22_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_22_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_22_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_2_LC_22_19_2  (
            .in0(_gnd_net_),
            .in1(N__80291),
            .in2(_gnd_net_),
            .in3(N__83009),
            .lcout(xy_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84085),
            .ce(N__80913),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_22_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_5_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__80109),
            .in2(_gnd_net_),
            .in3(N__83010),
            .lcout(xy_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84085),
            .ce(N__80913),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_22_19_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_22_19_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_22_19_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_7_LC_22_19_6  (
            .in0(_gnd_net_),
            .in1(N__79931),
            .in2(_gnd_net_),
            .in3(N__83011),
            .lcout(xy_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84085),
            .ce(N__80913),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_22_21_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_22_21_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_22_21_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_3_LC_22_21_3  (
            .in0(_gnd_net_),
            .in1(N__79724),
            .in2(_gnd_net_),
            .in3(N__83007),
            .lcout(xy_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84100),
            .ce(N__80914),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_3_LC_23_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_3_LC_23_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_3_LC_23_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_3_LC_23_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79575),
            .lcout(\pid_side.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84010),
            .ce(N__82460),
            .sr(N__82869));
    defparam \pid_side.error_d_reg_esr_4_LC_23_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_4_LC_23_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_4_LC_23_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_4_LC_23_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79542),
            .lcout(\pid_side.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84010),
            .ce(N__82460),
            .sr(N__82869));
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_17_LC_23_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81703),
            .lcout(\pid_side.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84024),
            .ce(N__81230),
            .sr(N__81149));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_14_3  (
            .in0(N__81383),
            .in1(N__80651),
            .in2(_gnd_net_),
            .in3(N__81664),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_18_LC_23_14_4  (
            .in0(N__81666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84024),
            .ce(N__81230),
            .sr(N__81149));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_14_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_14_5  (
            .in0(N__81384),
            .in1(N__80652),
            .in2(_gnd_net_),
            .in3(N__81665),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_23_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_23_14_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_23_14_6  (
            .in0(N__82190),
            .in1(N__82172),
            .in2(_gnd_net_),
            .in3(N__82126),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_19_LC_23_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_23_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_23_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_19_LC_23_14_7  (
            .in0(N__82127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84024),
            .ce(N__81230),
            .sr(N__81149));
    defparam \pid_side.error_d_reg_esr_11_LC_23_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_11_LC_23_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_11_LC_23_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_11_LC_23_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80598),
            .lcout(\pid_side.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84041),
            .ce(N__82464),
            .sr(N__82864));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_23_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_23_16_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_23_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__81304),
            .in3(N__82618),
            .lcout(\pid_side.N_1905_i ),
            .ltout(\pid_side.N_1905_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_0_12_LC_23_16_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_0_12_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_0_12_LC_23_16_2 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR3TQ1_0_12_LC_23_16_2  (
            .in0(N__81838),
            .in1(N__80546),
            .in2(N__80574),
            .in3(N__82059),
            .lcout(\pid_side.error_p_reg_esr_RNIR3TQ1_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_23_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_23_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_23_16_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_23_16_3  (
            .in0(_gnd_net_),
            .in1(N__82024),
            .in2(_gnd_net_),
            .in3(N__82084),
            .lcout(\pid_side.un1_pid_prereg_79 ),
            .ltout(\pid_side.un1_pid_prereg_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIVHA21_12_LC_23_16_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIVHA21_12_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIVHA21_12_LC_23_16_4 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIVHA21_12_LC_23_16_4  (
            .in0(N__81836),
            .in1(N__81288),
            .in2(N__80529),
            .in3(N__82619),
            .lcout(\pid_side.error_p_reg_esr_RNIVHA21Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIVKIO_12_LC_23_16_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIVKIO_12_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIVKIO_12_LC_23_16_5 .LUT_INIT=16'b1111111100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIVKIO_12_LC_23_16_5  (
            .in0(_gnd_net_),
            .in1(N__82617),
            .in2(N__81303),
            .in3(N__81837),
            .lcout(\pid_side.error_p_reg_esr_RNIVKIOZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_12_LC_23_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_23_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_23_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_12_LC_23_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82620),
            .lcout(\pid_side.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84056),
            .ce(N__81247),
            .sr(N__81147));
    defparam \pid_side.error_d_reg_prev_esr_11_LC_23_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_23_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_23_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_11_LC_23_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82101),
            .lcout(\pid_side.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84056),
            .ce(N__81247),
            .sr(N__81147));
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_23_19_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_23_19_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_23_19_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_6_LC_23_19_7  (
            .in0(_gnd_net_),
            .in1(N__81100),
            .in2(_gnd_net_),
            .in3(N__83012),
            .lcout(xy_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84093),
            .ce(N__80919),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_21_LC_24_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80844),
            .lcout(\pid_side.error_p_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_13_LC_24_10_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_13_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(N__80748),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_14_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80706),
            .lcout(\pid_side.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_8_LC_24_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_8_LC_24_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80676),
            .lcout(\pid_side.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_16_LC_24_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_16_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81498),
            .lcout(\pid_side.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_15_LC_24_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_15_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81474),
            .lcout(\pid_side.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_20_LC_24_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_20_LC_24_10_6  (
            .in0(N__81450),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_9_LC_24_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_9_LC_24_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_9_LC_24_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_9_LC_24_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81441),
            .lcout(\pid_side.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83975),
            .ce(N__82458),
            .sr(N__82879));
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_19_LC_24_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_19_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81420),
            .lcout(\pid_side.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_17_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81414),
            .lcout(\pid_side.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_18_LC_24_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_18_LC_24_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81390),
            .lcout(\pid_side.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_5_LC_24_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_5_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_5_LC_24_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_5_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81369),
            .lcout(\pid_side.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_7_LC_24_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_7_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81345),
            .lcout(\pid_side.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_10_LC_24_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_10_LC_24_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81816),
            .lcout(\pid_side.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__83991),
            .ce(N__82453),
            .sr(N__82876));
    defparam \pid_side.error_p_reg_esr_6_LC_24_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_6_LC_24_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_6_LC_24_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_6_LC_24_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81780),
            .lcout(\pid_side.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84011),
            .ce(N__82452),
            .sr(N__82873));
    defparam \pid_side.error_p_reg_esr_0_LC_24_13_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_0_LC_24_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_0_LC_24_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_0_LC_24_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81753),
            .lcout(\pid_side.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84025),
            .ce(N__82454),
            .sr(N__82871));
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_17_LC_24_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81717),
            .lcout(\pid_side.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84042),
            .ce(N__82459),
            .sr(N__82870));
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_18_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81675),
            .lcout(\pid_side.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84042),
            .ce(N__82459),
            .sr(N__82870));
    defparam \pid_side.error_d_reg_esr_16_LC_24_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_16_LC_24_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_16_LC_24_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_16_LC_24_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81654),
            .lcout(\pid_side.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84042),
            .ce(N__82459),
            .sr(N__82870));
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_15_LC_24_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_15_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81630),
            .lcout(\pid_side.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84042),
            .ce(N__82459),
            .sr(N__82870));
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_22_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81606),
            .lcout(\pid_side.error_d_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84042),
            .ce(N__82459),
            .sr(N__82870));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_24_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_24_15_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_24_15_0  (
            .in0(N__82191),
            .in1(N__82173),
            .in2(_gnd_net_),
            .in3(N__82128),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_19_LC_24_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_19_LC_24_15_2  (
            .in0(N__82137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84057),
            .ce(N__82455),
            .sr(N__82868));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_24_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_24_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_24_15_3  (
            .in0(N__82100),
            .in1(N__82026),
            .in2(_gnd_net_),
            .in3(N__82086),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHIO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_24_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_24_15_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_24_15_5  (
            .in0(N__82099),
            .in1(N__82025),
            .in2(_gnd_net_),
            .in3(N__82085),
            .lcout(\pid_side.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_11_LC_24_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_11_LC_24_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_11_LC_24_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_11_LC_24_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82038),
            .lcout(\pid_side.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84057),
            .ce(N__82455),
            .sr(N__82868));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_24_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_24_15_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_24_15_7  (
            .in0(N__82004),
            .in1(N__81987),
            .in2(_gnd_net_),
            .in3(N__82475),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_0_LC_24_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_0_LC_24_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_0_LC_24_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_0_LC_24_16_0  (
            .in0(N__81942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_1_LC_24_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_1_LC_24_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_1_LC_24_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_1_LC_24_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81906),
            .lcout(\pid_side.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_p_reg_esr_12_LC_24_16_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_12_LC_24_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_12_LC_24_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_12_LC_24_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81864),
            .lcout(\pid_side.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_12_LC_24_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_12_LC_24_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_12_LC_24_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_12_LC_24_16_3  (
            .in0(N__82650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_13_LC_24_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_13_LC_24_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_13_LC_24_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_esr_13_LC_24_16_4  (
            .in0(N__82590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_14_LC_24_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_14_LC_24_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_14_LC_24_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_14_LC_24_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82548),
            .lcout(\pid_side.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_21_LC_24_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_21_LC_24_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_21_LC_24_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_21_LC_24_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82521),
            .lcout(\pid_side.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_side.error_d_reg_esr_20_LC_24_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_20_LC_24_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_20_LC_24_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_20_LC_24_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82494),
            .lcout(\pid_side.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84075),
            .ce(N__82457),
            .sr(N__82865));
    defparam \pid_front.error_d_reg_esr_8_LC_24_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_8_LC_24_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_8_LC_24_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_8_LC_24_17_1  (
            .in0(N__82320),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84086),
            .ce(N__83202),
            .sr(N__82861));
    defparam \pid_front.error_d_reg_esr_17_LC_24_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_17_LC_24_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_17_LC_24_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_17_LC_24_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82272),
            .lcout(\pid_front.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84103),
            .ce(N__83203),
            .sr(N__82857));
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_18_LC_24_22_0  (
            .in0(N__82239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84106),
            .ce(N__83201),
            .sr(N__82856));
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_19_LC_24_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84444),
            .lcout(\pid_front.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84106),
            .ce(N__83201),
            .sr(N__82856));
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_20_LC_24_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_20_LC_24_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84411),
            .lcout(\pid_front.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84106),
            .ce(N__83201),
            .sr(N__82856));
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_21_LC_24_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84363),
            .lcout(\pid_front.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84106),
            .ce(N__83201),
            .sr(N__82856));
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_22_LC_24_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84315),
            .lcout(\pid_front.error_d_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84106),
            .ce(N__83201),
            .sr(N__82856));
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_16_LC_24_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_16_LC_24_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84204),
            .lcout(\pid_front.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84110),
            .ce(N__83204),
            .sr(N__82853));
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_15_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84171),
            .lcout(\pid_front.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84110),
            .ce(N__83204),
            .sr(N__82853));
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_14_LC_24_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_14_LC_24_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84141),
            .lcout(\pid_front.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__84113),
            .ce(N__83208),
            .sr(N__82851));
endmodule // Pc2drone
