// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Apr 3 2019 22:10:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_drone,
    uart_data_rdy_debug,
    ppm_output,
    uart_input_pc,
    uart_input_debug,
    drone_frame_decoder_data_rdy_debug,
    clk_system);

    input uart_input_drone;
    output uart_data_rdy_debug;
    output ppm_output;
    input uart_input_pc;
    output uart_input_debug;
    output drone_frame_decoder_data_rdy_debug;
    input clk_system;

    wire N__26456;
    wire N__26455;
    wire N__26454;
    wire N__26445;
    wire N__26444;
    wire N__26443;
    wire N__26436;
    wire N__26435;
    wire N__26434;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26418;
    wire N__26417;
    wire N__26416;
    wire N__26409;
    wire N__26408;
    wire N__26407;
    wire N__26400;
    wire N__26399;
    wire N__26398;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26363;
    wire N__26362;
    wire N__26361;
    wire N__26360;
    wire N__26359;
    wire N__26356;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26332;
    wire N__26325;
    wire N__26322;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26310;
    wire N__26309;
    wire N__26304;
    wire N__26301;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26258;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26234;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26176;
    wire N__26175;
    wire N__26172;
    wire N__26171;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26111;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26092;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26079;
    wire N__26074;
    wire N__26073;
    wire N__26072;
    wire N__26071;
    wire N__26068;
    wire N__26067;
    wire N__26066;
    wire N__26065;
    wire N__26064;
    wire N__26063;
    wire N__26062;
    wire N__26059;
    wire N__26052;
    wire N__26049;
    wire N__26048;
    wire N__26043;
    wire N__26040;
    wire N__26035;
    wire N__26032;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26015;
    wire N__26012;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25983;
    wire N__25980;
    wire N__25979;
    wire N__25978;
    wire N__25975;
    wire N__25968;
    wire N__25957;
    wire N__25952;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25936;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25909;
    wire N__25898;
    wire N__25897;
    wire N__25896;
    wire N__25895;
    wire N__25894;
    wire N__25893;
    wire N__25892;
    wire N__25891;
    wire N__25886;
    wire N__25885;
    wire N__25884;
    wire N__25883;
    wire N__25880;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25843;
    wire N__25840;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25824;
    wire N__25819;
    wire N__25808;
    wire N__25807;
    wire N__25806;
    wire N__25805;
    wire N__25804;
    wire N__25801;
    wire N__25800;
    wire N__25797;
    wire N__25796;
    wire N__25795;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25787;
    wire N__25786;
    wire N__25785;
    wire N__25782;
    wire N__25781;
    wire N__25778;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25733;
    wire N__25732;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25714;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25687;
    wire N__25674;
    wire N__25669;
    wire N__25658;
    wire N__25657;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25642;
    wire N__25639;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25554;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25544;
    wire N__25543;
    wire N__25542;
    wire N__25537;
    wire N__25534;
    wire N__25533;
    wire N__25530;
    wire N__25529;
    wire N__25528;
    wire N__25525;
    wire N__25524;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25520;
    wire N__25517;
    wire N__25516;
    wire N__25513;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25505;
    wire N__25502;
    wire N__25497;
    wire N__25496;
    wire N__25495;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25481;
    wire N__25478;
    wire N__25477;
    wire N__25474;
    wire N__25473;
    wire N__25468;
    wire N__25461;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25443;
    wire N__25438;
    wire N__25435;
    wire N__25434;
    wire N__25431;
    wire N__25430;
    wire N__25429;
    wire N__25426;
    wire N__25425;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25411;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25391;
    wire N__25386;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25362;
    wire N__25359;
    wire N__25346;
    wire N__25343;
    wire N__25338;
    wire N__25335;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25304;
    wire N__25303;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25299;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25295;
    wire N__25294;
    wire N__25293;
    wire N__25292;
    wire N__25291;
    wire N__25290;
    wire N__25289;
    wire N__25288;
    wire N__25287;
    wire N__25286;
    wire N__25285;
    wire N__25284;
    wire N__25283;
    wire N__25282;
    wire N__25281;
    wire N__25280;
    wire N__25279;
    wire N__25278;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25271;
    wire N__25270;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25265;
    wire N__25264;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25255;
    wire N__25254;
    wire N__25253;
    wire N__25252;
    wire N__25251;
    wire N__25250;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25246;
    wire N__25245;
    wire N__25244;
    wire N__25243;
    wire N__25242;
    wire N__25241;
    wire N__25240;
    wire N__25239;
    wire N__25238;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25231;
    wire N__25230;
    wire N__25229;
    wire N__25228;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25224;
    wire N__25223;
    wire N__25222;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25210;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25206;
    wire N__25205;
    wire N__25204;
    wire N__25203;
    wire N__25202;
    wire N__25201;
    wire N__25200;
    wire N__25199;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25195;
    wire N__25194;
    wire N__25193;
    wire N__25192;
    wire N__25191;
    wire N__25190;
    wire N__25189;
    wire N__25188;
    wire N__25187;
    wire N__25186;
    wire N__25185;
    wire N__25184;
    wire N__25183;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24931;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24920;
    wire N__24919;
    wire N__24918;
    wire N__24917;
    wire N__24916;
    wire N__24913;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24906;
    wire N__24905;
    wire N__24904;
    wire N__24903;
    wire N__24902;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24898;
    wire N__24897;
    wire N__24896;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24816;
    wire N__24813;
    wire N__24812;
    wire N__24811;
    wire N__24810;
    wire N__24809;
    wire N__24808;
    wire N__24807;
    wire N__24806;
    wire N__24805;
    wire N__24804;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24793;
    wire N__24792;
    wire N__24791;
    wire N__24790;
    wire N__24789;
    wire N__24788;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24783;
    wire N__24782;
    wire N__24781;
    wire N__24780;
    wire N__24779;
    wire N__24778;
    wire N__24777;
    wire N__24776;
    wire N__24775;
    wire N__24774;
    wire N__24773;
    wire N__24772;
    wire N__24771;
    wire N__24770;
    wire N__24769;
    wire N__24768;
    wire N__24767;
    wire N__24766;
    wire N__24765;
    wire N__24764;
    wire N__24763;
    wire N__24762;
    wire N__24761;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24757;
    wire N__24756;
    wire N__24755;
    wire N__24754;
    wire N__24753;
    wire N__24752;
    wire N__24751;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24747;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24460;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24406;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24367;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24350;
    wire N__24349;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24332;
    wire N__24331;
    wire N__24328;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24293;
    wire N__24292;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24280;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24257;
    wire N__24256;
    wire N__24253;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24222;
    wire N__24215;
    wire N__24214;
    wire N__24213;
    wire N__24212;
    wire N__24211;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24203;
    wire N__24200;
    wire N__24199;
    wire N__24196;
    wire N__24195;
    wire N__24194;
    wire N__24193;
    wire N__24192;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24177;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24165;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24141;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24120;
    wire N__24119;
    wire N__24118;
    wire N__24117;
    wire N__24116;
    wire N__24111;
    wire N__24106;
    wire N__24101;
    wire N__24098;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24077;
    wire N__24072;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24056;
    wire N__24051;
    wire N__24046;
    wire N__24029;
    wire N__24028;
    wire N__24027;
    wire N__24024;
    wire N__24023;
    wire N__24020;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23995;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23978;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23932;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23915;
    wire N__23914;
    wire N__23913;
    wire N__23910;
    wire N__23905;
    wire N__23904;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23900;
    wire N__23899;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23876;
    wire N__23867;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23823;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23813;
    wire N__23808;
    wire N__23801;
    wire N__23798;
    wire N__23793;
    wire N__23792;
    wire N__23789;
    wire N__23788;
    wire N__23787;
    wire N__23784;
    wire N__23779;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23744;
    wire N__23739;
    wire N__23734;
    wire N__23731;
    wire N__23726;
    wire N__23721;
    wire N__23714;
    wire N__23713;
    wire N__23712;
    wire N__23711;
    wire N__23710;
    wire N__23709;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23705;
    wire N__23702;
    wire N__23701;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23694;
    wire N__23693;
    wire N__23692;
    wire N__23691;
    wire N__23690;
    wire N__23689;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23684;
    wire N__23683;
    wire N__23682;
    wire N__23681;
    wire N__23680;
    wire N__23679;
    wire N__23678;
    wire N__23677;
    wire N__23676;
    wire N__23675;
    wire N__23664;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23631;
    wire N__23630;
    wire N__23629;
    wire N__23628;
    wire N__23627;
    wire N__23618;
    wire N__23607;
    wire N__23602;
    wire N__23595;
    wire N__23594;
    wire N__23593;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23569;
    wire N__23560;
    wire N__23557;
    wire N__23556;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23545;
    wire N__23540;
    wire N__23531;
    wire N__23522;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23486;
    wire N__23481;
    wire N__23478;
    wire N__23471;
    wire N__23462;
    wire N__23455;
    wire N__23448;
    wire N__23443;
    wire N__23430;
    wire N__23421;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23310;
    wire N__23309;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23301;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23281;
    wire N__23278;
    wire N__23277;
    wire N__23276;
    wire N__23275;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23259;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23251;
    wire N__23246;
    wire N__23237;
    wire N__23232;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23212;
    wire N__23211;
    wire N__23210;
    wire N__23209;
    wire N__23208;
    wire N__23207;
    wire N__23206;
    wire N__23205;
    wire N__23202;
    wire N__23193;
    wire N__23192;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23172;
    wire N__23167;
    wire N__23166;
    wire N__23161;
    wire N__23160;
    wire N__23157;
    wire N__23156;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23132;
    wire N__23129;
    wire N__23120;
    wire N__23117;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23109;
    wire N__23108;
    wire N__23105;
    wire N__23098;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23036;
    wire N__23035;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23018;
    wire N__23017;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22994;
    wire N__22993;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22976;
    wire N__22975;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22955;
    wire N__22954;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22910;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22862;
    wire N__22861;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22841;
    wire N__22840;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22824;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22819;
    wire N__22816;
    wire N__22815;
    wire N__22814;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22800;
    wire N__22797;
    wire N__22796;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22788;
    wire N__22787;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22772;
    wire N__22771;
    wire N__22770;
    wire N__22761;
    wire N__22760;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22752;
    wire N__22751;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22735;
    wire N__22724;
    wire N__22719;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22701;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22688;
    wire N__22687;
    wire N__22684;
    wire N__22683;
    wire N__22678;
    wire N__22665;
    wire N__22656;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22629;
    wire N__22622;
    wire N__22619;
    wire N__22614;
    wire N__22611;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22561;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22549;
    wire N__22548;
    wire N__22545;
    wire N__22540;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22516;
    wire N__22511;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22499;
    wire N__22494;
    wire N__22491;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22459;
    wire N__22458;
    wire N__22455;
    wire N__22450;
    wire N__22445;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22414;
    wire N__22413;
    wire N__22410;
    wire N__22405;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22389;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22344;
    wire N__22341;
    wire N__22336;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22234;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22210;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22137;
    wire N__22136;
    wire N__22133;
    wire N__22128;
    wire N__22125;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22102;
    wire N__22099;
    wire N__22098;
    wire N__22095;
    wire N__22090;
    wire N__22085;
    wire N__22082;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22043;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22028;
    wire N__22025;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21965;
    wire N__21964;
    wire N__21961;
    wire N__21956;
    wire N__21955;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21920;
    wire N__21917;
    wire N__21916;
    wire N__21913;
    wire N__21904;
    wire N__21897;
    wire N__21894;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21871;
    wire N__21868;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21850;
    wire N__21849;
    wire N__21848;
    wire N__21843;
    wire N__21840;
    wire N__21835;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21739;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21731;
    wire N__21730;
    wire N__21727;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21707;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21680;
    wire N__21675;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21527;
    wire N__21524;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21450;
    wire N__21447;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21362;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21338;
    wire N__21335;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21317;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21069;
    wire N__21066;
    wire N__21065;
    wire N__21056;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21033;
    wire N__21026;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21018;
    wire N__21017;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20990;
    wire N__20989;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20976;
    wire N__20975;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20942;
    wire N__20935;
    wire N__20932;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20897;
    wire N__20894;
    wire N__20893;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20865;
    wire N__20862;
    wire N__20855;
    wire N__20852;
    wire N__20851;
    wire N__20850;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20788;
    wire N__20781;
    wire N__20778;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20766;
    wire N__20761;
    wire N__20758;
    wire N__20753;
    wire N__20750;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20728;
    wire N__20727;
    wire N__20726;
    wire N__20725;
    wire N__20722;
    wire N__20721;
    wire N__20720;
    wire N__20717;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20674;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20659;
    wire N__20656;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20614;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20588;
    wire N__20585;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20560;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20536;
    wire N__20535;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20527;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20497;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20440;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20421;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20407;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20359;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20323;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20248;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20233;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20200;
    wire N__20199;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20169;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20165;
    wire N__20162;
    wire N__20153;
    wire N__20148;
    wire N__20145;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20102;
    wire N__20101;
    wire N__20100;
    wire N__20097;
    wire N__20096;
    wire N__20093;
    wire N__20088;
    wire N__20085;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20026;
    wire N__20025;
    wire N__20024;
    wire N__20021;
    wire N__20014;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19995;
    wire N__19990;
    wire N__19989;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19933;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19904;
    wire N__19901;
    wire N__19900;
    wire N__19899;
    wire N__19898;
    wire N__19895;
    wire N__19890;
    wire N__19887;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19702;
    wire N__19701;
    wire N__19700;
    wire N__19699;
    wire N__19696;
    wire N__19695;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19667;
    wire N__19666;
    wire N__19663;
    wire N__19658;
    wire N__19653;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19634;
    wire N__19629;
    wire N__19622;
    wire N__19613;
    wire N__19606;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19563;
    wire N__19562;
    wire N__19561;
    wire N__19558;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19527;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19501;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19491;
    wire N__19488;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19473;
    wire N__19470;
    wire N__19465;
    wire N__19460;
    wire N__19451;
    wire N__19446;
    wire N__19443;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19417;
    wire N__19412;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19397;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19147;
    wire N__19146;
    wire N__19143;
    wire N__19138;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19084;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19072;
    wire N__19071;
    wire N__19068;
    wire N__19063;
    wire N__19058;
    wire N__19055;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18988;
    wire N__18987;
    wire N__18984;
    wire N__18979;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18773;
    wire N__18770;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18692;
    wire N__18691;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18674;
    wire N__18673;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18665;
    wire N__18660;
    wire N__18657;
    wire N__18656;
    wire N__18653;
    wire N__18648;
    wire N__18645;
    wire N__18644;
    wire N__18643;
    wire N__18638;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18603;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18536;
    wire N__18535;
    wire N__18532;
    wire N__18531;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18517;
    wire N__18514;
    wire N__18513;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18505;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18455;
    wire N__18454;
    wire N__18453;
    wire N__18452;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18444;
    wire N__18441;
    wire N__18440;
    wire N__18437;
    wire N__18436;
    wire N__18435;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18073;
    wire N__18070;
    wire N__18069;
    wire N__18066;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18054;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18040;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18025;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18010;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17995;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17980;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17965;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17915;
    wire N__17908;
    wire N__17905;
    wire N__17900;
    wire N__17897;
    wire N__17896;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17819;
    wire N__17816;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17798;
    wire N__17795;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17762;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17747;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17552;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17330;
    wire N__17327;
    wire N__17326;
    wire N__17325;
    wire N__17318;
    wire N__17315;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17278;
    wire N__17277;
    wire N__17270;
    wire N__17267;
    wire N__17266;
    wire N__17265;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17248;
    wire N__17247;
    wire N__17240;
    wire N__17237;
    wire N__17236;
    wire N__17235;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17146;
    wire N__17145;
    wire N__17142;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17112;
    wire N__17107;
    wire N__17102;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17094;
    wire N__17089;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16993;
    wire N__16992;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16975;
    wire N__16974;
    wire N__16971;
    wire N__16966;
    wire N__16961;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16919;
    wire N__16918;
    wire N__16917;
    wire N__16914;
    wire N__16909;
    wire N__16904;
    wire N__16903;
    wire N__16900;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16880;
    wire N__16877;
    wire N__16876;
    wire N__16873;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16853;
    wire N__16850;
    wire N__16849;
    wire N__16846;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16826;
    wire N__16823;
    wire N__16822;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16804;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16786;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16768;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16635;
    wire N__16632;
    wire N__16627;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16611;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16599;
    wire N__16592;
    wire N__16591;
    wire N__16588;
    wire N__16587;
    wire N__16584;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16564;
    wire N__16561;
    wire N__16556;
    wire N__16555;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16537;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16503;
    wire N__16502;
    wire N__16499;
    wire N__16494;
    wire N__16491;
    wire N__16486;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16474;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16459;
    wire N__16456;
    wire N__16455;
    wire N__16452;
    wire N__16451;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16327;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16312;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16297;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16282;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16201;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16179;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16165;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16128;
    wire N__16127;
    wire N__16126;
    wire N__16125;
    wire N__16124;
    wire N__16123;
    wire N__16120;
    wire N__16115;
    wire N__16108;
    wire N__16103;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16055;
    wire N__16052;
    wire N__16051;
    wire N__16050;
    wire N__16047;
    wire N__16042;
    wire N__16037;
    wire N__16034;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16019;
    wire N__16018;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16001;
    wire N__15998;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15986;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15978;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15964;
    wire N__15961;
    wire N__15956;
    wire N__15955;
    wire N__15954;
    wire N__15951;
    wire N__15946;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15625;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15617;
    wire N__15616;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15604;
    wire N__15599;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15580;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15568;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15530;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15518;
    wire N__15515;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15437;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15425;
    wire N__15422;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15407;
    wire N__15404;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15392;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15351;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15328;
    wire N__15327;
    wire N__15322;
    wire N__15319;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15315;
    wire N__15310;
    wire N__15309;
    wire N__15306;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15281;
    wire N__15280;
    wire N__15275;
    wire N__15272;
    wire N__15271;
    wire N__15270;
    wire N__15269;
    wire N__15268;
    wire N__15267;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15253;
    wire N__15252;
    wire N__15251;
    wire N__15248;
    wire N__15247;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15225;
    wire N__15222;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15167;
    wire N__15166;
    wire N__15165;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15086;
    wire N__15085;
    wire N__15082;
    wire N__15081;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15047;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15039;
    wire N__15038;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15020;
    wire N__15017;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14981;
    wire N__14978;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14809;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14791;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14770;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14758;
    wire N__14753;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14725;
    wire N__14722;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14705;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14697;
    wire N__14694;
    wire N__14693;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14606;
    wire N__14603;
    wire N__14602;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14524;
    wire N__14521;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14513;
    wire N__14512;
    wire N__14511;
    wire N__14510;
    wire N__14509;
    wire N__14506;
    wire N__14499;
    wire N__14490;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14368;
    wire N__14367;
    wire N__14364;
    wire N__14361;
    wire N__14356;
    wire N__14351;
    wire N__14350;
    wire N__14349;
    wire N__14348;
    wire N__14345;
    wire N__14338;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14297;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14281;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14269;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14099;
    wire N__14098;
    wire N__14097;
    wire N__14094;
    wire N__14089;
    wire N__14084;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14072;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14057;
    wire N__14056;
    wire N__14055;
    wire N__14052;
    wire N__14047;
    wire N__14042;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14008;
    wire N__14005;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13981;
    wire N__13978;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13961;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13934;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13922;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13907;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13841;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13829;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13762;
    wire N__13761;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13749;
    wire N__13746;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13495;
    wire N__13494;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13352;
    wire N__13349;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13331;
    wire N__13328;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13310;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13292;
    wire N__13289;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13277;
    wire N__13274;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13262;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13226;
    wire N__13225;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13215;
    wire N__13210;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13183;
    wire N__13182;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13174;
    wire N__13173;
    wire N__13170;
    wire N__13169;
    wire N__13166;
    wire N__13165;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13133;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13076;
    wire N__13073;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13055;
    wire N__13054;
    wire N__13053;
    wire N__13050;
    wire N__13045;
    wire N__13040;
    wire N__13039;
    wire N__13036;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13001;
    wire N__12992;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12980;
    wire N__12977;
    wire N__12972;
    wire N__12969;
    wire N__12964;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12929;
    wire N__12928;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12917;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12909;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12901;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12883;
    wire N__12878;
    wire N__12869;
    wire N__12868;
    wire N__12867;
    wire N__12866;
    wire N__12865;
    wire N__12864;
    wire N__12863;
    wire N__12862;
    wire N__12859;
    wire N__12844;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12808;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12769;
    wire N__12768;
    wire N__12765;
    wire N__12760;
    wire N__12759;
    wire N__12758;
    wire N__12757;
    wire N__12756;
    wire N__12755;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12737;
    wire N__12734;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12704;
    wire N__12703;
    wire N__12702;
    wire N__12701;
    wire N__12700;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12685;
    wire N__12682;
    wire N__12671;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12659;
    wire N__12656;
    wire N__12647;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12635;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12623;
    wire N__12622;
    wire N__12621;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12616;
    wire N__12615;
    wire N__12610;
    wire N__12599;
    wire N__12598;
    wire N__12597;
    wire N__12592;
    wire N__12587;
    wire N__12582;
    wire N__12575;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12529;
    wire N__12528;
    wire N__12527;
    wire N__12524;
    wire N__12523;
    wire N__12522;
    wire N__12519;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12500;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12473;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12456;
    wire N__12449;
    wire N__12448;
    wire N__12447;
    wire N__12446;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12442;
    wire N__12441;
    wire N__12436;
    wire N__12431;
    wire N__12424;
    wire N__12423;
    wire N__12422;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12403;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12374;
    wire N__12373;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12363;
    wire N__12358;
    wire N__12353;
    wire N__12346;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12309;
    wire N__12304;
    wire N__12297;
    wire N__12296;
    wire N__12295;
    wire N__12292;
    wire N__12287;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12273;
    wire N__12270;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12238;
    wire N__12233;
    wire N__12230;
    wire N__12225;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12208;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12200;
    wire N__12197;
    wire N__12192;
    wire N__12187;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12153;
    wire N__12148;
    wire N__12137;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12130;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12122;
    wire N__12119;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12104;
    wire N__12101;
    wire N__12094;
    wire N__12083;
    wire N__12082;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12056;
    wire N__12055;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12018;
    wire N__12017;
    wire N__12016;
    wire N__12015;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11995;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11974;
    wire N__11971;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11947;
    wire N__11942;
    wire N__11941;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11934;
    wire N__11929;
    wire N__11928;
    wire N__11927;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11912;
    wire N__11905;
    wire N__11902;
    wire N__11891;
    wire N__11888;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11866;
    wire N__11861;
    wire N__11860;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11856;
    wire N__11855;
    wire N__11852;
    wire N__11847;
    wire N__11838;
    wire N__11831;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11756;
    wire N__11751;
    wire N__11746;
    wire N__11741;
    wire N__11740;
    wire N__11739;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11731;
    wire N__11726;
    wire N__11721;
    wire N__11714;
    wire N__11711;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11692;
    wire N__11689;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11645;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11630;
    wire N__11627;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11609;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11577;
    wire N__11572;
    wire N__11567;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11532;
    wire N__11529;
    wire N__11522;
    wire N__11521;
    wire N__11520;
    wire N__11517;
    wire N__11512;
    wire N__11507;
    wire N__11506;
    wire N__11503;
    wire N__11502;
    wire N__11501;
    wire N__11496;
    wire N__11491;
    wire N__11486;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11480;
    wire N__11475;
    wire N__11470;
    wire N__11465;
    wire N__11462;
    wire N__11461;
    wire N__11458;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11436;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11383;
    wire N__11380;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11330;
    wire N__11327;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11315;
    wire N__11312;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11297;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11233;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11182;
    wire N__11179;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11164;
    wire N__11161;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11141;
    wire N__11138;
    wire N__11137;
    wire N__11136;
    wire N__11135;
    wire N__11134;
    wire N__11131;
    wire N__11122;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11094;
    wire N__11093;
    wire N__11090;
    wire N__11081;
    wire N__11076;
    wire N__11069;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11050;
    wire N__11049;
    wire N__11046;
    wire N__11041;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11025;
    wire N__11020;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10988;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10973;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10961;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10898;
    wire N__10895;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10883;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10811;
    wire N__10808;
    wire N__10807;
    wire N__10802;
    wire N__10799;
    wire N__10798;
    wire N__10795;
    wire N__10790;
    wire N__10787;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10775;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10763;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10751;
    wire N__10748;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10736;
    wire N__10735;
    wire N__10730;
    wire N__10727;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10712;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10697;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10654;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10589;
    wire N__10586;
    wire N__10585;
    wire N__10582;
    wire N__10581;
    wire N__10578;
    wire N__10573;
    wire N__10568;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10560;
    wire N__10555;
    wire N__10550;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10535;
    wire N__10532;
    wire N__10531;
    wire N__10530;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10379;
    wire N__10376;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10364;
    wire N__10361;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10349;
    wire N__10346;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10334;
    wire N__10331;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10319;
    wire N__10316;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10276;
    wire N__10273;
    wire N__10272;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10247;
    wire N__10238;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10220;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10150;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10138;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10124;
    wire VCCG0;
    wire GNDG0;
    wire \frame_dron_decoder_1.stateZ0Z_2 ;
    wire \frame_dron_decoder_1.stateZ0Z_5 ;
    wire \frame_dron_decoder_1.stateZ0Z_4 ;
    wire \frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4 ;
    wire \frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_ ;
    wire \frame_dron_decoder_1.WDT10lt14_0_cascade_ ;
    wire \frame_dron_decoder_1.WDT10lt14_0 ;
    wire \frame_dron_decoder_1.WDT10lto13_1 ;
    wire \frame_dron_decoder_1.stateZ0Z_7 ;
    wire \frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_ ;
    wire \frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_ ;
    wire \frame_dron_decoder_1.N_229_cascade_ ;
    wire \frame_dron_decoder_1.state_ns_i_a2_0_2_0 ;
    wire \frame_dron_decoder_1.N_231 ;
    wire \frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_ ;
    wire \frame_dron_decoder_1.state_ns_0_a3_0_3_1 ;
    wire \frame_dron_decoder_1.N_249 ;
    wire \frame_dron_decoder_1.stateZ0Z_3 ;
    wire \frame_dron_decoder_1.WDT10_0_i ;
    wire \frame_dron_decoder_1.WDTZ0Z_0 ;
    wire bfn_2_14_0_;
    wire \frame_dron_decoder_1.WDTZ0Z_1 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_0 ;
    wire \frame_dron_decoder_1.WDTZ0Z_2 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_1 ;
    wire \frame_dron_decoder_1.WDTZ0Z_3 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_2 ;
    wire \frame_dron_decoder_1.WDTZ0Z_4 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_3 ;
    wire \frame_dron_decoder_1.WDTZ0Z_5 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_4 ;
    wire \frame_dron_decoder_1.WDTZ0Z_6 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_5 ;
    wire \frame_dron_decoder_1.WDTZ0Z_7 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_6 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_7 ;
    wire \frame_dron_decoder_1.WDTZ0Z_8 ;
    wire bfn_2_15_0_;
    wire \frame_dron_decoder_1.WDTZ0Z_9 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_8 ;
    wire \frame_dron_decoder_1.WDTZ0Z_10 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_9 ;
    wire \frame_dron_decoder_1.WDTZ0Z_11 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_10 ;
    wire \frame_dron_decoder_1.WDTZ0Z_12 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_11 ;
    wire \frame_dron_decoder_1.WDTZ0Z_13 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_12 ;
    wire \frame_dron_decoder_1.WDTZ0Z_14 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_13 ;
    wire \frame_dron_decoder_1.un1_WDT_cry_14 ;
    wire \frame_dron_decoder_1.WDTZ0Z_15 ;
    wire \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3 ;
    wire \frame_dron_decoder_1.stateZ0Z_1 ;
    wire uart_drone_data_4;
    wire \frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_ ;
    wire \frame_dron_decoder_1.state_ns_0_a3_0_3_3 ;
    wire \frame_dron_decoder_1.stateZ0Z_0 ;
    wire \frame_dron_decoder_1.state_ns_i_a2_1_2_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire bfn_2_17_0_;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire bfn_2_18_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_2_19_0_;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.reset6_3_cascade_ ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_11 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.reset6_15_cascade_ ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.countZ0Z_2 ;
    wire \frame_dron_decoder_1.stateZ0Z_6 ;
    wire drone_frame_decoder_data_rdy_debug_c;
    wire uart_drone_data_2;
    wire \frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ;
    wire \frame_dron_decoder_1.N_255 ;
    wire uart_data_rdy_debug_c;
    wire \frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire uart_drone_data_1;
    wire uart_drone_data_3;
    wire uart_drone_data_0;
    wire uart_drone_data_5;
    wire uart_drone_data_6;
    wire uart_drone_data_7;
    wire \uart_drone.state_1_sqmuxa_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_Auxce_0_0_4_cascade_ ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.state_1_sqmuxa ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire bfn_3_19_0_;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.state_srsts_0_0_0 ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \uart_drone.un1_state_2_0 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \uart_drone.N_143_cascade_ ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.N_144_1 ;
    wire \uart_drone.N_144_1_cascade_ ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_145 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.N_152 ;
    wire uart_input_debug_c;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.CO0 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.un1_state_4_0_cascade_ ;
    wire \uart_pc.CO0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1 ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire bfn_5_18_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \uart_pc.data_AuxZ0Z_1 ;
    wire \uart_pc.data_AuxZ0Z_0 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_AuxZ0Z_2 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ;
    wire \uart_frame_decoder.WDTZ0Z_0 ;
    wire bfn_7_15_0_;
    wire \uart_frame_decoder.WDTZ0Z_1 ;
    wire \uart_frame_decoder.un1_WDT_cry_0 ;
    wire \uart_frame_decoder.WDTZ0Z_2 ;
    wire \uart_frame_decoder.un1_WDT_cry_1 ;
    wire \uart_frame_decoder.WDTZ0Z_3 ;
    wire \uart_frame_decoder.un1_WDT_cry_2 ;
    wire \uart_frame_decoder.un1_WDT_cry_3 ;
    wire \uart_frame_decoder.un1_WDT_cry_4 ;
    wire \uart_frame_decoder.un1_WDT_cry_5 ;
    wire \uart_frame_decoder.un1_WDT_cry_6 ;
    wire \uart_frame_decoder.un1_WDT_cry_7 ;
    wire bfn_7_16_0_;
    wire \uart_frame_decoder.un1_WDT_cry_8 ;
    wire \uart_frame_decoder.un1_WDT_cry_9 ;
    wire \uart_frame_decoder.un1_WDT_cry_10 ;
    wire \uart_frame_decoder.un1_WDT_cry_11 ;
    wire \uart_frame_decoder.un1_WDT_cry_12 ;
    wire \uart_frame_decoder.un1_WDT_cry_13 ;
    wire \uart_frame_decoder.un1_WDT_cry_14 ;
    wire \uart_frame_decoder.source_offset1data_1_sqmuxa_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ;
    wire bfn_7_26_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire bfn_7_27_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_7_28_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.N_138_4 ;
    wire \uart_frame_decoder.N_138_4_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ;
    wire \uart_frame_decoder.state_1Z0Z_1 ;
    wire \uart_frame_decoder.state_1_RNO_2Z0Z_0 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ;
    wire \uart_frame_decoder.N_85_cascade_ ;
    wire \uart_frame_decoder.state_1Z0Z_6 ;
    wire \uart_frame_decoder.source_offset1data_1_sqmuxa ;
    wire \uart_frame_decoder.state_1Z0Z_7 ;
    wire \uart_frame_decoder.source_offset2data_1_sqmuxa ;
    wire \uart_frame_decoder.state_1Z0Z_8 ;
    wire \uart_frame_decoder.source_offset3data_1_sqmuxa ;
    wire \uart_frame_decoder.source_offset2data_1_sqmuxa_0 ;
    wire \uart_frame_decoder.source_offset3data_1_sqmuxa_0 ;
    wire \uart_frame_decoder.WDTZ0Z_6 ;
    wire \uart_frame_decoder.WDTZ0Z_11 ;
    wire \uart_frame_decoder.WDTZ0Z_10 ;
    wire \uart_frame_decoder.WDTZ0Z_13 ;
    wire \uart_frame_decoder.WDTZ0Z_12 ;
    wire \uart_frame_decoder.WDTZ0Z_7 ;
    wire \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ;
    wire \uart_frame_decoder.WDT8lto13_1 ;
    wire \uart_frame_decoder.WDT8lt14_0 ;
    wire \uart_frame_decoder.WDTZ0Z_14 ;
    wire \uart_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \uart_frame_decoder.WDTZ0Z_15 ;
    wire \uart_frame_decoder.WDT8_0_i ;
    wire \uart_frame_decoder.WDTZ0Z_8 ;
    wire \uart_frame_decoder.WDTZ0Z_5 ;
    wire \uart_frame_decoder.WDTZ0Z_9 ;
    wire \uart_frame_decoder.WDTZ0Z_4 ;
    wire \uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ;
    wire \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ;
    wire bfn_8_17_0_;
    wire frame_decoder_CH1data_1;
    wire frame_decoder_OFF1data_1;
    wire \scaler_1.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH1data_2;
    wire frame_decoder_OFF1data_2;
    wire \scaler_1.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH1data_3;
    wire frame_decoder_OFF1data_3;
    wire \scaler_1.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH1data_4;
    wire frame_decoder_OFF1data_4;
    wire \scaler_1.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH1data_5;
    wire frame_decoder_OFF1data_5;
    wire \scaler_1.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH1data_6;
    wire frame_decoder_OFF1data_6;
    wire \scaler_1.un3_source_data_0_cry_5 ;
    wire \scaler_1.un3_source_data_0_cry_6 ;
    wire \scaler_1.un3_source_data_0_cry_7 ;
    wire bfn_8_18_0_;
    wire \scaler_1.un3_source_data_0_cry_8 ;
    wire \scaler_1.un3_source_data_0_axb_7 ;
    wire frame_decoder_CH1data_7;
    wire frame_decoder_OFF1data_7;
    wire \scaler_1.N_508_i_l_ofxZ0 ;
    wire \uart_frame_decoder.count_RNIHJ501Z0Z_0 ;
    wire bfn_8_19_0_;
    wire \uart_frame_decoder.count8_axb_1 ;
    wire \uart_frame_decoder.count8_cry_0 ;
    wire \uart_frame_decoder.count_i_2 ;
    wire \uart_frame_decoder.count8_cry_1 ;
    wire \uart_frame_decoder.count8 ;
    wire \uart_frame_decoder.source_CH1data_1_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.N_299 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.PPM_STATE_62_d_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_11_0_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ;
    wire \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.state_1_sqmuxa_0 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_frame_decoder.state_1_ns_i_i_0_0 ;
    wire \uart_frame_decoder.N_39_i_1 ;
    wire \uart_frame_decoder.state_1Z0Z_0 ;
    wire \uart_frame_decoder.state_1Z0Z_9 ;
    wire \uart_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ;
    wire \uart_frame_decoder.countZ0Z_2 ;
    wire \uart_frame_decoder.countZ0Z_1 ;
    wire \uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_o2_0_10 ;
    wire bfn_9_14_0_;
    wire frame_decoder_CH2data_1;
    wire frame_decoder_OFF2data_1;
    wire \scaler_2.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH2data_2;
    wire frame_decoder_OFF2data_2;
    wire \scaler_2.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH2data_3;
    wire frame_decoder_OFF2data_3;
    wire \scaler_2.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH2data_4;
    wire frame_decoder_OFF2data_4;
    wire \scaler_2.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH2data_5;
    wire frame_decoder_OFF2data_5;
    wire \scaler_2.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH2data_6;
    wire frame_decoder_OFF2data_6;
    wire \scaler_2.un3_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_7 ;
    wire bfn_9_15_0_;
    wire \scaler_2.un3_source_data_0_cry_8 ;
    wire \uart_frame_decoder.state_1Z0Z_3 ;
    wire \uart_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ;
    wire \scaler_2.N_520_i_l_ofxZ0 ;
    wire scaler_1_data_5;
    wire scaler_3_data_5;
    wire scaler_1_data_4;
    wire frame_decoder_OFF2data_0;
    wire frame_decoder_CH2data_0;
    wire scaler_2_data_4;
    wire scaler_3_data_4;
    wire scaler_4_data_4;
    wire \uart_frame_decoder.state_1Z0Z_10 ;
    wire \uart_frame_decoder.count8_THRU_CO ;
    wire uart_input_pc_sync;
    wire \uart_pc.state_1_sqmuxa ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.N_306_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4 ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5 ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.N_300_cascade_ ;
    wire scaler_2_data_5;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire bfn_9_24_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.throttle_RNIALN65Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.throttle_RNI5V123Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.init_pulses_RNI60223Z0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.throttle_RNIONI96Z0Z_8 ;
    wire bfn_9_25_0_;
    wire \ppm_encoder_1.throttle_RNITSI96Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire bfn_9_26_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_162_d ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \scaler_2.un2_source_data_0_cry_1_c_RNO_0 ;
    wire bfn_10_13_0_;
    wire \scaler_2.un2_source_data_0 ;
    wire \scaler_2.un2_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_1_c_RNILSPH ;
    wire \scaler_2.un2_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ;
    wire \scaler_2.un2_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ;
    wire \scaler_2.un2_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ;
    wire \scaler_2.un2_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ;
    wire \scaler_2.un2_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ;
    wire \scaler_2.un2_source_data_0_cry_7 ;
    wire \scaler_2.un2_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ;
    wire \scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ;
    wire bfn_10_14_0_;
    wire \scaler_2.un2_source_data_0_cry_9 ;
    wire scaler_4_data_5;
    wire frame_decoder_OFF3data_0;
    wire bfn_10_15_0_;
    wire frame_decoder_OFF3data_1;
    wire \scaler_3.un3_source_data_0_cry_0 ;
    wire frame_decoder_OFF3data_2;
    wire \scaler_3.un3_source_data_0_cry_1 ;
    wire frame_decoder_OFF3data_3;
    wire \scaler_3.un3_source_data_0_cry_2 ;
    wire frame_decoder_OFF3data_4;
    wire \scaler_3.un3_source_data_0_cry_3 ;
    wire frame_decoder_OFF3data_5;
    wire \scaler_3.un3_source_data_0_cry_4 ;
    wire frame_decoder_OFF3data_6;
    wire \scaler_3.un3_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_axb_7 ;
    wire \scaler_3.un3_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_7 ;
    wire bfn_10_16_0_;
    wire \scaler_3.un3_source_data_0_cry_8 ;
    wire \uart_frame_decoder.count8_0_i ;
    wire frame_decoder_OFF3data_7;
    wire \scaler_3.N_532_i_l_ofxZ0 ;
    wire \uart_frame_decoder.state_1_RNINMHJZ0Z_10 ;
    wire \uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61 ;
    wire \uart_frame_decoder.count8_0 ;
    wire frame_decoder_OFF1data_0;
    wire frame_decoder_CH1data_0;
    wire \scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_10_17_0_;
    wire \scaler_1.un2_source_data_0 ;
    wire \scaler_1.un2_source_data_0_cry_1 ;
    wire \scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ;
    wire \scaler_1.un2_source_data_0_cry_2 ;
    wire \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ;
    wire \scaler_1.un2_source_data_0_cry_3 ;
    wire \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ;
    wire \scaler_1.un2_source_data_0_cry_4 ;
    wire \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ;
    wire \scaler_1.un2_source_data_0_cry_5 ;
    wire \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ;
    wire \scaler_1.un2_source_data_0_cry_6 ;
    wire \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ;
    wire \scaler_1.un2_source_data_0_cry_7 ;
    wire \scaler_1.un2_source_data_0_cry_8 ;
    wire \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ;
    wire \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ;
    wire bfn_10_18_0_;
    wire \scaler_1.un2_source_data_0_cry_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.N_303_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.N_307 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIJII96Z0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.N_302 ;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ;
    wire \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10 ;
    wire \ppm_encoder_1.N_305_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13 ;
    wire \ppm_encoder_1.N_308_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire bfn_10_27_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_10_28_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire bfn_11_12_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire bfn_11_13_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \uart_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire frame_decoder_CH4data_0;
    wire frame_decoder_OFF4data_0;
    wire \scaler_4.N_544_i_l_ofxZ0 ;
    wire frame_decoder_OFF2data_7;
    wire \scaler_2.un3_source_data_0_axb_7 ;
    wire frame_decoder_CH2data_7;
    wire \uart_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire \uart_frame_decoder.state_1Z0Z_5 ;
    wire \uart_frame_decoder.source_CH4data_1_sqmuxa ;
    wire frame_decoder_OFF4data_7;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_3.un2_source_data_0_cry_1_c_RNO_1 ;
    wire bfn_11_15_0_;
    wire \scaler_3.un2_source_data_0 ;
    wire \scaler_3.un2_source_data_0_cry_1 ;
    wire \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ;
    wire \scaler_3.un2_source_data_0_cry_2 ;
    wire \scaler_3.un3_source_data_0_cry_2_c_RNIR08I ;
    wire \scaler_3.un2_source_data_0_cry_3 ;
    wire \scaler_3.un3_source_data_0_cry_3_c_RNIU49I ;
    wire \scaler_3.un2_source_data_0_cry_4 ;
    wire \scaler_3.un3_source_data_0_cry_4_c_RNI19AI ;
    wire \scaler_3.un2_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ;
    wire \scaler_3.un2_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ;
    wire \scaler_3.un2_source_data_0_cry_7 ;
    wire \scaler_3.un2_source_data_0_cry_8 ;
    wire \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ;
    wire \scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ;
    wire bfn_11_16_0_;
    wire \scaler_3.un2_source_data_0_cry_9 ;
    wire bfn_11_17_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_11_18_0_;
    wire scaler_3_data_6;
    wire bfn_11_19_0_;
    wire scaler_3_data_7;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire scaler_3_data_8;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire scaler_3_data_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire scaler_3_data_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire scaler_3_data_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire scaler_3_data_12;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire scaler_3_data_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire scaler_3_data_14;
    wire bfn_11_20_0_;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ;
    wire \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire scaler_2_data_6;
    wire bfn_11_24_0_;
    wire scaler_2_data_7;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire scaler_2_data_8;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire scaler_2_data_9;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire scaler_2_data_10;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire scaler_2_data_11;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire scaler_2_data_12;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire scaler_2_data_14;
    wire bfn_11_25_0_;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.N_614_i ;
    wire bfn_11_28_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_11_29_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_11_30_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_228_g ;
    wire pc_frame_decoder_dv;
    wire pc_frame_decoder_dv_0;
    wire frame_decoder_OFF4data_4;
    wire \uart_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNO_2 ;
    wire bfn_12_13_0_;
    wire \scaler_4.un2_source_data_0 ;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ;
    wire scaler_4_data_7;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ;
    wire scaler_4_data_8;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNI15MI ;
    wire scaler_4_data_9;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNI49NI ;
    wire scaler_4_data_10;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire scaler_4_data_13;
    wire bfn_12_14_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire pc_frame_decoder_dv_0_g;
    wire uart_pc_data_0;
    wire frame_decoder_CH3data_0;
    wire uart_pc_data_1;
    wire frame_decoder_CH3data_1;
    wire uart_pc_data_2;
    wire frame_decoder_CH3data_2;
    wire uart_pc_data_3;
    wire frame_decoder_CH3data_3;
    wire uart_pc_data_4;
    wire frame_decoder_CH3data_4;
    wire uart_pc_data_6;
    wire frame_decoder_CH3data_6;
    wire uart_pc_data_7;
    wire frame_decoder_CH3data_7;
    wire \uart_frame_decoder.source_CH1data_1_sqmuxa ;
    wire scaler_1_data_6;
    wire bfn_12_17_0_;
    wire scaler_1_data_7;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire scaler_1_data_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire scaler_1_data_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire scaler_1_data_13;
    wire CONSTANT_ONE_NET;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire scaler_1_data_14;
    wire bfn_12_18_0_;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.scaler_1_dv_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire scaler_1_data_8;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire scaler_1_data_10;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.N_143_0 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire ppm_output_c;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire scaler_1_data_9;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.N_309 ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.N_301 ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.N_323_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.N_322 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.PPM_STATE_62_d ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.N_148_17_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \ppm_encoder_1.N_148_17 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.N_148 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \ppm_encoder_1.N_241 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire reset_system;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_2 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ;
    wire \uart_frame_decoder.N_85 ;
    wire \uart_frame_decoder.state_1Z0Z_2 ;
    wire \uart_frame_decoder.state_1Z0Z_4 ;
    wire uart_pc_data_rdy;
    wire \uart_frame_decoder.source_CH3data_1_sqmuxa ;
    wire uart_pc_data_5;
    wire frame_decoder_CH3data_5;
    wire \uart_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire scaler_4_data_6;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.N_614_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.N_230 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.N_304 ;
    wire scaler_2_data_13;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire scaler_1_dv;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire reset_system_g;

    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__26454),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__26456),
            .DIN(N__26455),
            .DOUT(N__26454),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__26456),
            .PADOUT(N__26455),
            .PADIN(N__26454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__26445),
            .DIN(N__26444),
            .DOUT(N__26443),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__26445),
            .PADOUT(N__26444),
            .PADIN(N__26443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__26436),
            .DIN(N__26435),
            .DOUT(N__26434),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__26436),
            .PADOUT(N__26435),
            .PADIN(N__26434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__26427),
            .DIN(N__26426),
            .DOUT(N__26425),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__26427),
            .PADOUT(N__26426),
            .PADIN(N__26425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam drone_frame_decoder_data_rdy_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD drone_frame_decoder_data_rdy_debug_obuf_iopad (
            .OE(N__26418),
            .DIN(N__26417),
            .DOUT(N__26416),
            .PACKAGEPIN(drone_frame_decoder_data_rdy_debug));
    defparam drone_frame_decoder_data_rdy_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam drone_frame_decoder_data_rdy_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO drone_frame_decoder_data_rdy_debug_obuf_preio (
            .PADOEN(N__26418),
            .PADOUT(N__26417),
            .PADIN(N__26416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_debug_obuf_iopad (
            .OE(N__26409),
            .DIN(N__26408),
            .DOUT(N__26407),
            .PACKAGEPIN(uart_input_debug));
    defparam uart_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_input_debug_obuf_preio (
            .PADOEN(N__26409),
            .PADOUT(N__26408),
            .PADIN(N__26407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_data_rdy_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_data_rdy_debug_obuf_iopad (
            .OE(N__26400),
            .DIN(N__26399),
            .DOUT(N__26398),
            .PACKAGEPIN(uart_data_rdy_debug));
    defparam uart_data_rdy_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_data_rdy_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_data_rdy_debug_obuf_preio (
            .PADOEN(N__26400),
            .PADOUT(N__26399),
            .PADIN(N__26398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__6282 (
            .O(N__26381),
            .I(N__26378));
    LocalMux I__6281 (
            .O(N__26378),
            .I(N__26375));
    Span4Mux_h I__6280 (
            .O(N__26375),
            .I(N__26371));
    InMux I__6279 (
            .O(N__26374),
            .I(N__26368));
    Odrv4 I__6278 (
            .O(N__26371),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa ));
    LocalMux I__6277 (
            .O(N__26368),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__6276 (
            .O(N__26363),
            .I(N__26356));
    InMux I__6275 (
            .O(N__26362),
            .I(N__26352));
    InMux I__6274 (
            .O(N__26361),
            .I(N__26349));
    InMux I__6273 (
            .O(N__26360),
            .I(N__26346));
    InMux I__6272 (
            .O(N__26359),
            .I(N__26343));
    LocalMux I__6271 (
            .O(N__26356),
            .I(N__26339));
    InMux I__6270 (
            .O(N__26355),
            .I(N__26336));
    LocalMux I__6269 (
            .O(N__26352),
            .I(N__26333));
    LocalMux I__6268 (
            .O(N__26349),
            .I(N__26325));
    LocalMux I__6267 (
            .O(N__26346),
            .I(N__26325));
    LocalMux I__6266 (
            .O(N__26343),
            .I(N__26325));
    InMux I__6265 (
            .O(N__26342),
            .I(N__26322));
    Span4Mux_v I__6264 (
            .O(N__26339),
            .I(N__26317));
    LocalMux I__6263 (
            .O(N__26336),
            .I(N__26317));
    Span4Mux_v I__6262 (
            .O(N__26333),
            .I(N__26314));
    InMux I__6261 (
            .O(N__26332),
            .I(N__26311));
    Span4Mux_v I__6260 (
            .O(N__26325),
            .I(N__26304));
    LocalMux I__6259 (
            .O(N__26322),
            .I(N__26304));
    Span4Mux_h I__6258 (
            .O(N__26317),
            .I(N__26301));
    Sp12to4 I__6257 (
            .O(N__26314),
            .I(N__26296));
    LocalMux I__6256 (
            .O(N__26311),
            .I(N__26296));
    InMux I__6255 (
            .O(N__26310),
            .I(N__26293));
    InMux I__6254 (
            .O(N__26309),
            .I(N__26290));
    Odrv4 I__6253 (
            .O(N__26304),
            .I(uart_pc_data_5));
    Odrv4 I__6252 (
            .O(N__26301),
            .I(uart_pc_data_5));
    Odrv12 I__6251 (
            .O(N__26296),
            .I(uart_pc_data_5));
    LocalMux I__6250 (
            .O(N__26293),
            .I(uart_pc_data_5));
    LocalMux I__6249 (
            .O(N__26290),
            .I(uart_pc_data_5));
    InMux I__6248 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__6247 (
            .O(N__26276),
            .I(N__26273));
    Odrv4 I__6246 (
            .O(N__26273),
            .I(frame_decoder_CH3data_5));
    CEMux I__6245 (
            .O(N__26270),
            .I(N__26266));
    CEMux I__6244 (
            .O(N__26269),
            .I(N__26263));
    LocalMux I__6243 (
            .O(N__26266),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    LocalMux I__6242 (
            .O(N__26263),
            .I(\uart_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__6241 (
            .O(N__26258),
            .I(N__26254));
    InMux I__6240 (
            .O(N__26257),
            .I(N__26251));
    LocalMux I__6239 (
            .O(N__26254),
            .I(N__26248));
    LocalMux I__6238 (
            .O(N__26251),
            .I(N__26245));
    Span4Mux_v I__6237 (
            .O(N__26248),
            .I(N__26242));
    Span4Mux_v I__6236 (
            .O(N__26245),
            .I(N__26239));
    Odrv4 I__6235 (
            .O(N__26242),
            .I(scaler_4_data_6));
    Odrv4 I__6234 (
            .O(N__26239),
            .I(scaler_4_data_6));
    InMux I__6233 (
            .O(N__26234),
            .I(N__26230));
    InMux I__6232 (
            .O(N__26233),
            .I(N__26227));
    LocalMux I__6231 (
            .O(N__26230),
            .I(N__26223));
    LocalMux I__6230 (
            .O(N__26227),
            .I(N__26220));
    InMux I__6229 (
            .O(N__26226),
            .I(N__26217));
    Span4Mux_v I__6228 (
            .O(N__26223),
            .I(N__26214));
    Span4Mux_v I__6227 (
            .O(N__26220),
            .I(N__26211));
    LocalMux I__6226 (
            .O(N__26217),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__6225 (
            .O(N__26214),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__6224 (
            .O(N__26211),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__6223 (
            .O(N__26204),
            .I(N__26201));
    LocalMux I__6222 (
            .O(N__26201),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__6221 (
            .O(N__26198),
            .I(N__26195));
    LocalMux I__6220 (
            .O(N__26195),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    InMux I__6219 (
            .O(N__26192),
            .I(N__26189));
    LocalMux I__6218 (
            .O(N__26189),
            .I(N__26186));
    Span4Mux_h I__6217 (
            .O(N__26186),
            .I(N__26183));
    Span4Mux_v I__6216 (
            .O(N__26183),
            .I(N__26180));
    Odrv4 I__6215 (
            .O(N__26180),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CEMux I__6214 (
            .O(N__26177),
            .I(N__26172));
    CEMux I__6213 (
            .O(N__26176),
            .I(N__26168));
    CEMux I__6212 (
            .O(N__26175),
            .I(N__26164));
    LocalMux I__6211 (
            .O(N__26172),
            .I(N__26161));
    CEMux I__6210 (
            .O(N__26171),
            .I(N__26157));
    LocalMux I__6209 (
            .O(N__26168),
            .I(N__26154));
    CEMux I__6208 (
            .O(N__26167),
            .I(N__26151));
    LocalMux I__6207 (
            .O(N__26164),
            .I(N__26148));
    Span4Mux_h I__6206 (
            .O(N__26161),
            .I(N__26145));
    CEMux I__6205 (
            .O(N__26160),
            .I(N__26142));
    LocalMux I__6204 (
            .O(N__26157),
            .I(N__26139));
    Span4Mux_h I__6203 (
            .O(N__26154),
            .I(N__26136));
    LocalMux I__6202 (
            .O(N__26151),
            .I(N__26133));
    Span4Mux_v I__6201 (
            .O(N__26148),
            .I(N__26130));
    Span4Mux_s1_v I__6200 (
            .O(N__26145),
            .I(N__26127));
    LocalMux I__6199 (
            .O(N__26142),
            .I(N__26124));
    Span4Mux_h I__6198 (
            .O(N__26139),
            .I(N__26121));
    Span4Mux_h I__6197 (
            .O(N__26136),
            .I(N__26118));
    Span4Mux_v I__6196 (
            .O(N__26133),
            .I(N__26111));
    Span4Mux_v I__6195 (
            .O(N__26130),
            .I(N__26111));
    Span4Mux_v I__6194 (
            .O(N__26127),
            .I(N__26111));
    Odrv4 I__6193 (
            .O(N__26124),
            .I(\ppm_encoder_1.N_614_0 ));
    Odrv4 I__6192 (
            .O(N__26121),
            .I(\ppm_encoder_1.N_614_0 ));
    Odrv4 I__6191 (
            .O(N__26118),
            .I(\ppm_encoder_1.N_614_0 ));
    Odrv4 I__6190 (
            .O(N__26111),
            .I(\ppm_encoder_1.N_614_0 ));
    InMux I__6189 (
            .O(N__26102),
            .I(N__26096));
    InMux I__6188 (
            .O(N__26101),
            .I(N__26093));
    CascadeMux I__6187 (
            .O(N__26100),
            .I(N__26087));
    InMux I__6186 (
            .O(N__26099),
            .I(N__26084));
    LocalMux I__6185 (
            .O(N__26096),
            .I(N__26079));
    LocalMux I__6184 (
            .O(N__26093),
            .I(N__26079));
    InMux I__6183 (
            .O(N__26092),
            .I(N__26074));
    InMux I__6182 (
            .O(N__26091),
            .I(N__26074));
    CascadeMux I__6181 (
            .O(N__26090),
            .I(N__26068));
    InMux I__6180 (
            .O(N__26087),
            .I(N__26059));
    LocalMux I__6179 (
            .O(N__26084),
            .I(N__26052));
    Span4Mux_h I__6178 (
            .O(N__26079),
            .I(N__26052));
    LocalMux I__6177 (
            .O(N__26074),
            .I(N__26052));
    InMux I__6176 (
            .O(N__26073),
            .I(N__26049));
    InMux I__6175 (
            .O(N__26072),
            .I(N__26043));
    InMux I__6174 (
            .O(N__26071),
            .I(N__26043));
    InMux I__6173 (
            .O(N__26068),
            .I(N__26040));
    InMux I__6172 (
            .O(N__26067),
            .I(N__26035));
    InMux I__6171 (
            .O(N__26066),
            .I(N__26035));
    CascadeMux I__6170 (
            .O(N__26065),
            .I(N__26032));
    InMux I__6169 (
            .O(N__26064),
            .I(N__26028));
    InMux I__6168 (
            .O(N__26063),
            .I(N__26025));
    InMux I__6167 (
            .O(N__26062),
            .I(N__26022));
    LocalMux I__6166 (
            .O(N__26059),
            .I(N__26015));
    Span4Mux_h I__6165 (
            .O(N__26052),
            .I(N__26015));
    LocalMux I__6164 (
            .O(N__26049),
            .I(N__26015));
    InMux I__6163 (
            .O(N__26048),
            .I(N__26012));
    LocalMux I__6162 (
            .O(N__26043),
            .I(N__26008));
    LocalMux I__6161 (
            .O(N__26040),
            .I(N__26005));
    LocalMux I__6160 (
            .O(N__26035),
            .I(N__26002));
    InMux I__6159 (
            .O(N__26032),
            .I(N__25997));
    InMux I__6158 (
            .O(N__26031),
            .I(N__25997));
    LocalMux I__6157 (
            .O(N__26028),
            .I(N__25994));
    LocalMux I__6156 (
            .O(N__26025),
            .I(N__25991));
    LocalMux I__6155 (
            .O(N__26022),
            .I(N__25988));
    Span4Mux_v I__6154 (
            .O(N__26015),
            .I(N__25983));
    LocalMux I__6153 (
            .O(N__26012),
            .I(N__25983));
    InMux I__6152 (
            .O(N__26011),
            .I(N__25980));
    Span12Mux_v I__6151 (
            .O(N__26008),
            .I(N__25975));
    Span4Mux_h I__6150 (
            .O(N__26005),
            .I(N__25968));
    Span4Mux_v I__6149 (
            .O(N__26002),
            .I(N__25968));
    LocalMux I__6148 (
            .O(N__25997),
            .I(N__25968));
    Span4Mux_v I__6147 (
            .O(N__25994),
            .I(N__25957));
    Span4Mux_h I__6146 (
            .O(N__25991),
            .I(N__25957));
    Span4Mux_v I__6145 (
            .O(N__25988),
            .I(N__25957));
    Span4Mux_v I__6144 (
            .O(N__25983),
            .I(N__25957));
    LocalMux I__6143 (
            .O(N__25980),
            .I(N__25957));
    InMux I__6142 (
            .O(N__25979),
            .I(N__25952));
    InMux I__6141 (
            .O(N__25978),
            .I(N__25952));
    Odrv12 I__6140 (
            .O(N__25975),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6139 (
            .O(N__25968),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__6138 (
            .O(N__25957),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__6137 (
            .O(N__25952),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__6136 (
            .O(N__25943),
            .I(N__25940));
    LocalMux I__6135 (
            .O(N__25940),
            .I(N__25937));
    Span4Mux_h I__6134 (
            .O(N__25937),
            .I(N__25933));
    CascadeMux I__6133 (
            .O(N__25936),
            .I(N__25926));
    Span4Mux_v I__6132 (
            .O(N__25933),
            .I(N__25923));
    InMux I__6131 (
            .O(N__25932),
            .I(N__25920));
    InMux I__6130 (
            .O(N__25931),
            .I(N__25917));
    InMux I__6129 (
            .O(N__25930),
            .I(N__25914));
    InMux I__6128 (
            .O(N__25929),
            .I(N__25909));
    InMux I__6127 (
            .O(N__25926),
            .I(N__25909));
    Odrv4 I__6126 (
            .O(N__25923),
            .I(\ppm_encoder_1.N_230 ));
    LocalMux I__6125 (
            .O(N__25920),
            .I(\ppm_encoder_1.N_230 ));
    LocalMux I__6124 (
            .O(N__25917),
            .I(\ppm_encoder_1.N_230 ));
    LocalMux I__6123 (
            .O(N__25914),
            .I(\ppm_encoder_1.N_230 ));
    LocalMux I__6122 (
            .O(N__25909),
            .I(\ppm_encoder_1.N_230 ));
    InMux I__6121 (
            .O(N__25898),
            .I(N__25886));
    InMux I__6120 (
            .O(N__25897),
            .I(N__25886));
    InMux I__6119 (
            .O(N__25896),
            .I(N__25880));
    InMux I__6118 (
            .O(N__25895),
            .I(N__25873));
    InMux I__6117 (
            .O(N__25894),
            .I(N__25873));
    InMux I__6116 (
            .O(N__25893),
            .I(N__25873));
    InMux I__6115 (
            .O(N__25892),
            .I(N__25870));
    InMux I__6114 (
            .O(N__25891),
            .I(N__25867));
    LocalMux I__6113 (
            .O(N__25886),
            .I(N__25864));
    InMux I__6112 (
            .O(N__25885),
            .I(N__25854));
    InMux I__6111 (
            .O(N__25884),
            .I(N__25854));
    InMux I__6110 (
            .O(N__25883),
            .I(N__25854));
    LocalMux I__6109 (
            .O(N__25880),
            .I(N__25851));
    LocalMux I__6108 (
            .O(N__25873),
            .I(N__25848));
    LocalMux I__6107 (
            .O(N__25870),
            .I(N__25843));
    LocalMux I__6106 (
            .O(N__25867),
            .I(N__25843));
    Span4Mux_v I__6105 (
            .O(N__25864),
            .I(N__25840));
    InMux I__6104 (
            .O(N__25863),
            .I(N__25835));
    InMux I__6103 (
            .O(N__25862),
            .I(N__25835));
    InMux I__6102 (
            .O(N__25861),
            .I(N__25832));
    LocalMux I__6101 (
            .O(N__25854),
            .I(N__25829));
    Span4Mux_v I__6100 (
            .O(N__25851),
            .I(N__25824));
    Span4Mux_h I__6099 (
            .O(N__25848),
            .I(N__25824));
    Span4Mux_h I__6098 (
            .O(N__25843),
            .I(N__25819));
    Span4Mux_h I__6097 (
            .O(N__25840),
            .I(N__25819));
    LocalMux I__6096 (
            .O(N__25835),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__6095 (
            .O(N__25832),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv4 I__6094 (
            .O(N__25829),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv4 I__6093 (
            .O(N__25824),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv4 I__6092 (
            .O(N__25819),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__6091 (
            .O(N__25808),
            .I(N__25801));
    CascadeMux I__6090 (
            .O(N__25807),
            .I(N__25797));
    InMux I__6089 (
            .O(N__25806),
            .I(N__25791));
    InMux I__6088 (
            .O(N__25805),
            .I(N__25788));
    CascadeMux I__6087 (
            .O(N__25804),
            .I(N__25782));
    LocalMux I__6086 (
            .O(N__25801),
            .I(N__25778));
    InMux I__6085 (
            .O(N__25800),
            .I(N__25774));
    InMux I__6084 (
            .O(N__25797),
            .I(N__25771));
    InMux I__6083 (
            .O(N__25796),
            .I(N__25768));
    InMux I__6082 (
            .O(N__25795),
            .I(N__25765));
    InMux I__6081 (
            .O(N__25794),
            .I(N__25762));
    LocalMux I__6080 (
            .O(N__25791),
            .I(N__25757));
    LocalMux I__6079 (
            .O(N__25788),
            .I(N__25757));
    InMux I__6078 (
            .O(N__25787),
            .I(N__25754));
    InMux I__6077 (
            .O(N__25786),
            .I(N__25751));
    InMux I__6076 (
            .O(N__25785),
            .I(N__25748));
    InMux I__6075 (
            .O(N__25782),
            .I(N__25742));
    InMux I__6074 (
            .O(N__25781),
            .I(N__25742));
    Span4Mux_v I__6073 (
            .O(N__25778),
            .I(N__25739));
    InMux I__6072 (
            .O(N__25777),
            .I(N__25736));
    LocalMux I__6071 (
            .O(N__25774),
            .I(N__25727));
    LocalMux I__6070 (
            .O(N__25771),
            .I(N__25727));
    LocalMux I__6069 (
            .O(N__25768),
            .I(N__25724));
    LocalMux I__6068 (
            .O(N__25765),
            .I(N__25721));
    LocalMux I__6067 (
            .O(N__25762),
            .I(N__25714));
    Span4Mux_v I__6066 (
            .O(N__25757),
            .I(N__25714));
    LocalMux I__6065 (
            .O(N__25754),
            .I(N__25714));
    LocalMux I__6064 (
            .O(N__25751),
            .I(N__25709));
    LocalMux I__6063 (
            .O(N__25748),
            .I(N__25709));
    InMux I__6062 (
            .O(N__25747),
            .I(N__25706));
    LocalMux I__6061 (
            .O(N__25742),
            .I(N__25703));
    Span4Mux_v I__6060 (
            .O(N__25739),
            .I(N__25698));
    LocalMux I__6059 (
            .O(N__25736),
            .I(N__25698));
    InMux I__6058 (
            .O(N__25735),
            .I(N__25695));
    InMux I__6057 (
            .O(N__25734),
            .I(N__25692));
    InMux I__6056 (
            .O(N__25733),
            .I(N__25687));
    InMux I__6055 (
            .O(N__25732),
            .I(N__25687));
    Span4Mux_h I__6054 (
            .O(N__25727),
            .I(N__25674));
    Span4Mux_v I__6053 (
            .O(N__25724),
            .I(N__25674));
    Span4Mux_v I__6052 (
            .O(N__25721),
            .I(N__25674));
    Span4Mux_v I__6051 (
            .O(N__25714),
            .I(N__25674));
    Span4Mux_v I__6050 (
            .O(N__25709),
            .I(N__25674));
    LocalMux I__6049 (
            .O(N__25706),
            .I(N__25674));
    Span4Mux_v I__6048 (
            .O(N__25703),
            .I(N__25669));
    Span4Mux_h I__6047 (
            .O(N__25698),
            .I(N__25669));
    LocalMux I__6046 (
            .O(N__25695),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__6045 (
            .O(N__25692),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__6044 (
            .O(N__25687),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__6043 (
            .O(N__25674),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__6042 (
            .O(N__25669),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__6041 (
            .O(N__25658),
            .I(N__25653));
    InMux I__6040 (
            .O(N__25657),
            .I(N__25650));
    CascadeMux I__6039 (
            .O(N__25656),
            .I(N__25647));
    LocalMux I__6038 (
            .O(N__25653),
            .I(N__25642));
    LocalMux I__6037 (
            .O(N__25650),
            .I(N__25642));
    InMux I__6036 (
            .O(N__25647),
            .I(N__25639));
    Odrv12 I__6035 (
            .O(N__25642),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__6034 (
            .O(N__25639),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__6033 (
            .O(N__25634),
            .I(N__25629));
    InMux I__6032 (
            .O(N__25633),
            .I(N__25626));
    InMux I__6031 (
            .O(N__25632),
            .I(N__25623));
    LocalMux I__6030 (
            .O(N__25629),
            .I(N__25620));
    LocalMux I__6029 (
            .O(N__25626),
            .I(N__25617));
    LocalMux I__6028 (
            .O(N__25623),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__6027 (
            .O(N__25620),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__6026 (
            .O(N__25617),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__6025 (
            .O(N__25610),
            .I(N__25607));
    LocalMux I__6024 (
            .O(N__25607),
            .I(N__25604));
    Span4Mux_h I__6023 (
            .O(N__25604),
            .I(N__25601));
    Odrv4 I__6022 (
            .O(N__25601),
            .I(\ppm_encoder_1.N_304 ));
    InMux I__6021 (
            .O(N__25598),
            .I(N__25595));
    LocalMux I__6020 (
            .O(N__25595),
            .I(N__25592));
    Span4Mux_v I__6019 (
            .O(N__25592),
            .I(N__25588));
    InMux I__6018 (
            .O(N__25591),
            .I(N__25585));
    Span4Mux_h I__6017 (
            .O(N__25588),
            .I(N__25580));
    LocalMux I__6016 (
            .O(N__25585),
            .I(N__25580));
    Span4Mux_v I__6015 (
            .O(N__25580),
            .I(N__25577));
    Span4Mux_v I__6014 (
            .O(N__25577),
            .I(N__25574));
    Odrv4 I__6013 (
            .O(N__25574),
            .I(scaler_2_data_13));
    InMux I__6012 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__6011 (
            .O(N__25568),
            .I(N__25565));
    Span4Mux_h I__6010 (
            .O(N__25565),
            .I(N__25562));
    Odrv4 I__6009 (
            .O(N__25562),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    CascadeMux I__6008 (
            .O(N__25559),
            .I(N__25555));
    CascadeMux I__6007 (
            .O(N__25558),
            .I(N__25551));
    InMux I__6006 (
            .O(N__25555),
            .I(N__25537));
    InMux I__6005 (
            .O(N__25554),
            .I(N__25537));
    InMux I__6004 (
            .O(N__25551),
            .I(N__25534));
    CascadeMux I__6003 (
            .O(N__25550),
            .I(N__25530));
    CascadeMux I__6002 (
            .O(N__25549),
            .I(N__25525));
    CascadeMux I__6001 (
            .O(N__25548),
            .I(N__25517));
    CascadeMux I__6000 (
            .O(N__25547),
            .I(N__25513));
    CascadeMux I__5999 (
            .O(N__25546),
            .I(N__25509));
    CascadeMux I__5998 (
            .O(N__25545),
            .I(N__25506));
    CascadeMux I__5997 (
            .O(N__25544),
            .I(N__25502));
    InMux I__5996 (
            .O(N__25543),
            .I(N__25497));
    InMux I__5995 (
            .O(N__25542),
            .I(N__25497));
    LocalMux I__5994 (
            .O(N__25537),
            .I(N__25491));
    LocalMux I__5993 (
            .O(N__25534),
            .I(N__25488));
    InMux I__5992 (
            .O(N__25533),
            .I(N__25485));
    InMux I__5991 (
            .O(N__25530),
            .I(N__25482));
    CascadeMux I__5990 (
            .O(N__25529),
            .I(N__25478));
    CascadeMux I__5989 (
            .O(N__25528),
            .I(N__25474));
    InMux I__5988 (
            .O(N__25525),
            .I(N__25468));
    InMux I__5987 (
            .O(N__25524),
            .I(N__25468));
    InMux I__5986 (
            .O(N__25523),
            .I(N__25461));
    InMux I__5985 (
            .O(N__25522),
            .I(N__25461));
    InMux I__5984 (
            .O(N__25521),
            .I(N__25461));
    InMux I__5983 (
            .O(N__25520),
            .I(N__25454));
    InMux I__5982 (
            .O(N__25517),
            .I(N__25454));
    InMux I__5981 (
            .O(N__25516),
            .I(N__25454));
    InMux I__5980 (
            .O(N__25513),
            .I(N__25451));
    InMux I__5979 (
            .O(N__25512),
            .I(N__25448));
    InMux I__5978 (
            .O(N__25509),
            .I(N__25443));
    InMux I__5977 (
            .O(N__25506),
            .I(N__25443));
    InMux I__5976 (
            .O(N__25505),
            .I(N__25438));
    InMux I__5975 (
            .O(N__25502),
            .I(N__25438));
    LocalMux I__5974 (
            .O(N__25497),
            .I(N__25435));
    CascadeMux I__5973 (
            .O(N__25496),
            .I(N__25431));
    CascadeMux I__5972 (
            .O(N__25495),
            .I(N__25426));
    CascadeMux I__5971 (
            .O(N__25494),
            .I(N__25421));
    Span4Mux_v I__5970 (
            .O(N__25491),
            .I(N__25418));
    Span4Mux_v I__5969 (
            .O(N__25488),
            .I(N__25411));
    LocalMux I__5968 (
            .O(N__25485),
            .I(N__25411));
    LocalMux I__5967 (
            .O(N__25482),
            .I(N__25411));
    InMux I__5966 (
            .O(N__25481),
            .I(N__25404));
    InMux I__5965 (
            .O(N__25478),
            .I(N__25404));
    InMux I__5964 (
            .O(N__25477),
            .I(N__25404));
    InMux I__5963 (
            .O(N__25474),
            .I(N__25401));
    InMux I__5962 (
            .O(N__25473),
            .I(N__25398));
    LocalMux I__5961 (
            .O(N__25468),
            .I(N__25391));
    LocalMux I__5960 (
            .O(N__25461),
            .I(N__25391));
    LocalMux I__5959 (
            .O(N__25454),
            .I(N__25391));
    LocalMux I__5958 (
            .O(N__25451),
            .I(N__25386));
    LocalMux I__5957 (
            .O(N__25448),
            .I(N__25386));
    LocalMux I__5956 (
            .O(N__25443),
            .I(N__25381));
    LocalMux I__5955 (
            .O(N__25438),
            .I(N__25381));
    Span4Mux_v I__5954 (
            .O(N__25435),
            .I(N__25378));
    InMux I__5953 (
            .O(N__25434),
            .I(N__25362));
    InMux I__5952 (
            .O(N__25431),
            .I(N__25362));
    InMux I__5951 (
            .O(N__25430),
            .I(N__25362));
    InMux I__5950 (
            .O(N__25429),
            .I(N__25362));
    InMux I__5949 (
            .O(N__25426),
            .I(N__25362));
    InMux I__5948 (
            .O(N__25425),
            .I(N__25362));
    InMux I__5947 (
            .O(N__25424),
            .I(N__25362));
    InMux I__5946 (
            .O(N__25421),
            .I(N__25359));
    Span4Mux_h I__5945 (
            .O(N__25418),
            .I(N__25346));
    Span4Mux_h I__5944 (
            .O(N__25411),
            .I(N__25346));
    LocalMux I__5943 (
            .O(N__25404),
            .I(N__25346));
    LocalMux I__5942 (
            .O(N__25401),
            .I(N__25346));
    LocalMux I__5941 (
            .O(N__25398),
            .I(N__25346));
    Span4Mux_v I__5940 (
            .O(N__25391),
            .I(N__25346));
    Span4Mux_h I__5939 (
            .O(N__25386),
            .I(N__25343));
    Span4Mux_v I__5938 (
            .O(N__25381),
            .I(N__25338));
    Span4Mux_v I__5937 (
            .O(N__25378),
            .I(N__25338));
    InMux I__5936 (
            .O(N__25377),
            .I(N__25335));
    LocalMux I__5935 (
            .O(N__25362),
            .I(scaler_1_dv));
    LocalMux I__5934 (
            .O(N__25359),
            .I(scaler_1_dv));
    Odrv4 I__5933 (
            .O(N__25346),
            .I(scaler_1_dv));
    Odrv4 I__5932 (
            .O(N__25343),
            .I(scaler_1_dv));
    Odrv4 I__5931 (
            .O(N__25338),
            .I(scaler_1_dv));
    LocalMux I__5930 (
            .O(N__25335),
            .I(scaler_1_dv));
    InMux I__5929 (
            .O(N__25322),
            .I(N__25315));
    InMux I__5928 (
            .O(N__25321),
            .I(N__25315));
    InMux I__5927 (
            .O(N__25320),
            .I(N__25312));
    LocalMux I__5926 (
            .O(N__25315),
            .I(N__25309));
    LocalMux I__5925 (
            .O(N__25312),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    Odrv12 I__5924 (
            .O(N__25309),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    ClkMux I__5923 (
            .O(N__25304),
            .I(N__24938));
    ClkMux I__5922 (
            .O(N__25303),
            .I(N__24938));
    ClkMux I__5921 (
            .O(N__25302),
            .I(N__24938));
    ClkMux I__5920 (
            .O(N__25301),
            .I(N__24938));
    ClkMux I__5919 (
            .O(N__25300),
            .I(N__24938));
    ClkMux I__5918 (
            .O(N__25299),
            .I(N__24938));
    ClkMux I__5917 (
            .O(N__25298),
            .I(N__24938));
    ClkMux I__5916 (
            .O(N__25297),
            .I(N__24938));
    ClkMux I__5915 (
            .O(N__25296),
            .I(N__24938));
    ClkMux I__5914 (
            .O(N__25295),
            .I(N__24938));
    ClkMux I__5913 (
            .O(N__25294),
            .I(N__24938));
    ClkMux I__5912 (
            .O(N__25293),
            .I(N__24938));
    ClkMux I__5911 (
            .O(N__25292),
            .I(N__24938));
    ClkMux I__5910 (
            .O(N__25291),
            .I(N__24938));
    ClkMux I__5909 (
            .O(N__25290),
            .I(N__24938));
    ClkMux I__5908 (
            .O(N__25289),
            .I(N__24938));
    ClkMux I__5907 (
            .O(N__25288),
            .I(N__24938));
    ClkMux I__5906 (
            .O(N__25287),
            .I(N__24938));
    ClkMux I__5905 (
            .O(N__25286),
            .I(N__24938));
    ClkMux I__5904 (
            .O(N__25285),
            .I(N__24938));
    ClkMux I__5903 (
            .O(N__25284),
            .I(N__24938));
    ClkMux I__5902 (
            .O(N__25283),
            .I(N__24938));
    ClkMux I__5901 (
            .O(N__25282),
            .I(N__24938));
    ClkMux I__5900 (
            .O(N__25281),
            .I(N__24938));
    ClkMux I__5899 (
            .O(N__25280),
            .I(N__24938));
    ClkMux I__5898 (
            .O(N__25279),
            .I(N__24938));
    ClkMux I__5897 (
            .O(N__25278),
            .I(N__24938));
    ClkMux I__5896 (
            .O(N__25277),
            .I(N__24938));
    ClkMux I__5895 (
            .O(N__25276),
            .I(N__24938));
    ClkMux I__5894 (
            .O(N__25275),
            .I(N__24938));
    ClkMux I__5893 (
            .O(N__25274),
            .I(N__24938));
    ClkMux I__5892 (
            .O(N__25273),
            .I(N__24938));
    ClkMux I__5891 (
            .O(N__25272),
            .I(N__24938));
    ClkMux I__5890 (
            .O(N__25271),
            .I(N__24938));
    ClkMux I__5889 (
            .O(N__25270),
            .I(N__24938));
    ClkMux I__5888 (
            .O(N__25269),
            .I(N__24938));
    ClkMux I__5887 (
            .O(N__25268),
            .I(N__24938));
    ClkMux I__5886 (
            .O(N__25267),
            .I(N__24938));
    ClkMux I__5885 (
            .O(N__25266),
            .I(N__24938));
    ClkMux I__5884 (
            .O(N__25265),
            .I(N__24938));
    ClkMux I__5883 (
            .O(N__25264),
            .I(N__24938));
    ClkMux I__5882 (
            .O(N__25263),
            .I(N__24938));
    ClkMux I__5881 (
            .O(N__25262),
            .I(N__24938));
    ClkMux I__5880 (
            .O(N__25261),
            .I(N__24938));
    ClkMux I__5879 (
            .O(N__25260),
            .I(N__24938));
    ClkMux I__5878 (
            .O(N__25259),
            .I(N__24938));
    ClkMux I__5877 (
            .O(N__25258),
            .I(N__24938));
    ClkMux I__5876 (
            .O(N__25257),
            .I(N__24938));
    ClkMux I__5875 (
            .O(N__25256),
            .I(N__24938));
    ClkMux I__5874 (
            .O(N__25255),
            .I(N__24938));
    ClkMux I__5873 (
            .O(N__25254),
            .I(N__24938));
    ClkMux I__5872 (
            .O(N__25253),
            .I(N__24938));
    ClkMux I__5871 (
            .O(N__25252),
            .I(N__24938));
    ClkMux I__5870 (
            .O(N__25251),
            .I(N__24938));
    ClkMux I__5869 (
            .O(N__25250),
            .I(N__24938));
    ClkMux I__5868 (
            .O(N__25249),
            .I(N__24938));
    ClkMux I__5867 (
            .O(N__25248),
            .I(N__24938));
    ClkMux I__5866 (
            .O(N__25247),
            .I(N__24938));
    ClkMux I__5865 (
            .O(N__25246),
            .I(N__24938));
    ClkMux I__5864 (
            .O(N__25245),
            .I(N__24938));
    ClkMux I__5863 (
            .O(N__25244),
            .I(N__24938));
    ClkMux I__5862 (
            .O(N__25243),
            .I(N__24938));
    ClkMux I__5861 (
            .O(N__25242),
            .I(N__24938));
    ClkMux I__5860 (
            .O(N__25241),
            .I(N__24938));
    ClkMux I__5859 (
            .O(N__25240),
            .I(N__24938));
    ClkMux I__5858 (
            .O(N__25239),
            .I(N__24938));
    ClkMux I__5857 (
            .O(N__25238),
            .I(N__24938));
    ClkMux I__5856 (
            .O(N__25237),
            .I(N__24938));
    ClkMux I__5855 (
            .O(N__25236),
            .I(N__24938));
    ClkMux I__5854 (
            .O(N__25235),
            .I(N__24938));
    ClkMux I__5853 (
            .O(N__25234),
            .I(N__24938));
    ClkMux I__5852 (
            .O(N__25233),
            .I(N__24938));
    ClkMux I__5851 (
            .O(N__25232),
            .I(N__24938));
    ClkMux I__5850 (
            .O(N__25231),
            .I(N__24938));
    ClkMux I__5849 (
            .O(N__25230),
            .I(N__24938));
    ClkMux I__5848 (
            .O(N__25229),
            .I(N__24938));
    ClkMux I__5847 (
            .O(N__25228),
            .I(N__24938));
    ClkMux I__5846 (
            .O(N__25227),
            .I(N__24938));
    ClkMux I__5845 (
            .O(N__25226),
            .I(N__24938));
    ClkMux I__5844 (
            .O(N__25225),
            .I(N__24938));
    ClkMux I__5843 (
            .O(N__25224),
            .I(N__24938));
    ClkMux I__5842 (
            .O(N__25223),
            .I(N__24938));
    ClkMux I__5841 (
            .O(N__25222),
            .I(N__24938));
    ClkMux I__5840 (
            .O(N__25221),
            .I(N__24938));
    ClkMux I__5839 (
            .O(N__25220),
            .I(N__24938));
    ClkMux I__5838 (
            .O(N__25219),
            .I(N__24938));
    ClkMux I__5837 (
            .O(N__25218),
            .I(N__24938));
    ClkMux I__5836 (
            .O(N__25217),
            .I(N__24938));
    ClkMux I__5835 (
            .O(N__25216),
            .I(N__24938));
    ClkMux I__5834 (
            .O(N__25215),
            .I(N__24938));
    ClkMux I__5833 (
            .O(N__25214),
            .I(N__24938));
    ClkMux I__5832 (
            .O(N__25213),
            .I(N__24938));
    ClkMux I__5831 (
            .O(N__25212),
            .I(N__24938));
    ClkMux I__5830 (
            .O(N__25211),
            .I(N__24938));
    ClkMux I__5829 (
            .O(N__25210),
            .I(N__24938));
    ClkMux I__5828 (
            .O(N__25209),
            .I(N__24938));
    ClkMux I__5827 (
            .O(N__25208),
            .I(N__24938));
    ClkMux I__5826 (
            .O(N__25207),
            .I(N__24938));
    ClkMux I__5825 (
            .O(N__25206),
            .I(N__24938));
    ClkMux I__5824 (
            .O(N__25205),
            .I(N__24938));
    ClkMux I__5823 (
            .O(N__25204),
            .I(N__24938));
    ClkMux I__5822 (
            .O(N__25203),
            .I(N__24938));
    ClkMux I__5821 (
            .O(N__25202),
            .I(N__24938));
    ClkMux I__5820 (
            .O(N__25201),
            .I(N__24938));
    ClkMux I__5819 (
            .O(N__25200),
            .I(N__24938));
    ClkMux I__5818 (
            .O(N__25199),
            .I(N__24938));
    ClkMux I__5817 (
            .O(N__25198),
            .I(N__24938));
    ClkMux I__5816 (
            .O(N__25197),
            .I(N__24938));
    ClkMux I__5815 (
            .O(N__25196),
            .I(N__24938));
    ClkMux I__5814 (
            .O(N__25195),
            .I(N__24938));
    ClkMux I__5813 (
            .O(N__25194),
            .I(N__24938));
    ClkMux I__5812 (
            .O(N__25193),
            .I(N__24938));
    ClkMux I__5811 (
            .O(N__25192),
            .I(N__24938));
    ClkMux I__5810 (
            .O(N__25191),
            .I(N__24938));
    ClkMux I__5809 (
            .O(N__25190),
            .I(N__24938));
    ClkMux I__5808 (
            .O(N__25189),
            .I(N__24938));
    ClkMux I__5807 (
            .O(N__25188),
            .I(N__24938));
    ClkMux I__5806 (
            .O(N__25187),
            .I(N__24938));
    ClkMux I__5805 (
            .O(N__25186),
            .I(N__24938));
    ClkMux I__5804 (
            .O(N__25185),
            .I(N__24938));
    ClkMux I__5803 (
            .O(N__25184),
            .I(N__24938));
    ClkMux I__5802 (
            .O(N__25183),
            .I(N__24938));
    GlobalMux I__5801 (
            .O(N__24938),
            .I(N__24935));
    gio2CtrlBuf I__5800 (
            .O(N__24935),
            .I(clk_system_c_g));
    CascadeMux I__5799 (
            .O(N__24932),
            .I(N__24924));
    CascadeMux I__5798 (
            .O(N__24931),
            .I(N__24921));
    CascadeMux I__5797 (
            .O(N__24930),
            .I(N__24913));
    InMux I__5796 (
            .O(N__24929),
            .I(N__24892));
    InMux I__5795 (
            .O(N__24928),
            .I(N__24889));
    InMux I__5794 (
            .O(N__24927),
            .I(N__24886));
    InMux I__5793 (
            .O(N__24924),
            .I(N__24881));
    InMux I__5792 (
            .O(N__24921),
            .I(N__24881));
    InMux I__5791 (
            .O(N__24920),
            .I(N__24878));
    InMux I__5790 (
            .O(N__24919),
            .I(N__24875));
    InMux I__5789 (
            .O(N__24918),
            .I(N__24872));
    InMux I__5788 (
            .O(N__24917),
            .I(N__24869));
    InMux I__5787 (
            .O(N__24916),
            .I(N__24862));
    InMux I__5786 (
            .O(N__24913),
            .I(N__24862));
    InMux I__5785 (
            .O(N__24912),
            .I(N__24862));
    InMux I__5784 (
            .O(N__24911),
            .I(N__24859));
    InMux I__5783 (
            .O(N__24910),
            .I(N__24856));
    InMux I__5782 (
            .O(N__24909),
            .I(N__24853));
    InMux I__5781 (
            .O(N__24908),
            .I(N__24850));
    InMux I__5780 (
            .O(N__24907),
            .I(N__24847));
    InMux I__5779 (
            .O(N__24906),
            .I(N__24842));
    InMux I__5778 (
            .O(N__24905),
            .I(N__24842));
    InMux I__5777 (
            .O(N__24904),
            .I(N__24839));
    InMux I__5776 (
            .O(N__24903),
            .I(N__24836));
    InMux I__5775 (
            .O(N__24902),
            .I(N__24833));
    InMux I__5774 (
            .O(N__24901),
            .I(N__24830));
    InMux I__5773 (
            .O(N__24900),
            .I(N__24827));
    InMux I__5772 (
            .O(N__24899),
            .I(N__24824));
    InMux I__5771 (
            .O(N__24898),
            .I(N__24821));
    InMux I__5770 (
            .O(N__24897),
            .I(N__24816));
    InMux I__5769 (
            .O(N__24896),
            .I(N__24816));
    InMux I__5768 (
            .O(N__24895),
            .I(N__24813));
    LocalMux I__5767 (
            .O(N__24892),
            .I(N__24737));
    LocalMux I__5766 (
            .O(N__24889),
            .I(N__24734));
    LocalMux I__5765 (
            .O(N__24886),
            .I(N__24731));
    LocalMux I__5764 (
            .O(N__24881),
            .I(N__24728));
    LocalMux I__5763 (
            .O(N__24878),
            .I(N__24725));
    LocalMux I__5762 (
            .O(N__24875),
            .I(N__24722));
    LocalMux I__5761 (
            .O(N__24872),
            .I(N__24719));
    LocalMux I__5760 (
            .O(N__24869),
            .I(N__24716));
    LocalMux I__5759 (
            .O(N__24862),
            .I(N__24713));
    LocalMux I__5758 (
            .O(N__24859),
            .I(N__24710));
    LocalMux I__5757 (
            .O(N__24856),
            .I(N__24707));
    LocalMux I__5756 (
            .O(N__24853),
            .I(N__24704));
    LocalMux I__5755 (
            .O(N__24850),
            .I(N__24701));
    LocalMux I__5754 (
            .O(N__24847),
            .I(N__24698));
    LocalMux I__5753 (
            .O(N__24842),
            .I(N__24695));
    LocalMux I__5752 (
            .O(N__24839),
            .I(N__24692));
    LocalMux I__5751 (
            .O(N__24836),
            .I(N__24689));
    LocalMux I__5750 (
            .O(N__24833),
            .I(N__24686));
    LocalMux I__5749 (
            .O(N__24830),
            .I(N__24683));
    LocalMux I__5748 (
            .O(N__24827),
            .I(N__24680));
    LocalMux I__5747 (
            .O(N__24824),
            .I(N__24677));
    LocalMux I__5746 (
            .O(N__24821),
            .I(N__24674));
    LocalMux I__5745 (
            .O(N__24816),
            .I(N__24671));
    LocalMux I__5744 (
            .O(N__24813),
            .I(N__24668));
    SRMux I__5743 (
            .O(N__24812),
            .I(N__24473));
    SRMux I__5742 (
            .O(N__24811),
            .I(N__24473));
    SRMux I__5741 (
            .O(N__24810),
            .I(N__24473));
    SRMux I__5740 (
            .O(N__24809),
            .I(N__24473));
    SRMux I__5739 (
            .O(N__24808),
            .I(N__24473));
    SRMux I__5738 (
            .O(N__24807),
            .I(N__24473));
    SRMux I__5737 (
            .O(N__24806),
            .I(N__24473));
    SRMux I__5736 (
            .O(N__24805),
            .I(N__24473));
    SRMux I__5735 (
            .O(N__24804),
            .I(N__24473));
    SRMux I__5734 (
            .O(N__24803),
            .I(N__24473));
    SRMux I__5733 (
            .O(N__24802),
            .I(N__24473));
    SRMux I__5732 (
            .O(N__24801),
            .I(N__24473));
    SRMux I__5731 (
            .O(N__24800),
            .I(N__24473));
    SRMux I__5730 (
            .O(N__24799),
            .I(N__24473));
    SRMux I__5729 (
            .O(N__24798),
            .I(N__24473));
    SRMux I__5728 (
            .O(N__24797),
            .I(N__24473));
    SRMux I__5727 (
            .O(N__24796),
            .I(N__24473));
    SRMux I__5726 (
            .O(N__24795),
            .I(N__24473));
    SRMux I__5725 (
            .O(N__24794),
            .I(N__24473));
    SRMux I__5724 (
            .O(N__24793),
            .I(N__24473));
    SRMux I__5723 (
            .O(N__24792),
            .I(N__24473));
    SRMux I__5722 (
            .O(N__24791),
            .I(N__24473));
    SRMux I__5721 (
            .O(N__24790),
            .I(N__24473));
    SRMux I__5720 (
            .O(N__24789),
            .I(N__24473));
    SRMux I__5719 (
            .O(N__24788),
            .I(N__24473));
    SRMux I__5718 (
            .O(N__24787),
            .I(N__24473));
    SRMux I__5717 (
            .O(N__24786),
            .I(N__24473));
    SRMux I__5716 (
            .O(N__24785),
            .I(N__24473));
    SRMux I__5715 (
            .O(N__24784),
            .I(N__24473));
    SRMux I__5714 (
            .O(N__24783),
            .I(N__24473));
    SRMux I__5713 (
            .O(N__24782),
            .I(N__24473));
    SRMux I__5712 (
            .O(N__24781),
            .I(N__24473));
    SRMux I__5711 (
            .O(N__24780),
            .I(N__24473));
    SRMux I__5710 (
            .O(N__24779),
            .I(N__24473));
    SRMux I__5709 (
            .O(N__24778),
            .I(N__24473));
    SRMux I__5708 (
            .O(N__24777),
            .I(N__24473));
    SRMux I__5707 (
            .O(N__24776),
            .I(N__24473));
    SRMux I__5706 (
            .O(N__24775),
            .I(N__24473));
    SRMux I__5705 (
            .O(N__24774),
            .I(N__24473));
    SRMux I__5704 (
            .O(N__24773),
            .I(N__24473));
    SRMux I__5703 (
            .O(N__24772),
            .I(N__24473));
    SRMux I__5702 (
            .O(N__24771),
            .I(N__24473));
    SRMux I__5701 (
            .O(N__24770),
            .I(N__24473));
    SRMux I__5700 (
            .O(N__24769),
            .I(N__24473));
    SRMux I__5699 (
            .O(N__24768),
            .I(N__24473));
    SRMux I__5698 (
            .O(N__24767),
            .I(N__24473));
    SRMux I__5697 (
            .O(N__24766),
            .I(N__24473));
    SRMux I__5696 (
            .O(N__24765),
            .I(N__24473));
    SRMux I__5695 (
            .O(N__24764),
            .I(N__24473));
    SRMux I__5694 (
            .O(N__24763),
            .I(N__24473));
    SRMux I__5693 (
            .O(N__24762),
            .I(N__24473));
    SRMux I__5692 (
            .O(N__24761),
            .I(N__24473));
    SRMux I__5691 (
            .O(N__24760),
            .I(N__24473));
    SRMux I__5690 (
            .O(N__24759),
            .I(N__24473));
    SRMux I__5689 (
            .O(N__24758),
            .I(N__24473));
    SRMux I__5688 (
            .O(N__24757),
            .I(N__24473));
    SRMux I__5687 (
            .O(N__24756),
            .I(N__24473));
    SRMux I__5686 (
            .O(N__24755),
            .I(N__24473));
    SRMux I__5685 (
            .O(N__24754),
            .I(N__24473));
    SRMux I__5684 (
            .O(N__24753),
            .I(N__24473));
    SRMux I__5683 (
            .O(N__24752),
            .I(N__24473));
    SRMux I__5682 (
            .O(N__24751),
            .I(N__24473));
    SRMux I__5681 (
            .O(N__24750),
            .I(N__24473));
    SRMux I__5680 (
            .O(N__24749),
            .I(N__24473));
    SRMux I__5679 (
            .O(N__24748),
            .I(N__24473));
    SRMux I__5678 (
            .O(N__24747),
            .I(N__24473));
    SRMux I__5677 (
            .O(N__24746),
            .I(N__24473));
    SRMux I__5676 (
            .O(N__24745),
            .I(N__24473));
    SRMux I__5675 (
            .O(N__24744),
            .I(N__24473));
    SRMux I__5674 (
            .O(N__24743),
            .I(N__24473));
    SRMux I__5673 (
            .O(N__24742),
            .I(N__24473));
    SRMux I__5672 (
            .O(N__24741),
            .I(N__24473));
    SRMux I__5671 (
            .O(N__24740),
            .I(N__24473));
    Glb2LocalMux I__5670 (
            .O(N__24737),
            .I(N__24473));
    Glb2LocalMux I__5669 (
            .O(N__24734),
            .I(N__24473));
    Glb2LocalMux I__5668 (
            .O(N__24731),
            .I(N__24473));
    Glb2LocalMux I__5667 (
            .O(N__24728),
            .I(N__24473));
    Glb2LocalMux I__5666 (
            .O(N__24725),
            .I(N__24473));
    Glb2LocalMux I__5665 (
            .O(N__24722),
            .I(N__24473));
    Glb2LocalMux I__5664 (
            .O(N__24719),
            .I(N__24473));
    Glb2LocalMux I__5663 (
            .O(N__24716),
            .I(N__24473));
    Glb2LocalMux I__5662 (
            .O(N__24713),
            .I(N__24473));
    Glb2LocalMux I__5661 (
            .O(N__24710),
            .I(N__24473));
    Glb2LocalMux I__5660 (
            .O(N__24707),
            .I(N__24473));
    Glb2LocalMux I__5659 (
            .O(N__24704),
            .I(N__24473));
    Glb2LocalMux I__5658 (
            .O(N__24701),
            .I(N__24473));
    Glb2LocalMux I__5657 (
            .O(N__24698),
            .I(N__24473));
    Glb2LocalMux I__5656 (
            .O(N__24695),
            .I(N__24473));
    Glb2LocalMux I__5655 (
            .O(N__24692),
            .I(N__24473));
    Glb2LocalMux I__5654 (
            .O(N__24689),
            .I(N__24473));
    Glb2LocalMux I__5653 (
            .O(N__24686),
            .I(N__24473));
    Glb2LocalMux I__5652 (
            .O(N__24683),
            .I(N__24473));
    Glb2LocalMux I__5651 (
            .O(N__24680),
            .I(N__24473));
    Glb2LocalMux I__5650 (
            .O(N__24677),
            .I(N__24473));
    Glb2LocalMux I__5649 (
            .O(N__24674),
            .I(N__24473));
    Glb2LocalMux I__5648 (
            .O(N__24671),
            .I(N__24473));
    Glb2LocalMux I__5647 (
            .O(N__24668),
            .I(N__24473));
    GlobalMux I__5646 (
            .O(N__24473),
            .I(N__24470));
    gio2CtrlBuf I__5645 (
            .O(N__24470),
            .I(reset_system_g));
    InMux I__5644 (
            .O(N__24467),
            .I(N__24464));
    LocalMux I__5643 (
            .O(N__24464),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ));
    InMux I__5642 (
            .O(N__24461),
            .I(N__24456));
    InMux I__5641 (
            .O(N__24460),
            .I(N__24453));
    InMux I__5640 (
            .O(N__24459),
            .I(N__24450));
    LocalMux I__5639 (
            .O(N__24456),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__5638 (
            .O(N__24453),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__5637 (
            .O(N__24450),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    CascadeMux I__5636 (
            .O(N__24443),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ));
    InMux I__5635 (
            .O(N__24440),
            .I(N__24435));
    InMux I__5634 (
            .O(N__24439),
            .I(N__24432));
    InMux I__5633 (
            .O(N__24438),
            .I(N__24429));
    LocalMux I__5632 (
            .O(N__24435),
            .I(N__24426));
    LocalMux I__5631 (
            .O(N__24432),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__5630 (
            .O(N__24429),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__5629 (
            .O(N__24426),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    CascadeMux I__5628 (
            .O(N__24419),
            .I(\ppm_encoder_1.N_148_17_cascade_ ));
    InMux I__5627 (
            .O(N__24416),
            .I(N__24413));
    LocalMux I__5626 (
            .O(N__24413),
            .I(N__24410));
    Odrv12 I__5625 (
            .O(N__24410),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    InMux I__5624 (
            .O(N__24407),
            .I(N__24401));
    InMux I__5623 (
            .O(N__24406),
            .I(N__24401));
    LocalMux I__5622 (
            .O(N__24401),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    InMux I__5621 (
            .O(N__24398),
            .I(N__24395));
    LocalMux I__5620 (
            .O(N__24395),
            .I(\ppm_encoder_1.N_148_17 ));
    CascadeMux I__5619 (
            .O(N__24392),
            .I(N__24389));
    InMux I__5618 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__5617 (
            .O(N__24386),
            .I(N__24383));
    Odrv4 I__5616 (
            .O(N__24383),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    InMux I__5615 (
            .O(N__24380),
            .I(N__24377));
    LocalMux I__5614 (
            .O(N__24377),
            .I(N__24374));
    Span12Mux_v I__5613 (
            .O(N__24374),
            .I(N__24371));
    Odrv12 I__5612 (
            .O(N__24371),
            .I(\ppm_encoder_1.N_148 ));
    InMux I__5611 (
            .O(N__24368),
            .I(N__24363));
    InMux I__5610 (
            .O(N__24367),
            .I(N__24360));
    InMux I__5609 (
            .O(N__24366),
            .I(N__24357));
    LocalMux I__5608 (
            .O(N__24363),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__5607 (
            .O(N__24360),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__5606 (
            .O(N__24357),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__5605 (
            .O(N__24350),
            .I(N__24345));
    InMux I__5604 (
            .O(N__24349),
            .I(N__24342));
    InMux I__5603 (
            .O(N__24348),
            .I(N__24339));
    LocalMux I__5602 (
            .O(N__24345),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__5601 (
            .O(N__24342),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__5600 (
            .O(N__24339),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    CascadeMux I__5599 (
            .O(N__24332),
            .I(N__24328));
    InMux I__5598 (
            .O(N__24331),
            .I(N__24324));
    InMux I__5597 (
            .O(N__24328),
            .I(N__24321));
    InMux I__5596 (
            .O(N__24327),
            .I(N__24318));
    LocalMux I__5595 (
            .O(N__24324),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__5594 (
            .O(N__24321),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__5593 (
            .O(N__24318),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__5592 (
            .O(N__24311),
            .I(N__24306));
    InMux I__5591 (
            .O(N__24310),
            .I(N__24303));
    InMux I__5590 (
            .O(N__24309),
            .I(N__24300));
    LocalMux I__5589 (
            .O(N__24306),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__5588 (
            .O(N__24303),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__5587 (
            .O(N__24300),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__5586 (
            .O(N__24293),
            .I(N__24287));
    InMux I__5585 (
            .O(N__24292),
            .I(N__24287));
    LocalMux I__5584 (
            .O(N__24287),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    CascadeMux I__5583 (
            .O(N__24284),
            .I(N__24281));
    InMux I__5582 (
            .O(N__24281),
            .I(N__24275));
    InMux I__5581 (
            .O(N__24280),
            .I(N__24275));
    LocalMux I__5580 (
            .O(N__24275),
            .I(N__24272));
    Span4Mux_h I__5579 (
            .O(N__24272),
            .I(N__24269));
    Span4Mux_v I__5578 (
            .O(N__24269),
            .I(N__24265));
    InMux I__5577 (
            .O(N__24268),
            .I(N__24262));
    Odrv4 I__5576 (
            .O(N__24265),
            .I(\ppm_encoder_1.N_241 ));
    LocalMux I__5575 (
            .O(N__24262),
            .I(\ppm_encoder_1.N_241 ));
    InMux I__5574 (
            .O(N__24257),
            .I(N__24253));
    InMux I__5573 (
            .O(N__24256),
            .I(N__24249));
    LocalMux I__5572 (
            .O(N__24253),
            .I(N__24246));
    InMux I__5571 (
            .O(N__24252),
            .I(N__24243));
    LocalMux I__5570 (
            .O(N__24249),
            .I(N__24240));
    Span4Mux_v I__5569 (
            .O(N__24246),
            .I(N__24236));
    LocalMux I__5568 (
            .O(N__24243),
            .I(N__24233));
    Span4Mux_v I__5567 (
            .O(N__24240),
            .I(N__24230));
    InMux I__5566 (
            .O(N__24239),
            .I(N__24227));
    Span4Mux_v I__5565 (
            .O(N__24236),
            .I(N__24222));
    Span4Mux_s2_v I__5564 (
            .O(N__24233),
            .I(N__24222));
    Odrv4 I__5563 (
            .O(N__24230),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__5562 (
            .O(N__24227),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__5561 (
            .O(N__24222),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__5560 (
            .O(N__24215),
            .I(N__24207));
    InMux I__5559 (
            .O(N__24214),
            .I(N__24204));
    IoInMux I__5558 (
            .O(N__24213),
            .I(N__24200));
    CascadeMux I__5557 (
            .O(N__24212),
            .I(N__24196));
    CascadeMux I__5556 (
            .O(N__24211),
            .I(N__24188));
    CascadeMux I__5555 (
            .O(N__24210),
            .I(N__24185));
    LocalMux I__5554 (
            .O(N__24207),
            .I(N__24181));
    LocalMux I__5553 (
            .O(N__24204),
            .I(N__24178));
    CascadeMux I__5552 (
            .O(N__24203),
            .I(N__24174));
    LocalMux I__5551 (
            .O(N__24200),
            .I(N__24170));
    CascadeMux I__5550 (
            .O(N__24199),
            .I(N__24165));
    InMux I__5549 (
            .O(N__24196),
            .I(N__24160));
    InMux I__5548 (
            .O(N__24195),
            .I(N__24160));
    InMux I__5547 (
            .O(N__24194),
            .I(N__24157));
    InMux I__5546 (
            .O(N__24193),
            .I(N__24154));
    InMux I__5545 (
            .O(N__24192),
            .I(N__24151));
    InMux I__5544 (
            .O(N__24191),
            .I(N__24148));
    InMux I__5543 (
            .O(N__24188),
            .I(N__24141));
    InMux I__5542 (
            .O(N__24185),
            .I(N__24141));
    InMux I__5541 (
            .O(N__24184),
            .I(N__24141));
    Span4Mux_v I__5540 (
            .O(N__24181),
            .I(N__24136));
    Span4Mux_v I__5539 (
            .O(N__24178),
            .I(N__24136));
    InMux I__5538 (
            .O(N__24177),
            .I(N__24133));
    InMux I__5537 (
            .O(N__24174),
            .I(N__24130));
    InMux I__5536 (
            .O(N__24173),
            .I(N__24127));
    IoSpan4Mux I__5535 (
            .O(N__24170),
            .I(N__24124));
    CascadeMux I__5534 (
            .O(N__24169),
            .I(N__24121));
    InMux I__5533 (
            .O(N__24168),
            .I(N__24111));
    InMux I__5532 (
            .O(N__24165),
            .I(N__24111));
    LocalMux I__5531 (
            .O(N__24160),
            .I(N__24106));
    LocalMux I__5530 (
            .O(N__24157),
            .I(N__24106));
    LocalMux I__5529 (
            .O(N__24154),
            .I(N__24101));
    LocalMux I__5528 (
            .O(N__24151),
            .I(N__24101));
    LocalMux I__5527 (
            .O(N__24148),
            .I(N__24098));
    LocalMux I__5526 (
            .O(N__24141),
            .I(N__24091));
    Sp12to4 I__5525 (
            .O(N__24136),
            .I(N__24091));
    LocalMux I__5524 (
            .O(N__24133),
            .I(N__24091));
    LocalMux I__5523 (
            .O(N__24130),
            .I(N__24088));
    LocalMux I__5522 (
            .O(N__24127),
            .I(N__24085));
    Sp12to4 I__5521 (
            .O(N__24124),
            .I(N__24082));
    InMux I__5520 (
            .O(N__24121),
            .I(N__24077));
    InMux I__5519 (
            .O(N__24120),
            .I(N__24077));
    InMux I__5518 (
            .O(N__24119),
            .I(N__24072));
    InMux I__5517 (
            .O(N__24118),
            .I(N__24072));
    InMux I__5516 (
            .O(N__24117),
            .I(N__24067));
    InMux I__5515 (
            .O(N__24116),
            .I(N__24067));
    LocalMux I__5514 (
            .O(N__24111),
            .I(N__24064));
    Span4Mux_h I__5513 (
            .O(N__24106),
            .I(N__24061));
    Span4Mux_h I__5512 (
            .O(N__24101),
            .I(N__24056));
    Span4Mux_s3_h I__5511 (
            .O(N__24098),
            .I(N__24056));
    Span12Mux_h I__5510 (
            .O(N__24091),
            .I(N__24051));
    Span12Mux_h I__5509 (
            .O(N__24088),
            .I(N__24051));
    Span12Mux_h I__5508 (
            .O(N__24085),
            .I(N__24046));
    Span12Mux_s9_v I__5507 (
            .O(N__24082),
            .I(N__24046));
    LocalMux I__5506 (
            .O(N__24077),
            .I(reset_system));
    LocalMux I__5505 (
            .O(N__24072),
            .I(reset_system));
    LocalMux I__5504 (
            .O(N__24067),
            .I(reset_system));
    Odrv4 I__5503 (
            .O(N__24064),
            .I(reset_system));
    Odrv4 I__5502 (
            .O(N__24061),
            .I(reset_system));
    Odrv4 I__5501 (
            .O(N__24056),
            .I(reset_system));
    Odrv12 I__5500 (
            .O(N__24051),
            .I(reset_system));
    Odrv12 I__5499 (
            .O(N__24046),
            .I(reset_system));
    InMux I__5498 (
            .O(N__24029),
            .I(N__24024));
    InMux I__5497 (
            .O(N__24028),
            .I(N__24020));
    CascadeMux I__5496 (
            .O(N__24027),
            .I(N__24016));
    LocalMux I__5495 (
            .O(N__24024),
            .I(N__24013));
    InMux I__5494 (
            .O(N__24023),
            .I(N__24010));
    LocalMux I__5493 (
            .O(N__24020),
            .I(N__24007));
    InMux I__5492 (
            .O(N__24019),
            .I(N__24002));
    InMux I__5491 (
            .O(N__24016),
            .I(N__24002));
    Span4Mux_v I__5490 (
            .O(N__24013),
            .I(N__23999));
    LocalMux I__5489 (
            .O(N__24010),
            .I(N__23996));
    Span4Mux_h I__5488 (
            .O(N__24007),
            .I(N__23991));
    LocalMux I__5487 (
            .O(N__24002),
            .I(N__23986));
    Span4Mux_h I__5486 (
            .O(N__23999),
            .I(N__23986));
    Span12Mux_s7_v I__5485 (
            .O(N__23996),
            .I(N__23983));
    InMux I__5484 (
            .O(N__23995),
            .I(N__23978));
    InMux I__5483 (
            .O(N__23994),
            .I(N__23978));
    Odrv4 I__5482 (
            .O(N__23991),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__5481 (
            .O(N__23986),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv12 I__5480 (
            .O(N__23983),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__5479 (
            .O(N__23978),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    IoInMux I__5478 (
            .O(N__23969),
            .I(N__23966));
    LocalMux I__5477 (
            .O(N__23966),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__5476 (
            .O(N__23963),
            .I(N__23960));
    LocalMux I__5475 (
            .O(N__23960),
            .I(N__23957));
    Span4Mux_h I__5474 (
            .O(N__23957),
            .I(N__23954));
    Span4Mux_h I__5473 (
            .O(N__23954),
            .I(N__23950));
    InMux I__5472 (
            .O(N__23953),
            .I(N__23947));
    Odrv4 I__5471 (
            .O(N__23950),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ));
    LocalMux I__5470 (
            .O(N__23947),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ));
    InMux I__5469 (
            .O(N__23942),
            .I(N__23939));
    LocalMux I__5468 (
            .O(N__23939),
            .I(N__23936));
    Span4Mux_h I__5467 (
            .O(N__23936),
            .I(N__23933));
    Span4Mux_h I__5466 (
            .O(N__23933),
            .I(N__23928));
    InMux I__5465 (
            .O(N__23932),
            .I(N__23925));
    InMux I__5464 (
            .O(N__23931),
            .I(N__23922));
    Odrv4 I__5463 (
            .O(N__23928),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ));
    LocalMux I__5462 (
            .O(N__23925),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ));
    LocalMux I__5461 (
            .O(N__23922),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ));
    InMux I__5460 (
            .O(N__23915),
            .I(N__23910));
    InMux I__5459 (
            .O(N__23914),
            .I(N__23905));
    InMux I__5458 (
            .O(N__23913),
            .I(N__23905));
    LocalMux I__5457 (
            .O(N__23910),
            .I(N__23895));
    LocalMux I__5456 (
            .O(N__23905),
            .I(N__23892));
    InMux I__5455 (
            .O(N__23904),
            .I(N__23889));
    InMux I__5454 (
            .O(N__23903),
            .I(N__23876));
    InMux I__5453 (
            .O(N__23902),
            .I(N__23876));
    InMux I__5452 (
            .O(N__23901),
            .I(N__23876));
    InMux I__5451 (
            .O(N__23900),
            .I(N__23876));
    InMux I__5450 (
            .O(N__23899),
            .I(N__23876));
    InMux I__5449 (
            .O(N__23898),
            .I(N__23876));
    Odrv12 I__5448 (
            .O(N__23895),
            .I(\uart_frame_decoder.N_85 ));
    Odrv4 I__5447 (
            .O(N__23892),
            .I(\uart_frame_decoder.N_85 ));
    LocalMux I__5446 (
            .O(N__23889),
            .I(\uart_frame_decoder.N_85 ));
    LocalMux I__5445 (
            .O(N__23876),
            .I(\uart_frame_decoder.N_85 ));
    CascadeMux I__5444 (
            .O(N__23867),
            .I(N__23863));
    InMux I__5443 (
            .O(N__23866),
            .I(N__23860));
    InMux I__5442 (
            .O(N__23863),
            .I(N__23857));
    LocalMux I__5441 (
            .O(N__23860),
            .I(N__23854));
    LocalMux I__5440 (
            .O(N__23857),
            .I(N__23849));
    Span4Mux_v I__5439 (
            .O(N__23854),
            .I(N__23849));
    Odrv4 I__5438 (
            .O(N__23849),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    InMux I__5437 (
            .O(N__23846),
            .I(N__23842));
    InMux I__5436 (
            .O(N__23845),
            .I(N__23839));
    LocalMux I__5435 (
            .O(N__23842),
            .I(N__23836));
    LocalMux I__5434 (
            .O(N__23839),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    Odrv12 I__5433 (
            .O(N__23836),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    CascadeMux I__5432 (
            .O(N__23831),
            .I(N__23828));
    InMux I__5431 (
            .O(N__23828),
            .I(N__23813));
    InMux I__5430 (
            .O(N__23827),
            .I(N__23808));
    InMux I__5429 (
            .O(N__23826),
            .I(N__23808));
    InMux I__5428 (
            .O(N__23825),
            .I(N__23801));
    InMux I__5427 (
            .O(N__23824),
            .I(N__23801));
    InMux I__5426 (
            .O(N__23823),
            .I(N__23801));
    InMux I__5425 (
            .O(N__23822),
            .I(N__23798));
    InMux I__5424 (
            .O(N__23821),
            .I(N__23793));
    InMux I__5423 (
            .O(N__23820),
            .I(N__23793));
    InMux I__5422 (
            .O(N__23819),
            .I(N__23789));
    CascadeMux I__5421 (
            .O(N__23818),
            .I(N__23784));
    InMux I__5420 (
            .O(N__23817),
            .I(N__23779));
    InMux I__5419 (
            .O(N__23816),
            .I(N__23779));
    LocalMux I__5418 (
            .O(N__23813),
            .I(N__23772));
    LocalMux I__5417 (
            .O(N__23808),
            .I(N__23772));
    LocalMux I__5416 (
            .O(N__23801),
            .I(N__23772));
    LocalMux I__5415 (
            .O(N__23798),
            .I(N__23769));
    LocalMux I__5414 (
            .O(N__23793),
            .I(N__23766));
    InMux I__5413 (
            .O(N__23792),
            .I(N__23763));
    LocalMux I__5412 (
            .O(N__23789),
            .I(N__23760));
    InMux I__5411 (
            .O(N__23788),
            .I(N__23757));
    CascadeMux I__5410 (
            .O(N__23787),
            .I(N__23754));
    InMux I__5409 (
            .O(N__23784),
            .I(N__23751));
    LocalMux I__5408 (
            .O(N__23779),
            .I(N__23744));
    Span4Mux_v I__5407 (
            .O(N__23772),
            .I(N__23744));
    Span4Mux_h I__5406 (
            .O(N__23769),
            .I(N__23744));
    Span4Mux_h I__5405 (
            .O(N__23766),
            .I(N__23739));
    LocalMux I__5404 (
            .O(N__23763),
            .I(N__23739));
    Span4Mux_v I__5403 (
            .O(N__23760),
            .I(N__23734));
    LocalMux I__5402 (
            .O(N__23757),
            .I(N__23734));
    InMux I__5401 (
            .O(N__23754),
            .I(N__23731));
    LocalMux I__5400 (
            .O(N__23751),
            .I(N__23726));
    Span4Mux_v I__5399 (
            .O(N__23744),
            .I(N__23726));
    Span4Mux_v I__5398 (
            .O(N__23739),
            .I(N__23721));
    Span4Mux_h I__5397 (
            .O(N__23734),
            .I(N__23721));
    LocalMux I__5396 (
            .O(N__23731),
            .I(uart_pc_data_rdy));
    Odrv4 I__5395 (
            .O(N__23726),
            .I(uart_pc_data_rdy));
    Odrv4 I__5394 (
            .O(N__23721),
            .I(uart_pc_data_rdy));
    CascadeMux I__5393 (
            .O(N__23714),
            .I(N__23702));
    CascadeMux I__5392 (
            .O(N__23713),
            .I(N__23695));
    InMux I__5391 (
            .O(N__23712),
            .I(N__23664));
    InMux I__5390 (
            .O(N__23711),
            .I(N__23664));
    InMux I__5389 (
            .O(N__23710),
            .I(N__23664));
    InMux I__5388 (
            .O(N__23709),
            .I(N__23664));
    InMux I__5387 (
            .O(N__23708),
            .I(N__23664));
    InMux I__5386 (
            .O(N__23707),
            .I(N__23657));
    InMux I__5385 (
            .O(N__23706),
            .I(N__23657));
    InMux I__5384 (
            .O(N__23705),
            .I(N__23657));
    InMux I__5383 (
            .O(N__23702),
            .I(N__23644));
    InMux I__5382 (
            .O(N__23701),
            .I(N__23644));
    InMux I__5381 (
            .O(N__23700),
            .I(N__23644));
    InMux I__5380 (
            .O(N__23699),
            .I(N__23644));
    InMux I__5379 (
            .O(N__23698),
            .I(N__23641));
    InMux I__5378 (
            .O(N__23695),
            .I(N__23638));
    InMux I__5377 (
            .O(N__23694),
            .I(N__23635));
    CascadeMux I__5376 (
            .O(N__23693),
            .I(N__23632));
    InMux I__5375 (
            .O(N__23692),
            .I(N__23618));
    InMux I__5374 (
            .O(N__23691),
            .I(N__23618));
    InMux I__5373 (
            .O(N__23690),
            .I(N__23618));
    InMux I__5372 (
            .O(N__23689),
            .I(N__23618));
    InMux I__5371 (
            .O(N__23688),
            .I(N__23607));
    InMux I__5370 (
            .O(N__23687),
            .I(N__23607));
    InMux I__5369 (
            .O(N__23686),
            .I(N__23607));
    InMux I__5368 (
            .O(N__23685),
            .I(N__23607));
    InMux I__5367 (
            .O(N__23684),
            .I(N__23607));
    InMux I__5366 (
            .O(N__23683),
            .I(N__23602));
    InMux I__5365 (
            .O(N__23682),
            .I(N__23602));
    InMux I__5364 (
            .O(N__23681),
            .I(N__23595));
    InMux I__5363 (
            .O(N__23680),
            .I(N__23595));
    InMux I__5362 (
            .O(N__23679),
            .I(N__23595));
    CascadeMux I__5361 (
            .O(N__23678),
            .I(N__23585));
    CascadeMux I__5360 (
            .O(N__23677),
            .I(N__23582));
    CascadeMux I__5359 (
            .O(N__23676),
            .I(N__23579));
    InMux I__5358 (
            .O(N__23675),
            .I(N__23576));
    LocalMux I__5357 (
            .O(N__23664),
            .I(N__23573));
    LocalMux I__5356 (
            .O(N__23657),
            .I(N__23569));
    InMux I__5355 (
            .O(N__23656),
            .I(N__23560));
    InMux I__5354 (
            .O(N__23655),
            .I(N__23560));
    InMux I__5353 (
            .O(N__23654),
            .I(N__23560));
    InMux I__5352 (
            .O(N__23653),
            .I(N__23560));
    LocalMux I__5351 (
            .O(N__23644),
            .I(N__23557));
    LocalMux I__5350 (
            .O(N__23641),
            .I(N__23550));
    LocalMux I__5349 (
            .O(N__23638),
            .I(N__23545));
    LocalMux I__5348 (
            .O(N__23635),
            .I(N__23545));
    InMux I__5347 (
            .O(N__23632),
            .I(N__23540));
    InMux I__5346 (
            .O(N__23631),
            .I(N__23540));
    InMux I__5345 (
            .O(N__23630),
            .I(N__23531));
    InMux I__5344 (
            .O(N__23629),
            .I(N__23531));
    InMux I__5343 (
            .O(N__23628),
            .I(N__23531));
    InMux I__5342 (
            .O(N__23627),
            .I(N__23531));
    LocalMux I__5341 (
            .O(N__23618),
            .I(N__23522));
    LocalMux I__5340 (
            .O(N__23607),
            .I(N__23522));
    LocalMux I__5339 (
            .O(N__23602),
            .I(N__23522));
    LocalMux I__5338 (
            .O(N__23595),
            .I(N__23522));
    InMux I__5337 (
            .O(N__23594),
            .I(N__23513));
    InMux I__5336 (
            .O(N__23593),
            .I(N__23513));
    InMux I__5335 (
            .O(N__23592),
            .I(N__23513));
    InMux I__5334 (
            .O(N__23591),
            .I(N__23513));
    CascadeMux I__5333 (
            .O(N__23590),
            .I(N__23500));
    InMux I__5332 (
            .O(N__23589),
            .I(N__23496));
    InMux I__5331 (
            .O(N__23588),
            .I(N__23493));
    InMux I__5330 (
            .O(N__23585),
            .I(N__23486));
    InMux I__5329 (
            .O(N__23582),
            .I(N__23486));
    InMux I__5328 (
            .O(N__23579),
            .I(N__23486));
    LocalMux I__5327 (
            .O(N__23576),
            .I(N__23481));
    Span4Mux_v I__5326 (
            .O(N__23573),
            .I(N__23481));
    InMux I__5325 (
            .O(N__23572),
            .I(N__23478));
    Span4Mux_v I__5324 (
            .O(N__23569),
            .I(N__23471));
    LocalMux I__5323 (
            .O(N__23560),
            .I(N__23471));
    Span4Mux_h I__5322 (
            .O(N__23557),
            .I(N__23471));
    InMux I__5321 (
            .O(N__23556),
            .I(N__23462));
    InMux I__5320 (
            .O(N__23555),
            .I(N__23462));
    InMux I__5319 (
            .O(N__23554),
            .I(N__23462));
    InMux I__5318 (
            .O(N__23553),
            .I(N__23462));
    Span4Mux_v I__5317 (
            .O(N__23550),
            .I(N__23455));
    Span4Mux_v I__5316 (
            .O(N__23545),
            .I(N__23455));
    LocalMux I__5315 (
            .O(N__23540),
            .I(N__23455));
    LocalMux I__5314 (
            .O(N__23531),
            .I(N__23448));
    Span4Mux_v I__5313 (
            .O(N__23522),
            .I(N__23448));
    LocalMux I__5312 (
            .O(N__23513),
            .I(N__23448));
    InMux I__5311 (
            .O(N__23512),
            .I(N__23443));
    InMux I__5310 (
            .O(N__23511),
            .I(N__23443));
    InMux I__5309 (
            .O(N__23510),
            .I(N__23430));
    InMux I__5308 (
            .O(N__23509),
            .I(N__23430));
    InMux I__5307 (
            .O(N__23508),
            .I(N__23430));
    InMux I__5306 (
            .O(N__23507),
            .I(N__23430));
    InMux I__5305 (
            .O(N__23506),
            .I(N__23430));
    InMux I__5304 (
            .O(N__23505),
            .I(N__23430));
    InMux I__5303 (
            .O(N__23504),
            .I(N__23421));
    InMux I__5302 (
            .O(N__23503),
            .I(N__23421));
    InMux I__5301 (
            .O(N__23500),
            .I(N__23421));
    InMux I__5300 (
            .O(N__23499),
            .I(N__23421));
    LocalMux I__5299 (
            .O(N__23496),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5298 (
            .O(N__23493),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5297 (
            .O(N__23486),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    Odrv4 I__5296 (
            .O(N__23481),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5295 (
            .O(N__23478),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    Odrv4 I__5294 (
            .O(N__23471),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5293 (
            .O(N__23462),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    Odrv4 I__5292 (
            .O(N__23455),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    Odrv4 I__5291 (
            .O(N__23448),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5290 (
            .O(N__23443),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5289 (
            .O(N__23430),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    LocalMux I__5288 (
            .O(N__23421),
            .I(\ppm_encoder_1.PPM_STATE_62_d ));
    InMux I__5287 (
            .O(N__23396),
            .I(N__23393));
    LocalMux I__5286 (
            .O(N__23393),
            .I(N__23390));
    Span12Mux_s10_v I__5285 (
            .O(N__23390),
            .I(N__23387));
    Odrv12 I__5284 (
            .O(N__23387),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__5283 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__5282 (
            .O(N__23381),
            .I(N__23378));
    Span4Mux_v I__5281 (
            .O(N__23378),
            .I(N__23375));
    Odrv4 I__5280 (
            .O(N__23375),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    CascadeMux I__5279 (
            .O(N__23372),
            .I(N__23369));
    InMux I__5278 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__5277 (
            .O(N__23366),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__5276 (
            .O(N__23363),
            .I(N__23360));
    LocalMux I__5275 (
            .O(N__23360),
            .I(N__23357));
    Odrv4 I__5274 (
            .O(N__23357),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__5273 (
            .O(N__23354),
            .I(N__23351));
    LocalMux I__5272 (
            .O(N__23351),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__5271 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__5270 (
            .O(N__23345),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__5269 (
            .O(N__23342),
            .I(N__23339));
    LocalMux I__5268 (
            .O(N__23339),
            .I(N__23336));
    Span4Mux_v I__5267 (
            .O(N__23336),
            .I(N__23333));
    Span4Mux_v I__5266 (
            .O(N__23333),
            .I(N__23330));
    Sp12to4 I__5265 (
            .O(N__23330),
            .I(N__23327));
    Odrv12 I__5264 (
            .O(N__23327),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__5263 (
            .O(N__23324),
            .I(N__23321));
    LocalMux I__5262 (
            .O(N__23321),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    InMux I__5261 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__5260 (
            .O(N__23315),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    CascadeMux I__5259 (
            .O(N__23312),
            .I(N__23305));
    CascadeMux I__5258 (
            .O(N__23311),
            .I(N__23302));
    InMux I__5257 (
            .O(N__23310),
            .I(N__23296));
    InMux I__5256 (
            .O(N__23309),
            .I(N__23293));
    InMux I__5255 (
            .O(N__23308),
            .I(N__23290));
    InMux I__5254 (
            .O(N__23305),
            .I(N__23281));
    InMux I__5253 (
            .O(N__23302),
            .I(N__23281));
    InMux I__5252 (
            .O(N__23301),
            .I(N__23281));
    InMux I__5251 (
            .O(N__23300),
            .I(N__23281));
    CascadeMux I__5250 (
            .O(N__23299),
            .I(N__23278));
    LocalMux I__5249 (
            .O(N__23296),
            .I(N__23266));
    LocalMux I__5248 (
            .O(N__23293),
            .I(N__23266));
    LocalMux I__5247 (
            .O(N__23290),
            .I(N__23266));
    LocalMux I__5246 (
            .O(N__23281),
            .I(N__23266));
    InMux I__5245 (
            .O(N__23278),
            .I(N__23263));
    CascadeMux I__5244 (
            .O(N__23277),
            .I(N__23260));
    CascadeMux I__5243 (
            .O(N__23276),
            .I(N__23255));
    CascadeMux I__5242 (
            .O(N__23275),
            .I(N__23252));
    Span4Mux_v I__5241 (
            .O(N__23266),
            .I(N__23246));
    LocalMux I__5240 (
            .O(N__23263),
            .I(N__23246));
    InMux I__5239 (
            .O(N__23260),
            .I(N__23237));
    InMux I__5238 (
            .O(N__23259),
            .I(N__23237));
    InMux I__5237 (
            .O(N__23258),
            .I(N__23237));
    InMux I__5236 (
            .O(N__23255),
            .I(N__23237));
    InMux I__5235 (
            .O(N__23252),
            .I(N__23232));
    InMux I__5234 (
            .O(N__23251),
            .I(N__23232));
    Odrv4 I__5233 (
            .O(N__23246),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__5232 (
            .O(N__23237),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__5231 (
            .O(N__23232),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    InMux I__5230 (
            .O(N__23225),
            .I(N__23216));
    InMux I__5229 (
            .O(N__23224),
            .I(N__23213));
    InMux I__5228 (
            .O(N__23223),
            .I(N__23202));
    InMux I__5227 (
            .O(N__23222),
            .I(N__23193));
    InMux I__5226 (
            .O(N__23221),
            .I(N__23193));
    InMux I__5225 (
            .O(N__23220),
            .I(N__23193));
    InMux I__5224 (
            .O(N__23219),
            .I(N__23193));
    LocalMux I__5223 (
            .O(N__23216),
            .I(N__23187));
    LocalMux I__5222 (
            .O(N__23213),
            .I(N__23187));
    InMux I__5221 (
            .O(N__23212),
            .I(N__23184));
    InMux I__5220 (
            .O(N__23211),
            .I(N__23181));
    InMux I__5219 (
            .O(N__23210),
            .I(N__23172));
    InMux I__5218 (
            .O(N__23209),
            .I(N__23172));
    InMux I__5217 (
            .O(N__23208),
            .I(N__23172));
    InMux I__5216 (
            .O(N__23207),
            .I(N__23172));
    InMux I__5215 (
            .O(N__23206),
            .I(N__23167));
    InMux I__5214 (
            .O(N__23205),
            .I(N__23167));
    LocalMux I__5213 (
            .O(N__23202),
            .I(N__23161));
    LocalMux I__5212 (
            .O(N__23193),
            .I(N__23161));
    CascadeMux I__5211 (
            .O(N__23192),
            .I(N__23157));
    Span4Mux_v I__5210 (
            .O(N__23187),
            .I(N__23145));
    LocalMux I__5209 (
            .O(N__23184),
            .I(N__23145));
    LocalMux I__5208 (
            .O(N__23181),
            .I(N__23145));
    LocalMux I__5207 (
            .O(N__23172),
            .I(N__23145));
    LocalMux I__5206 (
            .O(N__23167),
            .I(N__23145));
    InMux I__5205 (
            .O(N__23166),
            .I(N__23142));
    Span4Mux_h I__5204 (
            .O(N__23161),
            .I(N__23139));
    InMux I__5203 (
            .O(N__23160),
            .I(N__23132));
    InMux I__5202 (
            .O(N__23157),
            .I(N__23132));
    InMux I__5201 (
            .O(N__23156),
            .I(N__23132));
    Span4Mux_v I__5200 (
            .O(N__23145),
            .I(N__23129));
    LocalMux I__5199 (
            .O(N__23142),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5198 (
            .O(N__23139),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__5197 (
            .O(N__23132),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__5196 (
            .O(N__23129),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    CascadeMux I__5195 (
            .O(N__23120),
            .I(N__23117));
    InMux I__5194 (
            .O(N__23117),
            .I(N__23113));
    CascadeMux I__5193 (
            .O(N__23116),
            .I(N__23110));
    LocalMux I__5192 (
            .O(N__23113),
            .I(N__23105));
    InMux I__5191 (
            .O(N__23110),
            .I(N__23098));
    InMux I__5190 (
            .O(N__23109),
            .I(N__23098));
    InMux I__5189 (
            .O(N__23108),
            .I(N__23098));
    Span4Mux_v I__5188 (
            .O(N__23105),
            .I(N__23093));
    LocalMux I__5187 (
            .O(N__23098),
            .I(N__23093));
    Odrv4 I__5186 (
            .O(N__23093),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    InMux I__5185 (
            .O(N__23090),
            .I(N__23087));
    LocalMux I__5184 (
            .O(N__23087),
            .I(N__23083));
    InMux I__5183 (
            .O(N__23086),
            .I(N__23080));
    Span4Mux_v I__5182 (
            .O(N__23083),
            .I(N__23076));
    LocalMux I__5181 (
            .O(N__23080),
            .I(N__23073));
    InMux I__5180 (
            .O(N__23079),
            .I(N__23070));
    Odrv4 I__5179 (
            .O(N__23076),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv4 I__5178 (
            .O(N__23073),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__5177 (
            .O(N__23070),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__5176 (
            .O(N__23063),
            .I(N__23060));
    LocalMux I__5175 (
            .O(N__23060),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    InMux I__5174 (
            .O(N__23057),
            .I(N__23052));
    InMux I__5173 (
            .O(N__23056),
            .I(N__23049));
    InMux I__5172 (
            .O(N__23055),
            .I(N__23046));
    LocalMux I__5171 (
            .O(N__23052),
            .I(N__23043));
    LocalMux I__5170 (
            .O(N__23049),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__5169 (
            .O(N__23046),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__5168 (
            .O(N__23043),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__5167 (
            .O(N__23036),
            .I(N__23031));
    InMux I__5166 (
            .O(N__23035),
            .I(N__23028));
    InMux I__5165 (
            .O(N__23034),
            .I(N__23025));
    LocalMux I__5164 (
            .O(N__23031),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__5163 (
            .O(N__23028),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__5162 (
            .O(N__23025),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    CascadeMux I__5161 (
            .O(N__23018),
            .I(N__23013));
    InMux I__5160 (
            .O(N__23017),
            .I(N__23010));
    InMux I__5159 (
            .O(N__23016),
            .I(N__23007));
    InMux I__5158 (
            .O(N__23013),
            .I(N__23004));
    LocalMux I__5157 (
            .O(N__23010),
            .I(N__23001));
    LocalMux I__5156 (
            .O(N__23007),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__5155 (
            .O(N__23004),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__5154 (
            .O(N__23001),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__5153 (
            .O(N__22994),
            .I(N__22989));
    InMux I__5152 (
            .O(N__22993),
            .I(N__22986));
    InMux I__5151 (
            .O(N__22992),
            .I(N__22983));
    LocalMux I__5150 (
            .O(N__22989),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__5149 (
            .O(N__22986),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__5148 (
            .O(N__22983),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__5147 (
            .O(N__22976),
            .I(N__22971));
    InMux I__5146 (
            .O(N__22975),
            .I(N__22968));
    InMux I__5145 (
            .O(N__22974),
            .I(N__22965));
    LocalMux I__5144 (
            .O(N__22971),
            .I(N__22962));
    LocalMux I__5143 (
            .O(N__22968),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__5142 (
            .O(N__22965),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__5141 (
            .O(N__22962),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__5140 (
            .O(N__22955),
            .I(N__22950));
    InMux I__5139 (
            .O(N__22954),
            .I(N__22947));
    InMux I__5138 (
            .O(N__22953),
            .I(N__22944));
    LocalMux I__5137 (
            .O(N__22950),
            .I(N__22941));
    LocalMux I__5136 (
            .O(N__22947),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__5135 (
            .O(N__22944),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__5134 (
            .O(N__22941),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    CascadeMux I__5133 (
            .O(N__22934),
            .I(N__22929));
    InMux I__5132 (
            .O(N__22933),
            .I(N__22926));
    InMux I__5131 (
            .O(N__22932),
            .I(N__22923));
    InMux I__5130 (
            .O(N__22929),
            .I(N__22920));
    LocalMux I__5129 (
            .O(N__22926),
            .I(N__22917));
    LocalMux I__5128 (
            .O(N__22923),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__5127 (
            .O(N__22920),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv4 I__5126 (
            .O(N__22917),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__5125 (
            .O(N__22910),
            .I(N__22907));
    LocalMux I__5124 (
            .O(N__22907),
            .I(N__22902));
    InMux I__5123 (
            .O(N__22906),
            .I(N__22899));
    InMux I__5122 (
            .O(N__22905),
            .I(N__22896));
    Span4Mux_h I__5121 (
            .O(N__22902),
            .I(N__22893));
    LocalMux I__5120 (
            .O(N__22899),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__5119 (
            .O(N__22896),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    Odrv4 I__5118 (
            .O(N__22893),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__5117 (
            .O(N__22886),
            .I(N__22883));
    LocalMux I__5116 (
            .O(N__22883),
            .I(N__22878));
    InMux I__5115 (
            .O(N__22882),
            .I(N__22875));
    InMux I__5114 (
            .O(N__22881),
            .I(N__22872));
    Span4Mux_h I__5113 (
            .O(N__22878),
            .I(N__22869));
    LocalMux I__5112 (
            .O(N__22875),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__5111 (
            .O(N__22872),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__5110 (
            .O(N__22869),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__5109 (
            .O(N__22862),
            .I(N__22857));
    InMux I__5108 (
            .O(N__22861),
            .I(N__22854));
    InMux I__5107 (
            .O(N__22860),
            .I(N__22851));
    LocalMux I__5106 (
            .O(N__22857),
            .I(N__22848));
    LocalMux I__5105 (
            .O(N__22854),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__5104 (
            .O(N__22851),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__5103 (
            .O(N__22848),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__5102 (
            .O(N__22841),
            .I(N__22834));
    CascadeMux I__5101 (
            .O(N__22840),
            .I(N__22831));
    CascadeMux I__5100 (
            .O(N__22839),
            .I(N__22828));
    CascadeMux I__5099 (
            .O(N__22838),
            .I(N__22816));
    InMux I__5098 (
            .O(N__22837),
            .I(N__22810));
    LocalMux I__5097 (
            .O(N__22834),
            .I(N__22807));
    InMux I__5096 (
            .O(N__22831),
            .I(N__22800));
    InMux I__5095 (
            .O(N__22828),
            .I(N__22800));
    InMux I__5094 (
            .O(N__22827),
            .I(N__22800));
    CascadeMux I__5093 (
            .O(N__22826),
            .I(N__22797));
    CascadeMux I__5092 (
            .O(N__22825),
            .I(N__22793));
    CascadeMux I__5091 (
            .O(N__22824),
            .I(N__22788));
    CascadeMux I__5090 (
            .O(N__22823),
            .I(N__22783));
    CascadeMux I__5089 (
            .O(N__22822),
            .I(N__22780));
    CascadeMux I__5088 (
            .O(N__22821),
            .I(N__22776));
    CascadeMux I__5087 (
            .O(N__22820),
            .I(N__22773));
    InMux I__5086 (
            .O(N__22819),
            .I(N__22761));
    InMux I__5085 (
            .O(N__22816),
            .I(N__22761));
    InMux I__5084 (
            .O(N__22815),
            .I(N__22761));
    InMux I__5083 (
            .O(N__22814),
            .I(N__22761));
    InMux I__5082 (
            .O(N__22813),
            .I(N__22756));
    LocalMux I__5081 (
            .O(N__22810),
            .I(N__22753));
    Span4Mux_v I__5080 (
            .O(N__22807),
            .I(N__22747));
    LocalMux I__5079 (
            .O(N__22800),
            .I(N__22744));
    InMux I__5078 (
            .O(N__22797),
            .I(N__22735));
    InMux I__5077 (
            .O(N__22796),
            .I(N__22735));
    InMux I__5076 (
            .O(N__22793),
            .I(N__22735));
    InMux I__5075 (
            .O(N__22792),
            .I(N__22735));
    InMux I__5074 (
            .O(N__22791),
            .I(N__22724));
    InMux I__5073 (
            .O(N__22788),
            .I(N__22724));
    InMux I__5072 (
            .O(N__22787),
            .I(N__22724));
    InMux I__5071 (
            .O(N__22786),
            .I(N__22724));
    InMux I__5070 (
            .O(N__22783),
            .I(N__22724));
    InMux I__5069 (
            .O(N__22780),
            .I(N__22719));
    InMux I__5068 (
            .O(N__22779),
            .I(N__22719));
    InMux I__5067 (
            .O(N__22776),
            .I(N__22712));
    InMux I__5066 (
            .O(N__22773),
            .I(N__22712));
    InMux I__5065 (
            .O(N__22772),
            .I(N__22712));
    CascadeMux I__5064 (
            .O(N__22771),
            .I(N__22709));
    CascadeMux I__5063 (
            .O(N__22770),
            .I(N__22706));
    LocalMux I__5062 (
            .O(N__22761),
            .I(N__22701));
    InMux I__5061 (
            .O(N__22760),
            .I(N__22696));
    InMux I__5060 (
            .O(N__22759),
            .I(N__22696));
    LocalMux I__5059 (
            .O(N__22756),
            .I(N__22688));
    Span4Mux_s3_v I__5058 (
            .O(N__22753),
            .I(N__22688));
    CascadeMux I__5057 (
            .O(N__22752),
            .I(N__22684));
    InMux I__5056 (
            .O(N__22751),
            .I(N__22678));
    InMux I__5055 (
            .O(N__22750),
            .I(N__22678));
    Span4Mux_h I__5054 (
            .O(N__22747),
            .I(N__22665));
    Span4Mux_s3_v I__5053 (
            .O(N__22744),
            .I(N__22665));
    LocalMux I__5052 (
            .O(N__22735),
            .I(N__22665));
    LocalMux I__5051 (
            .O(N__22724),
            .I(N__22665));
    LocalMux I__5050 (
            .O(N__22719),
            .I(N__22665));
    LocalMux I__5049 (
            .O(N__22712),
            .I(N__22665));
    InMux I__5048 (
            .O(N__22709),
            .I(N__22656));
    InMux I__5047 (
            .O(N__22706),
            .I(N__22656));
    InMux I__5046 (
            .O(N__22705),
            .I(N__22656));
    InMux I__5045 (
            .O(N__22704),
            .I(N__22656));
    Span4Mux_v I__5044 (
            .O(N__22701),
            .I(N__22651));
    LocalMux I__5043 (
            .O(N__22696),
            .I(N__22651));
    CascadeMux I__5042 (
            .O(N__22695),
            .I(N__22646));
    InMux I__5041 (
            .O(N__22694),
            .I(N__22643));
    InMux I__5040 (
            .O(N__22693),
            .I(N__22640));
    Span4Mux_v I__5039 (
            .O(N__22688),
            .I(N__22637));
    InMux I__5038 (
            .O(N__22687),
            .I(N__22634));
    InMux I__5037 (
            .O(N__22684),
            .I(N__22629));
    InMux I__5036 (
            .O(N__22683),
            .I(N__22629));
    LocalMux I__5035 (
            .O(N__22678),
            .I(N__22622));
    Span4Mux_v I__5034 (
            .O(N__22665),
            .I(N__22622));
    LocalMux I__5033 (
            .O(N__22656),
            .I(N__22622));
    Span4Mux_h I__5032 (
            .O(N__22651),
            .I(N__22619));
    InMux I__5031 (
            .O(N__22650),
            .I(N__22614));
    InMux I__5030 (
            .O(N__22649),
            .I(N__22614));
    InMux I__5029 (
            .O(N__22646),
            .I(N__22611));
    LocalMux I__5028 (
            .O(N__22643),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__5027 (
            .O(N__22640),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__5026 (
            .O(N__22637),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__5025 (
            .O(N__22634),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__5024 (
            .O(N__22629),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__5023 (
            .O(N__22622),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__5022 (
            .O(N__22619),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__5021 (
            .O(N__22614),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__5020 (
            .O(N__22611),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    InMux I__5019 (
            .O(N__22592),
            .I(N__22589));
    LocalMux I__5018 (
            .O(N__22589),
            .I(N__22586));
    Span4Mux_h I__5017 (
            .O(N__22586),
            .I(N__22583));
    Odrv4 I__5016 (
            .O(N__22583),
            .I(\ppm_encoder_1.N_301 ));
    InMux I__5015 (
            .O(N__22580),
            .I(N__22577));
    LocalMux I__5014 (
            .O(N__22577),
            .I(N__22574));
    Sp12to4 I__5013 (
            .O(N__22574),
            .I(N__22571));
    Span12Mux_s7_v I__5012 (
            .O(N__22571),
            .I(N__22566));
    InMux I__5011 (
            .O(N__22570),
            .I(N__22561));
    InMux I__5010 (
            .O(N__22569),
            .I(N__22561));
    Odrv12 I__5009 (
            .O(N__22566),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    LocalMux I__5008 (
            .O(N__22561),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__5007 (
            .O(N__22556),
            .I(N__22553));
    LocalMux I__5006 (
            .O(N__22553),
            .I(N__22550));
    Span4Mux_v I__5005 (
            .O(N__22550),
            .I(N__22545));
    InMux I__5004 (
            .O(N__22549),
            .I(N__22540));
    InMux I__5003 (
            .O(N__22548),
            .I(N__22540));
    Odrv4 I__5002 (
            .O(N__22545),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__5001 (
            .O(N__22540),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__5000 (
            .O(N__22535),
            .I(N__22532));
    LocalMux I__4999 (
            .O(N__22532),
            .I(N__22527));
    InMux I__4998 (
            .O(N__22531),
            .I(N__22524));
    InMux I__4997 (
            .O(N__22530),
            .I(N__22521));
    Span4Mux_v I__4996 (
            .O(N__22527),
            .I(N__22516));
    LocalMux I__4995 (
            .O(N__22524),
            .I(N__22516));
    LocalMux I__4994 (
            .O(N__22521),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__4993 (
            .O(N__22516),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    CascadeMux I__4992 (
            .O(N__22511),
            .I(N__22507));
    CascadeMux I__4991 (
            .O(N__22510),
            .I(N__22504));
    InMux I__4990 (
            .O(N__22507),
            .I(N__22499));
    InMux I__4989 (
            .O(N__22504),
            .I(N__22494));
    InMux I__4988 (
            .O(N__22503),
            .I(N__22494));
    InMux I__4987 (
            .O(N__22502),
            .I(N__22491));
    LocalMux I__4986 (
            .O(N__22499),
            .I(N__22486));
    LocalMux I__4985 (
            .O(N__22494),
            .I(N__22486));
    LocalMux I__4984 (
            .O(N__22491),
            .I(N__22483));
    Span4Mux_h I__4983 (
            .O(N__22486),
            .I(N__22480));
    Odrv4 I__4982 (
            .O(N__22483),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__4981 (
            .O(N__22480),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__4980 (
            .O(N__22475),
            .I(N__22472));
    LocalMux I__4979 (
            .O(N__22472),
            .I(N__22469));
    Span4Mux_h I__4978 (
            .O(N__22469),
            .I(N__22466));
    Odrv4 I__4977 (
            .O(N__22466),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    InMux I__4976 (
            .O(N__22463),
            .I(N__22460));
    LocalMux I__4975 (
            .O(N__22460),
            .I(N__22455));
    InMux I__4974 (
            .O(N__22459),
            .I(N__22450));
    InMux I__4973 (
            .O(N__22458),
            .I(N__22450));
    Odrv12 I__4972 (
            .O(N__22455),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    LocalMux I__4971 (
            .O(N__22450),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__4970 (
            .O(N__22445),
            .I(N__22440));
    InMux I__4969 (
            .O(N__22444),
            .I(N__22437));
    InMux I__4968 (
            .O(N__22443),
            .I(N__22434));
    LocalMux I__4967 (
            .O(N__22440),
            .I(N__22431));
    LocalMux I__4966 (
            .O(N__22437),
            .I(N__22428));
    LocalMux I__4965 (
            .O(N__22434),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv12 I__4964 (
            .O(N__22431),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__4963 (
            .O(N__22428),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__4962 (
            .O(N__22421),
            .I(\ppm_encoder_1.N_323_cascade_ ));
    InMux I__4961 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__4960 (
            .O(N__22415),
            .I(N__22410));
    InMux I__4959 (
            .O(N__22414),
            .I(N__22405));
    InMux I__4958 (
            .O(N__22413),
            .I(N__22405));
    Odrv12 I__4957 (
            .O(N__22410),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__4956 (
            .O(N__22405),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__4955 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__4954 (
            .O(N__22397),
            .I(N__22393));
    InMux I__4953 (
            .O(N__22396),
            .I(N__22390));
    Span4Mux_h I__4952 (
            .O(N__22393),
            .I(N__22384));
    LocalMux I__4951 (
            .O(N__22390),
            .I(N__22384));
    InMux I__4950 (
            .O(N__22389),
            .I(N__22381));
    Span4Mux_v I__4949 (
            .O(N__22384),
            .I(N__22378));
    LocalMux I__4948 (
            .O(N__22381),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__4947 (
            .O(N__22378),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__4946 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__4945 (
            .O(N__22370),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    InMux I__4944 (
            .O(N__22367),
            .I(N__22364));
    LocalMux I__4943 (
            .O(N__22364),
            .I(\ppm_encoder_1.N_322 ));
    InMux I__4942 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__4941 (
            .O(N__22358),
            .I(N__22355));
    Span4Mux_v I__4940 (
            .O(N__22355),
            .I(N__22352));
    Odrv4 I__4939 (
            .O(N__22352),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    InMux I__4938 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__4937 (
            .O(N__22346),
            .I(N__22341));
    InMux I__4936 (
            .O(N__22345),
            .I(N__22336));
    InMux I__4935 (
            .O(N__22344),
            .I(N__22336));
    Odrv12 I__4934 (
            .O(N__22341),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__4933 (
            .O(N__22336),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    InMux I__4932 (
            .O(N__22331),
            .I(N__22327));
    InMux I__4931 (
            .O(N__22330),
            .I(N__22324));
    LocalMux I__4930 (
            .O(N__22327),
            .I(N__22321));
    LocalMux I__4929 (
            .O(N__22324),
            .I(N__22318));
    Span4Mux_h I__4928 (
            .O(N__22321),
            .I(N__22314));
    Span4Mux_v I__4927 (
            .O(N__22318),
            .I(N__22311));
    InMux I__4926 (
            .O(N__22317),
            .I(N__22308));
    Odrv4 I__4925 (
            .O(N__22314),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__4924 (
            .O(N__22311),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    LocalMux I__4923 (
            .O(N__22308),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    CascadeMux I__4922 (
            .O(N__22301),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ));
    InMux I__4921 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__4920 (
            .O(N__22295),
            .I(N__22291));
    InMux I__4919 (
            .O(N__22294),
            .I(N__22288));
    Span4Mux_v I__4918 (
            .O(N__22291),
            .I(N__22285));
    LocalMux I__4917 (
            .O(N__22288),
            .I(N__22282));
    Odrv4 I__4916 (
            .O(N__22285),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv12 I__4915 (
            .O(N__22282),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__4914 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__4913 (
            .O(N__22274),
            .I(\ppm_encoder_1.N_309 ));
    InMux I__4912 (
            .O(N__22271),
            .I(N__22267));
    InMux I__4911 (
            .O(N__22270),
            .I(N__22264));
    LocalMux I__4910 (
            .O(N__22267),
            .I(N__22261));
    LocalMux I__4909 (
            .O(N__22264),
            .I(N__22258));
    Odrv4 I__4908 (
            .O(N__22261),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    Odrv4 I__4907 (
            .O(N__22258),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    InMux I__4906 (
            .O(N__22253),
            .I(N__22250));
    LocalMux I__4905 (
            .O(N__22250),
            .I(N__22246));
    InMux I__4904 (
            .O(N__22249),
            .I(N__22243));
    Span4Mux_v I__4903 (
            .O(N__22246),
            .I(N__22234));
    LocalMux I__4902 (
            .O(N__22243),
            .I(N__22234));
    InMux I__4901 (
            .O(N__22242),
            .I(N__22230));
    InMux I__4900 (
            .O(N__22241),
            .I(N__22227));
    InMux I__4899 (
            .O(N__22240),
            .I(N__22224));
    InMux I__4898 (
            .O(N__22239),
            .I(N__22221));
    Span4Mux_h I__4897 (
            .O(N__22234),
            .I(N__22218));
    InMux I__4896 (
            .O(N__22233),
            .I(N__22215));
    LocalMux I__4895 (
            .O(N__22230),
            .I(N__22210));
    LocalMux I__4894 (
            .O(N__22227),
            .I(N__22210));
    LocalMux I__4893 (
            .O(N__22224),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__4892 (
            .O(N__22221),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__4891 (
            .O(N__22218),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__4890 (
            .O(N__22215),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__4889 (
            .O(N__22210),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__4888 (
            .O(N__22199),
            .I(N__22196));
    LocalMux I__4887 (
            .O(N__22196),
            .I(N__22191));
    CascadeMux I__4886 (
            .O(N__22195),
            .I(N__22185));
    InMux I__4885 (
            .O(N__22194),
            .I(N__22182));
    Span4Mux_h I__4884 (
            .O(N__22191),
            .I(N__22179));
    CascadeMux I__4883 (
            .O(N__22190),
            .I(N__22176));
    InMux I__4882 (
            .O(N__22189),
            .I(N__22171));
    InMux I__4881 (
            .O(N__22188),
            .I(N__22171));
    InMux I__4880 (
            .O(N__22185),
            .I(N__22168));
    LocalMux I__4879 (
            .O(N__22182),
            .I(N__22165));
    Span4Mux_h I__4878 (
            .O(N__22179),
            .I(N__22162));
    InMux I__4877 (
            .O(N__22176),
            .I(N__22159));
    LocalMux I__4876 (
            .O(N__22171),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4875 (
            .O(N__22168),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv12 I__4874 (
            .O(N__22165),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__4873 (
            .O(N__22162),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__4872 (
            .O(N__22159),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__4871 (
            .O(N__22148),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ));
    InMux I__4870 (
            .O(N__22145),
            .I(N__22142));
    LocalMux I__4869 (
            .O(N__22142),
            .I(N__22139));
    Span4Mux_h I__4868 (
            .O(N__22139),
            .I(N__22133));
    InMux I__4867 (
            .O(N__22138),
            .I(N__22128));
    InMux I__4866 (
            .O(N__22137),
            .I(N__22128));
    InMux I__4865 (
            .O(N__22136),
            .I(N__22125));
    Odrv4 I__4864 (
            .O(N__22133),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__4863 (
            .O(N__22128),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__4862 (
            .O(N__22125),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    InMux I__4861 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__4860 (
            .O(N__22115),
            .I(N__22112));
    Span4Mux_h I__4859 (
            .O(N__22112),
            .I(N__22109));
    Span4Mux_v I__4858 (
            .O(N__22109),
            .I(N__22106));
    Odrv4 I__4857 (
            .O(N__22106),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    CascadeMux I__4856 (
            .O(N__22103),
            .I(N__22099));
    InMux I__4855 (
            .O(N__22102),
            .I(N__22095));
    InMux I__4854 (
            .O(N__22099),
            .I(N__22090));
    InMux I__4853 (
            .O(N__22098),
            .I(N__22090));
    LocalMux I__4852 (
            .O(N__22095),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    LocalMux I__4851 (
            .O(N__22090),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__4850 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__4849 (
            .O(N__22082),
            .I(N__22078));
    InMux I__4848 (
            .O(N__22081),
            .I(N__22075));
    Span4Mux_h I__4847 (
            .O(N__22078),
            .I(N__22070));
    LocalMux I__4846 (
            .O(N__22075),
            .I(N__22070));
    Span4Mux_h I__4845 (
            .O(N__22070),
            .I(N__22067));
    Odrv4 I__4844 (
            .O(N__22067),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__4843 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__4842 (
            .O(N__22061),
            .I(N__22058));
    Odrv4 I__4841 (
            .O(N__22058),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__4840 (
            .O(N__22055),
            .I(N__22051));
    InMux I__4839 (
            .O(N__22054),
            .I(N__22048));
    LocalMux I__4838 (
            .O(N__22051),
            .I(N__22043));
    LocalMux I__4837 (
            .O(N__22048),
            .I(N__22043));
    Span4Mux_h I__4836 (
            .O(N__22043),
            .I(N__22039));
    InMux I__4835 (
            .O(N__22042),
            .I(N__22036));
    Span4Mux_v I__4834 (
            .O(N__22039),
            .I(N__22033));
    LocalMux I__4833 (
            .O(N__22036),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__4832 (
            .O(N__22033),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__4831 (
            .O(N__22028),
            .I(N__22025));
    LocalMux I__4830 (
            .O(N__22025),
            .I(N__22021));
    InMux I__4829 (
            .O(N__22024),
            .I(N__22018));
    Span4Mux_h I__4828 (
            .O(N__22021),
            .I(N__22014));
    LocalMux I__4827 (
            .O(N__22018),
            .I(N__22011));
    InMux I__4826 (
            .O(N__22017),
            .I(N__22008));
    Odrv4 I__4825 (
            .O(N__22014),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv12 I__4824 (
            .O(N__22011),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    LocalMux I__4823 (
            .O(N__22008),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__4822 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__4821 (
            .O(N__21998),
            .I(N__21995));
    Span4Mux_s2_v I__4820 (
            .O(N__21995),
            .I(N__21992));
    Span4Mux_v I__4819 (
            .O(N__21992),
            .I(N__21989));
    Odrv4 I__4818 (
            .O(N__21989),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__4817 (
            .O(N__21986),
            .I(N__21982));
    InMux I__4816 (
            .O(N__21985),
            .I(N__21979));
    LocalMux I__4815 (
            .O(N__21982),
            .I(N__21976));
    LocalMux I__4814 (
            .O(N__21979),
            .I(N__21973));
    Span4Mux_v I__4813 (
            .O(N__21976),
            .I(N__21970));
    Odrv12 I__4812 (
            .O(N__21973),
            .I(scaler_1_data_13));
    Odrv4 I__4811 (
            .O(N__21970),
            .I(scaler_1_data_13));
    CascadeMux I__4810 (
            .O(N__21965),
            .I(N__21961));
    InMux I__4809 (
            .O(N__21964),
            .I(N__21956));
    InMux I__4808 (
            .O(N__21961),
            .I(N__21956));
    LocalMux I__4807 (
            .O(N__21956),
            .I(N__21945));
    CascadeMux I__4806 (
            .O(N__21955),
            .I(N__21942));
    CascadeMux I__4805 (
            .O(N__21954),
            .I(N__21939));
    CascadeMux I__4804 (
            .O(N__21953),
            .I(N__21936));
    CascadeMux I__4803 (
            .O(N__21952),
            .I(N__21933));
    CascadeMux I__4802 (
            .O(N__21951),
            .I(N__21930));
    CascadeMux I__4801 (
            .O(N__21950),
            .I(N__21927));
    CascadeMux I__4800 (
            .O(N__21949),
            .I(N__21924));
    CascadeMux I__4799 (
            .O(N__21948),
            .I(N__21917));
    Span4Mux_v I__4798 (
            .O(N__21945),
            .I(N__21913));
    InMux I__4797 (
            .O(N__21942),
            .I(N__21904));
    InMux I__4796 (
            .O(N__21939),
            .I(N__21904));
    InMux I__4795 (
            .O(N__21936),
            .I(N__21904));
    InMux I__4794 (
            .O(N__21933),
            .I(N__21904));
    InMux I__4793 (
            .O(N__21930),
            .I(N__21897));
    InMux I__4792 (
            .O(N__21927),
            .I(N__21897));
    InMux I__4791 (
            .O(N__21924),
            .I(N__21897));
    CascadeMux I__4790 (
            .O(N__21923),
            .I(N__21894));
    CascadeMux I__4789 (
            .O(N__21922),
            .I(N__21890));
    CascadeMux I__4788 (
            .O(N__21921),
            .I(N__21887));
    CascadeMux I__4787 (
            .O(N__21920),
            .I(N__21884));
    InMux I__4786 (
            .O(N__21917),
            .I(N__21881));
    CascadeMux I__4785 (
            .O(N__21916),
            .I(N__21878));
    Span4Mux_s1_v I__4784 (
            .O(N__21913),
            .I(N__21871));
    LocalMux I__4783 (
            .O(N__21904),
            .I(N__21871));
    LocalMux I__4782 (
            .O(N__21897),
            .I(N__21871));
    InMux I__4781 (
            .O(N__21894),
            .I(N__21868));
    InMux I__4780 (
            .O(N__21893),
            .I(N__21863));
    InMux I__4779 (
            .O(N__21890),
            .I(N__21863));
    InMux I__4778 (
            .O(N__21887),
            .I(N__21860));
    InMux I__4777 (
            .O(N__21884),
            .I(N__21857));
    LocalMux I__4776 (
            .O(N__21881),
            .I(N__21854));
    InMux I__4775 (
            .O(N__21878),
            .I(N__21851));
    Sp12to4 I__4774 (
            .O(N__21871),
            .I(N__21843));
    LocalMux I__4773 (
            .O(N__21868),
            .I(N__21843));
    LocalMux I__4772 (
            .O(N__21863),
            .I(N__21840));
    LocalMux I__4771 (
            .O(N__21860),
            .I(N__21835));
    LocalMux I__4770 (
            .O(N__21857),
            .I(N__21835));
    Span4Mux_h I__4769 (
            .O(N__21854),
            .I(N__21830));
    LocalMux I__4768 (
            .O(N__21851),
            .I(N__21830));
    CascadeMux I__4767 (
            .O(N__21850),
            .I(N__21827));
    InMux I__4766 (
            .O(N__21849),
            .I(N__21824));
    CascadeMux I__4765 (
            .O(N__21848),
            .I(N__21821));
    Span12Mux_s11_v I__4764 (
            .O(N__21843),
            .I(N__21818));
    Span4Mux_v I__4763 (
            .O(N__21840),
            .I(N__21815));
    Span4Mux_h I__4762 (
            .O(N__21835),
            .I(N__21810));
    Span4Mux_v I__4761 (
            .O(N__21830),
            .I(N__21810));
    InMux I__4760 (
            .O(N__21827),
            .I(N__21807));
    LocalMux I__4759 (
            .O(N__21824),
            .I(N__21804));
    InMux I__4758 (
            .O(N__21821),
            .I(N__21801));
    Odrv12 I__4757 (
            .O(N__21818),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4756 (
            .O(N__21815),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4755 (
            .O(N__21810),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4754 (
            .O(N__21807),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4753 (
            .O(N__21804),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4752 (
            .O(N__21801),
            .I(CONSTANT_ONE_NET));
    InMux I__4751 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__4750 (
            .O(N__21785),
            .I(N__21782));
    Span4Mux_v I__4749 (
            .O(N__21782),
            .I(N__21779));
    Span4Mux_v I__4748 (
            .O(N__21779),
            .I(N__21776));
    Odrv4 I__4747 (
            .O(N__21776),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__4746 (
            .O(N__21773),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__4745 (
            .O(N__21770),
            .I(N__21767));
    LocalMux I__4744 (
            .O(N__21767),
            .I(N__21764));
    Odrv4 I__4743 (
            .O(N__21764),
            .I(scaler_1_data_14));
    InMux I__4742 (
            .O(N__21761),
            .I(bfn_12_18_0_));
    InMux I__4741 (
            .O(N__21758),
            .I(N__21754));
    InMux I__4740 (
            .O(N__21757),
            .I(N__21751));
    LocalMux I__4739 (
            .O(N__21754),
            .I(N__21746));
    LocalMux I__4738 (
            .O(N__21751),
            .I(N__21746));
    Span4Mux_v I__4737 (
            .O(N__21746),
            .I(N__21743));
    Odrv4 I__4736 (
            .O(N__21743),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CEMux I__4735 (
            .O(N__21740),
            .I(N__21735));
    CEMux I__4734 (
            .O(N__21739),
            .I(N__21732));
    CEMux I__4733 (
            .O(N__21738),
            .I(N__21727));
    LocalMux I__4732 (
            .O(N__21735),
            .I(N__21723));
    LocalMux I__4731 (
            .O(N__21732),
            .I(N__21720));
    CEMux I__4730 (
            .O(N__21731),
            .I(N__21717));
    CEMux I__4729 (
            .O(N__21730),
            .I(N__21714));
    LocalMux I__4728 (
            .O(N__21727),
            .I(N__21711));
    CEMux I__4727 (
            .O(N__21726),
            .I(N__21708));
    Span4Mux_h I__4726 (
            .O(N__21723),
            .I(N__21700));
    Span4Mux_h I__4725 (
            .O(N__21720),
            .I(N__21700));
    LocalMux I__4724 (
            .O(N__21717),
            .I(N__21700));
    LocalMux I__4723 (
            .O(N__21714),
            .I(N__21697));
    Span4Mux_h I__4722 (
            .O(N__21711),
            .I(N__21694));
    LocalMux I__4721 (
            .O(N__21708),
            .I(N__21691));
    CEMux I__4720 (
            .O(N__21707),
            .I(N__21688));
    Sp12to4 I__4719 (
            .O(N__21700),
            .I(N__21685));
    Span4Mux_h I__4718 (
            .O(N__21697),
            .I(N__21680));
    Span4Mux_h I__4717 (
            .O(N__21694),
            .I(N__21680));
    Span4Mux_h I__4716 (
            .O(N__21691),
            .I(N__21675));
    LocalMux I__4715 (
            .O(N__21688),
            .I(N__21675));
    Odrv12 I__4714 (
            .O(N__21685),
            .I(\ppm_encoder_1.scaler_1_dv_0 ));
    Odrv4 I__4713 (
            .O(N__21680),
            .I(\ppm_encoder_1.scaler_1_dv_0 ));
    Odrv4 I__4712 (
            .O(N__21675),
            .I(\ppm_encoder_1.scaler_1_dv_0 ));
    InMux I__4711 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__4710 (
            .O(N__21665),
            .I(N__21662));
    Odrv4 I__4709 (
            .O(N__21662),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__4708 (
            .O(N__21659),
            .I(N__21656));
    LocalMux I__4707 (
            .O(N__21656),
            .I(N__21652));
    InMux I__4706 (
            .O(N__21655),
            .I(N__21649));
    Span4Mux_v I__4705 (
            .O(N__21652),
            .I(N__21644));
    LocalMux I__4704 (
            .O(N__21649),
            .I(N__21644));
    Odrv4 I__4703 (
            .O(N__21644),
            .I(scaler_1_data_8));
    InMux I__4702 (
            .O(N__21641),
            .I(N__21637));
    InMux I__4701 (
            .O(N__21640),
            .I(N__21634));
    LocalMux I__4700 (
            .O(N__21637),
            .I(N__21630));
    LocalMux I__4699 (
            .O(N__21634),
            .I(N__21627));
    InMux I__4698 (
            .O(N__21633),
            .I(N__21624));
    Span4Mux_h I__4697 (
            .O(N__21630),
            .I(N__21621));
    Span4Mux_v I__4696 (
            .O(N__21627),
            .I(N__21618));
    LocalMux I__4695 (
            .O(N__21624),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__4694 (
            .O(N__21621),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__4693 (
            .O(N__21618),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__4692 (
            .O(N__21611),
            .I(N__21608));
    LocalMux I__4691 (
            .O(N__21608),
            .I(N__21604));
    InMux I__4690 (
            .O(N__21607),
            .I(N__21601));
    Span4Mux_v I__4689 (
            .O(N__21604),
            .I(N__21596));
    LocalMux I__4688 (
            .O(N__21601),
            .I(N__21596));
    Span4Mux_v I__4687 (
            .O(N__21596),
            .I(N__21593));
    Odrv4 I__4686 (
            .O(N__21593),
            .I(scaler_4_data_11));
    InMux I__4685 (
            .O(N__21590),
            .I(N__21587));
    LocalMux I__4684 (
            .O(N__21587),
            .I(N__21584));
    Odrv4 I__4683 (
            .O(N__21584),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__4682 (
            .O(N__21581),
            .I(N__21578));
    LocalMux I__4681 (
            .O(N__21578),
            .I(N__21575));
    Odrv4 I__4680 (
            .O(N__21575),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__4679 (
            .O(N__21572),
            .I(N__21569));
    LocalMux I__4678 (
            .O(N__21569),
            .I(N__21565));
    InMux I__4677 (
            .O(N__21568),
            .I(N__21562));
    Span4Mux_h I__4676 (
            .O(N__21565),
            .I(N__21559));
    LocalMux I__4675 (
            .O(N__21562),
            .I(N__21556));
    Odrv4 I__4674 (
            .O(N__21559),
            .I(scaler_1_data_10));
    Odrv12 I__4673 (
            .O(N__21556),
            .I(scaler_1_data_10));
    InMux I__4672 (
            .O(N__21551),
            .I(N__21544));
    InMux I__4671 (
            .O(N__21550),
            .I(N__21544));
    CascadeMux I__4670 (
            .O(N__21549),
            .I(N__21541));
    LocalMux I__4669 (
            .O(N__21544),
            .I(N__21538));
    InMux I__4668 (
            .O(N__21541),
            .I(N__21535));
    Span4Mux_v I__4667 (
            .O(N__21538),
            .I(N__21532));
    LocalMux I__4666 (
            .O(N__21535),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__4665 (
            .O(N__21532),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__4664 (
            .O(N__21527),
            .I(N__21524));
    LocalMux I__4663 (
            .O(N__21524),
            .I(N__21520));
    InMux I__4662 (
            .O(N__21523),
            .I(N__21517));
    Span4Mux_v I__4661 (
            .O(N__21520),
            .I(N__21514));
    LocalMux I__4660 (
            .O(N__21517),
            .I(N__21511));
    Span4Mux_v I__4659 (
            .O(N__21514),
            .I(N__21506));
    Span4Mux_v I__4658 (
            .O(N__21511),
            .I(N__21506));
    Odrv4 I__4657 (
            .O(N__21506),
            .I(scaler_4_data_12));
    InMux I__4656 (
            .O(N__21503),
            .I(N__21500));
    LocalMux I__4655 (
            .O(N__21500),
            .I(N__21497));
    Span4Mux_v I__4654 (
            .O(N__21497),
            .I(N__21494));
    Odrv4 I__4653 (
            .O(N__21494),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__4652 (
            .O(N__21491),
            .I(N__21488));
    LocalMux I__4651 (
            .O(N__21488),
            .I(\ppm_encoder_1.N_143_0 ));
    CascadeMux I__4650 (
            .O(N__21485),
            .I(N__21482));
    InMux I__4649 (
            .O(N__21482),
            .I(N__21478));
    InMux I__4648 (
            .O(N__21481),
            .I(N__21475));
    LocalMux I__4647 (
            .O(N__21478),
            .I(N__21472));
    LocalMux I__4646 (
            .O(N__21475),
            .I(N__21469));
    Span4Mux_h I__4645 (
            .O(N__21472),
            .I(N__21464));
    Span4Mux_h I__4644 (
            .O(N__21469),
            .I(N__21461));
    CascadeMux I__4643 (
            .O(N__21468),
            .I(N__21458));
    InMux I__4642 (
            .O(N__21467),
            .I(N__21455));
    Span4Mux_h I__4641 (
            .O(N__21464),
            .I(N__21450));
    Span4Mux_v I__4640 (
            .O(N__21461),
            .I(N__21450));
    InMux I__4639 (
            .O(N__21458),
            .I(N__21447));
    LocalMux I__4638 (
            .O(N__21455),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv4 I__4637 (
            .O(N__21450),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__4636 (
            .O(N__21447),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    IoInMux I__4635 (
            .O(N__21440),
            .I(N__21437));
    LocalMux I__4634 (
            .O(N__21437),
            .I(N__21434));
    IoSpan4Mux I__4633 (
            .O(N__21434),
            .I(N__21431));
    Span4Mux_s2_v I__4632 (
            .O(N__21431),
            .I(N__21428));
    Sp12to4 I__4631 (
            .O(N__21428),
            .I(N__21425));
    Span12Mux_s10_v I__4630 (
            .O(N__21425),
            .I(N__21421));
    InMux I__4629 (
            .O(N__21424),
            .I(N__21418));
    Odrv12 I__4628 (
            .O(N__21421),
            .I(ppm_output_c));
    LocalMux I__4627 (
            .O(N__21418),
            .I(ppm_output_c));
    InMux I__4626 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__4625 (
            .O(N__21410),
            .I(N__21407));
    Odrv12 I__4624 (
            .O(N__21407),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__4623 (
            .O(N__21404),
            .I(N__21401));
    LocalMux I__4622 (
            .O(N__21401),
            .I(N__21397));
    InMux I__4621 (
            .O(N__21400),
            .I(N__21394));
    Span4Mux_v I__4620 (
            .O(N__21397),
            .I(N__21391));
    LocalMux I__4619 (
            .O(N__21394),
            .I(N__21388));
    Odrv4 I__4618 (
            .O(N__21391),
            .I(scaler_1_data_9));
    Odrv4 I__4617 (
            .O(N__21388),
            .I(scaler_1_data_9));
    InMux I__4616 (
            .O(N__21383),
            .I(N__21380));
    LocalMux I__4615 (
            .O(N__21380),
            .I(N__21376));
    InMux I__4614 (
            .O(N__21379),
            .I(N__21373));
    Span4Mux_h I__4613 (
            .O(N__21376),
            .I(N__21370));
    LocalMux I__4612 (
            .O(N__21373),
            .I(N__21367));
    Odrv4 I__4611 (
            .O(N__21370),
            .I(frame_decoder_CH3data_7));
    Odrv4 I__4610 (
            .O(N__21367),
            .I(frame_decoder_CH3data_7));
    InMux I__4609 (
            .O(N__21362),
            .I(N__21358));
    InMux I__4608 (
            .O(N__21361),
            .I(N__21355));
    LocalMux I__4607 (
            .O(N__21358),
            .I(N__21352));
    LocalMux I__4606 (
            .O(N__21355),
            .I(N__21349));
    Span4Mux_v I__4605 (
            .O(N__21352),
            .I(N__21346));
    Span4Mux_v I__4604 (
            .O(N__21349),
            .I(N__21343));
    Span4Mux_h I__4603 (
            .O(N__21346),
            .I(N__21338));
    Span4Mux_h I__4602 (
            .O(N__21343),
            .I(N__21338));
    Odrv4 I__4601 (
            .O(N__21338),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa ));
    InMux I__4600 (
            .O(N__21335),
            .I(N__21331));
    InMux I__4599 (
            .O(N__21334),
            .I(N__21328));
    LocalMux I__4598 (
            .O(N__21331),
            .I(N__21325));
    LocalMux I__4597 (
            .O(N__21328),
            .I(N__21322));
    Odrv12 I__4596 (
            .O(N__21325),
            .I(scaler_1_data_6));
    Odrv4 I__4595 (
            .O(N__21322),
            .I(scaler_1_data_6));
    InMux I__4594 (
            .O(N__21317),
            .I(N__21313));
    InMux I__4593 (
            .O(N__21316),
            .I(N__21310));
    LocalMux I__4592 (
            .O(N__21313),
            .I(N__21307));
    LocalMux I__4591 (
            .O(N__21310),
            .I(N__21304));
    Odrv4 I__4590 (
            .O(N__21307),
            .I(scaler_1_data_7));
    Odrv4 I__4589 (
            .O(N__21304),
            .I(scaler_1_data_7));
    InMux I__4588 (
            .O(N__21299),
            .I(N__21296));
    LocalMux I__4587 (
            .O(N__21296),
            .I(N__21293));
    Span4Mux_h I__4586 (
            .O(N__21293),
            .I(N__21290));
    Odrv4 I__4585 (
            .O(N__21290),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__4584 (
            .O(N__21287),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__4583 (
            .O(N__21284),
            .I(\ppm_encoder_1.un1_throttle_cry_7 ));
    InMux I__4582 (
            .O(N__21281),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__4581 (
            .O(N__21278),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__4580 (
            .O(N__21275),
            .I(N__21271));
    InMux I__4579 (
            .O(N__21274),
            .I(N__21268));
    LocalMux I__4578 (
            .O(N__21271),
            .I(N__21265));
    LocalMux I__4577 (
            .O(N__21268),
            .I(N__21262));
    Odrv12 I__4576 (
            .O(N__21265),
            .I(scaler_1_data_11));
    Odrv12 I__4575 (
            .O(N__21262),
            .I(scaler_1_data_11));
    InMux I__4574 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__4573 (
            .O(N__21254),
            .I(N__21251));
    Span4Mux_h I__4572 (
            .O(N__21251),
            .I(N__21248));
    Odrv4 I__4571 (
            .O(N__21248),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__4570 (
            .O(N__21245),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__4569 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__4568 (
            .O(N__21239),
            .I(N__21235));
    CascadeMux I__4567 (
            .O(N__21238),
            .I(N__21232));
    Span4Mux_h I__4566 (
            .O(N__21235),
            .I(N__21229));
    InMux I__4565 (
            .O(N__21232),
            .I(N__21226));
    Span4Mux_v I__4564 (
            .O(N__21229),
            .I(N__21221));
    LocalMux I__4563 (
            .O(N__21226),
            .I(N__21221));
    Odrv4 I__4562 (
            .O(N__21221),
            .I(scaler_1_data_12));
    InMux I__4561 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__4560 (
            .O(N__21215),
            .I(N__21212));
    Span4Mux_v I__4559 (
            .O(N__21212),
            .I(N__21209));
    Odrv4 I__4558 (
            .O(N__21209),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__4557 (
            .O(N__21206),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__4556 (
            .O(N__21203),
            .I(N__21199));
    InMux I__4555 (
            .O(N__21202),
            .I(N__21196));
    LocalMux I__4554 (
            .O(N__21199),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ));
    LocalMux I__4553 (
            .O(N__21196),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ));
    CascadeMux I__4552 (
            .O(N__21191),
            .I(N__21188));
    InMux I__4551 (
            .O(N__21188),
            .I(N__21185));
    LocalMux I__4550 (
            .O(N__21185),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__4549 (
            .O(N__21182),
            .I(N__21179));
    LocalMux I__4548 (
            .O(N__21179),
            .I(N__21175));
    InMux I__4547 (
            .O(N__21178),
            .I(N__21172));
    Span4Mux_v I__4546 (
            .O(N__21175),
            .I(N__21167));
    LocalMux I__4545 (
            .O(N__21172),
            .I(N__21167));
    Span4Mux_v I__4544 (
            .O(N__21167),
            .I(N__21164));
    Odrv4 I__4543 (
            .O(N__21164),
            .I(scaler_4_data_13));
    InMux I__4542 (
            .O(N__21161),
            .I(bfn_12_14_0_));
    InMux I__4541 (
            .O(N__21158),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__4540 (
            .O(N__21155),
            .I(N__21152));
    LocalMux I__4539 (
            .O(N__21152),
            .I(N__21149));
    Span4Mux_v I__4538 (
            .O(N__21149),
            .I(N__21146));
    Odrv4 I__4537 (
            .O(N__21146),
            .I(scaler_4_data_14));
    CEMux I__4536 (
            .O(N__21143),
            .I(N__21116));
    CEMux I__4535 (
            .O(N__21142),
            .I(N__21116));
    CEMux I__4534 (
            .O(N__21141),
            .I(N__21116));
    CEMux I__4533 (
            .O(N__21140),
            .I(N__21116));
    CEMux I__4532 (
            .O(N__21139),
            .I(N__21116));
    CEMux I__4531 (
            .O(N__21138),
            .I(N__21116));
    CEMux I__4530 (
            .O(N__21137),
            .I(N__21116));
    CEMux I__4529 (
            .O(N__21136),
            .I(N__21116));
    CEMux I__4528 (
            .O(N__21135),
            .I(N__21116));
    GlobalMux I__4527 (
            .O(N__21116),
            .I(N__21113));
    gio2CtrlBuf I__4526 (
            .O(N__21113),
            .I(pc_frame_decoder_dv_0_g));
    InMux I__4525 (
            .O(N__21110),
            .I(N__21104));
    InMux I__4524 (
            .O(N__21109),
            .I(N__21098));
    InMux I__4523 (
            .O(N__21108),
            .I(N__21095));
    InMux I__4522 (
            .O(N__21107),
            .I(N__21091));
    LocalMux I__4521 (
            .O(N__21104),
            .I(N__21088));
    InMux I__4520 (
            .O(N__21103),
            .I(N__21085));
    InMux I__4519 (
            .O(N__21102),
            .I(N__21082));
    InMux I__4518 (
            .O(N__21101),
            .I(N__21079));
    LocalMux I__4517 (
            .O(N__21098),
            .I(N__21076));
    LocalMux I__4516 (
            .O(N__21095),
            .I(N__21073));
    InMux I__4515 (
            .O(N__21094),
            .I(N__21070));
    LocalMux I__4514 (
            .O(N__21091),
            .I(N__21066));
    Span4Mux_v I__4513 (
            .O(N__21088),
            .I(N__21056));
    LocalMux I__4512 (
            .O(N__21085),
            .I(N__21056));
    LocalMux I__4511 (
            .O(N__21082),
            .I(N__21056));
    LocalMux I__4510 (
            .O(N__21079),
            .I(N__21056));
    Span4Mux_v I__4509 (
            .O(N__21076),
            .I(N__21049));
    Span4Mux_v I__4508 (
            .O(N__21073),
            .I(N__21049));
    LocalMux I__4507 (
            .O(N__21070),
            .I(N__21049));
    InMux I__4506 (
            .O(N__21069),
            .I(N__21046));
    Span4Mux_h I__4505 (
            .O(N__21066),
            .I(N__21043));
    InMux I__4504 (
            .O(N__21065),
            .I(N__21040));
    Span4Mux_v I__4503 (
            .O(N__21056),
            .I(N__21033));
    Span4Mux_h I__4502 (
            .O(N__21049),
            .I(N__21033));
    LocalMux I__4501 (
            .O(N__21046),
            .I(N__21033));
    Odrv4 I__4500 (
            .O(N__21043),
            .I(uart_pc_data_0));
    LocalMux I__4499 (
            .O(N__21040),
            .I(uart_pc_data_0));
    Odrv4 I__4498 (
            .O(N__21033),
            .I(uart_pc_data_0));
    InMux I__4497 (
            .O(N__21026),
            .I(N__21022));
    InMux I__4496 (
            .O(N__21025),
            .I(N__21019));
    LocalMux I__4495 (
            .O(N__21022),
            .I(N__21012));
    LocalMux I__4494 (
            .O(N__21019),
            .I(N__21012));
    InMux I__4493 (
            .O(N__21018),
            .I(N__21009));
    InMux I__4492 (
            .O(N__21017),
            .I(N__21006));
    Span4Mux_v I__4491 (
            .O(N__21012),
            .I(N__21001));
    LocalMux I__4490 (
            .O(N__21009),
            .I(N__21001));
    LocalMux I__4489 (
            .O(N__21006),
            .I(N__20998));
    Span4Mux_h I__4488 (
            .O(N__21001),
            .I(N__20995));
    Odrv4 I__4487 (
            .O(N__20998),
            .I(frame_decoder_CH3data_0));
    Odrv4 I__4486 (
            .O(N__20995),
            .I(frame_decoder_CH3data_0));
    InMux I__4485 (
            .O(N__20990),
            .I(N__20985));
    InMux I__4484 (
            .O(N__20989),
            .I(N__20982));
    InMux I__4483 (
            .O(N__20988),
            .I(N__20977));
    LocalMux I__4482 (
            .O(N__20985),
            .I(N__20971));
    LocalMux I__4481 (
            .O(N__20982),
            .I(N__20968));
    InMux I__4480 (
            .O(N__20981),
            .I(N__20965));
    InMux I__4479 (
            .O(N__20980),
            .I(N__20962));
    LocalMux I__4478 (
            .O(N__20977),
            .I(N__20959));
    InMux I__4477 (
            .O(N__20976),
            .I(N__20956));
    InMux I__4476 (
            .O(N__20975),
            .I(N__20952));
    InMux I__4475 (
            .O(N__20974),
            .I(N__20949));
    Span4Mux_v I__4474 (
            .O(N__20971),
            .I(N__20942));
    Span4Mux_v I__4473 (
            .O(N__20968),
            .I(N__20942));
    LocalMux I__4472 (
            .O(N__20965),
            .I(N__20942));
    LocalMux I__4471 (
            .O(N__20962),
            .I(N__20935));
    Span4Mux_h I__4470 (
            .O(N__20959),
            .I(N__20935));
    LocalMux I__4469 (
            .O(N__20956),
            .I(N__20935));
    InMux I__4468 (
            .O(N__20955),
            .I(N__20932));
    LocalMux I__4467 (
            .O(N__20952),
            .I(N__20927));
    LocalMux I__4466 (
            .O(N__20949),
            .I(N__20927));
    Span4Mux_h I__4465 (
            .O(N__20942),
            .I(N__20924));
    Span4Mux_v I__4464 (
            .O(N__20935),
            .I(N__20921));
    LocalMux I__4463 (
            .O(N__20932),
            .I(N__20918));
    Odrv12 I__4462 (
            .O(N__20927),
            .I(uart_pc_data_1));
    Odrv4 I__4461 (
            .O(N__20924),
            .I(uart_pc_data_1));
    Odrv4 I__4460 (
            .O(N__20921),
            .I(uart_pc_data_1));
    Odrv4 I__4459 (
            .O(N__20918),
            .I(uart_pc_data_1));
    InMux I__4458 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__4457 (
            .O(N__20906),
            .I(N__20903));
    Odrv4 I__4456 (
            .O(N__20903),
            .I(frame_decoder_CH3data_1));
    InMux I__4455 (
            .O(N__20900),
            .I(N__20894));
    InMux I__4454 (
            .O(N__20899),
            .I(N__20889));
    InMux I__4453 (
            .O(N__20898),
            .I(N__20886));
    InMux I__4452 (
            .O(N__20897),
            .I(N__20883));
    LocalMux I__4451 (
            .O(N__20894),
            .I(N__20879));
    InMux I__4450 (
            .O(N__20893),
            .I(N__20876));
    InMux I__4449 (
            .O(N__20892),
            .I(N__20873));
    LocalMux I__4448 (
            .O(N__20889),
            .I(N__20865));
    LocalMux I__4447 (
            .O(N__20886),
            .I(N__20865));
    LocalMux I__4446 (
            .O(N__20883),
            .I(N__20865));
    InMux I__4445 (
            .O(N__20882),
            .I(N__20862));
    Span4Mux_h I__4444 (
            .O(N__20879),
            .I(N__20855));
    LocalMux I__4443 (
            .O(N__20876),
            .I(N__20855));
    LocalMux I__4442 (
            .O(N__20873),
            .I(N__20855));
    InMux I__4441 (
            .O(N__20872),
            .I(N__20852));
    Span4Mux_v I__4440 (
            .O(N__20865),
            .I(N__20845));
    LocalMux I__4439 (
            .O(N__20862),
            .I(N__20845));
    Span4Mux_v I__4438 (
            .O(N__20855),
            .I(N__20842));
    LocalMux I__4437 (
            .O(N__20852),
            .I(N__20839));
    InMux I__4436 (
            .O(N__20851),
            .I(N__20836));
    InMux I__4435 (
            .O(N__20850),
            .I(N__20833));
    Odrv4 I__4434 (
            .O(N__20845),
            .I(uart_pc_data_2));
    Odrv4 I__4433 (
            .O(N__20842),
            .I(uart_pc_data_2));
    Odrv12 I__4432 (
            .O(N__20839),
            .I(uart_pc_data_2));
    LocalMux I__4431 (
            .O(N__20836),
            .I(uart_pc_data_2));
    LocalMux I__4430 (
            .O(N__20833),
            .I(uart_pc_data_2));
    InMux I__4429 (
            .O(N__20822),
            .I(N__20819));
    LocalMux I__4428 (
            .O(N__20819),
            .I(N__20816));
    Odrv4 I__4427 (
            .O(N__20816),
            .I(frame_decoder_CH3data_2));
    InMux I__4426 (
            .O(N__20813),
            .I(N__20805));
    InMux I__4425 (
            .O(N__20812),
            .I(N__20802));
    InMux I__4424 (
            .O(N__20811),
            .I(N__20799));
    InMux I__4423 (
            .O(N__20810),
            .I(N__20795));
    InMux I__4422 (
            .O(N__20809),
            .I(N__20792));
    InMux I__4421 (
            .O(N__20808),
            .I(N__20789));
    LocalMux I__4420 (
            .O(N__20805),
            .I(N__20781));
    LocalMux I__4419 (
            .O(N__20802),
            .I(N__20781));
    LocalMux I__4418 (
            .O(N__20799),
            .I(N__20781));
    InMux I__4417 (
            .O(N__20798),
            .I(N__20778));
    LocalMux I__4416 (
            .O(N__20795),
            .I(N__20773));
    LocalMux I__4415 (
            .O(N__20792),
            .I(N__20773));
    LocalMux I__4414 (
            .O(N__20789),
            .I(N__20770));
    InMux I__4413 (
            .O(N__20788),
            .I(N__20767));
    Span4Mux_v I__4412 (
            .O(N__20781),
            .I(N__20761));
    LocalMux I__4411 (
            .O(N__20778),
            .I(N__20761));
    Span4Mux_v I__4410 (
            .O(N__20773),
            .I(N__20758));
    Span12Mux_v I__4409 (
            .O(N__20770),
            .I(N__20753));
    LocalMux I__4408 (
            .O(N__20767),
            .I(N__20753));
    InMux I__4407 (
            .O(N__20766),
            .I(N__20750));
    Odrv4 I__4406 (
            .O(N__20761),
            .I(uart_pc_data_3));
    Odrv4 I__4405 (
            .O(N__20758),
            .I(uart_pc_data_3));
    Odrv12 I__4404 (
            .O(N__20753),
            .I(uart_pc_data_3));
    LocalMux I__4403 (
            .O(N__20750),
            .I(uart_pc_data_3));
    CascadeMux I__4402 (
            .O(N__20741),
            .I(N__20738));
    InMux I__4401 (
            .O(N__20738),
            .I(N__20735));
    LocalMux I__4400 (
            .O(N__20735),
            .I(N__20732));
    Odrv4 I__4399 (
            .O(N__20732),
            .I(frame_decoder_CH3data_3));
    InMux I__4398 (
            .O(N__20729),
            .I(N__20722));
    InMux I__4397 (
            .O(N__20728),
            .I(N__20717));
    InMux I__4396 (
            .O(N__20727),
            .I(N__20713));
    InMux I__4395 (
            .O(N__20726),
            .I(N__20710));
    InMux I__4394 (
            .O(N__20725),
            .I(N__20707));
    LocalMux I__4393 (
            .O(N__20722),
            .I(N__20704));
    InMux I__4392 (
            .O(N__20721),
            .I(N__20701));
    InMux I__4391 (
            .O(N__20720),
            .I(N__20698));
    LocalMux I__4390 (
            .O(N__20717),
            .I(N__20695));
    InMux I__4389 (
            .O(N__20716),
            .I(N__20692));
    LocalMux I__4388 (
            .O(N__20713),
            .I(N__20685));
    LocalMux I__4387 (
            .O(N__20710),
            .I(N__20685));
    LocalMux I__4386 (
            .O(N__20707),
            .I(N__20685));
    Span4Mux_h I__4385 (
            .O(N__20704),
            .I(N__20682));
    LocalMux I__4384 (
            .O(N__20701),
            .I(N__20679));
    LocalMux I__4383 (
            .O(N__20698),
            .I(N__20674));
    Span4Mux_h I__4382 (
            .O(N__20695),
            .I(N__20674));
    LocalMux I__4381 (
            .O(N__20692),
            .I(N__20670));
    Span4Mux_v I__4380 (
            .O(N__20685),
            .I(N__20667));
    Span4Mux_h I__4379 (
            .O(N__20682),
            .I(N__20664));
    Span4Mux_h I__4378 (
            .O(N__20679),
            .I(N__20659));
    Span4Mux_v I__4377 (
            .O(N__20674),
            .I(N__20659));
    InMux I__4376 (
            .O(N__20673),
            .I(N__20656));
    Odrv12 I__4375 (
            .O(N__20670),
            .I(uart_pc_data_4));
    Odrv4 I__4374 (
            .O(N__20667),
            .I(uart_pc_data_4));
    Odrv4 I__4373 (
            .O(N__20664),
            .I(uart_pc_data_4));
    Odrv4 I__4372 (
            .O(N__20659),
            .I(uart_pc_data_4));
    LocalMux I__4371 (
            .O(N__20656),
            .I(uart_pc_data_4));
    CascadeMux I__4370 (
            .O(N__20645),
            .I(N__20642));
    InMux I__4369 (
            .O(N__20642),
            .I(N__20639));
    LocalMux I__4368 (
            .O(N__20639),
            .I(N__20636));
    Odrv4 I__4367 (
            .O(N__20636),
            .I(frame_decoder_CH3data_4));
    InMux I__4366 (
            .O(N__20633),
            .I(N__20628));
    InMux I__4365 (
            .O(N__20632),
            .I(N__20625));
    InMux I__4364 (
            .O(N__20631),
            .I(N__20622));
    LocalMux I__4363 (
            .O(N__20628),
            .I(N__20614));
    LocalMux I__4362 (
            .O(N__20625),
            .I(N__20614));
    LocalMux I__4361 (
            .O(N__20622),
            .I(N__20610));
    InMux I__4360 (
            .O(N__20621),
            .I(N__20607));
    InMux I__4359 (
            .O(N__20620),
            .I(N__20603));
    InMux I__4358 (
            .O(N__20619),
            .I(N__20600));
    Span4Mux_v I__4357 (
            .O(N__20614),
            .I(N__20596));
    InMux I__4356 (
            .O(N__20613),
            .I(N__20593));
    Span4Mux_v I__4355 (
            .O(N__20610),
            .I(N__20588));
    LocalMux I__4354 (
            .O(N__20607),
            .I(N__20588));
    InMux I__4353 (
            .O(N__20606),
            .I(N__20585));
    LocalMux I__4352 (
            .O(N__20603),
            .I(N__20580));
    LocalMux I__4351 (
            .O(N__20600),
            .I(N__20580));
    InMux I__4350 (
            .O(N__20599),
            .I(N__20577));
    Span4Mux_v I__4349 (
            .O(N__20596),
            .I(N__20574));
    LocalMux I__4348 (
            .O(N__20593),
            .I(N__20571));
    Span4Mux_h I__4347 (
            .O(N__20588),
            .I(N__20568));
    LocalMux I__4346 (
            .O(N__20585),
            .I(N__20565));
    Span4Mux_v I__4345 (
            .O(N__20580),
            .I(N__20560));
    LocalMux I__4344 (
            .O(N__20577),
            .I(N__20560));
    Odrv4 I__4343 (
            .O(N__20574),
            .I(uart_pc_data_6));
    Odrv4 I__4342 (
            .O(N__20571),
            .I(uart_pc_data_6));
    Odrv4 I__4341 (
            .O(N__20568),
            .I(uart_pc_data_6));
    Odrv12 I__4340 (
            .O(N__20565),
            .I(uart_pc_data_6));
    Odrv4 I__4339 (
            .O(N__20560),
            .I(uart_pc_data_6));
    CascadeMux I__4338 (
            .O(N__20549),
            .I(N__20546));
    InMux I__4337 (
            .O(N__20546),
            .I(N__20543));
    LocalMux I__4336 (
            .O(N__20543),
            .I(N__20540));
    Odrv4 I__4335 (
            .O(N__20540),
            .I(frame_decoder_CH3data_6));
    InMux I__4334 (
            .O(N__20537),
            .I(N__20532));
    InMux I__4333 (
            .O(N__20536),
            .I(N__20528));
    InMux I__4332 (
            .O(N__20535),
            .I(N__20523));
    LocalMux I__4331 (
            .O(N__20532),
            .I(N__20520));
    InMux I__4330 (
            .O(N__20531),
            .I(N__20517));
    LocalMux I__4329 (
            .O(N__20528),
            .I(N__20514));
    InMux I__4328 (
            .O(N__20527),
            .I(N__20511));
    InMux I__4327 (
            .O(N__20526),
            .I(N__20508));
    LocalMux I__4326 (
            .O(N__20523),
            .I(N__20502));
    Span4Mux_v I__4325 (
            .O(N__20520),
            .I(N__20497));
    LocalMux I__4324 (
            .O(N__20517),
            .I(N__20497));
    Span4Mux_v I__4323 (
            .O(N__20514),
            .I(N__20490));
    LocalMux I__4322 (
            .O(N__20511),
            .I(N__20490));
    LocalMux I__4321 (
            .O(N__20508),
            .I(N__20490));
    InMux I__4320 (
            .O(N__20507),
            .I(N__20487));
    InMux I__4319 (
            .O(N__20506),
            .I(N__20484));
    CascadeMux I__4318 (
            .O(N__20505),
            .I(N__20480));
    Span4Mux_h I__4317 (
            .O(N__20502),
            .I(N__20477));
    Span4Mux_h I__4316 (
            .O(N__20497),
            .I(N__20470));
    Span4Mux_v I__4315 (
            .O(N__20490),
            .I(N__20470));
    LocalMux I__4314 (
            .O(N__20487),
            .I(N__20470));
    LocalMux I__4313 (
            .O(N__20484),
            .I(N__20467));
    InMux I__4312 (
            .O(N__20483),
            .I(N__20464));
    InMux I__4311 (
            .O(N__20480),
            .I(N__20461));
    Odrv4 I__4310 (
            .O(N__20477),
            .I(uart_pc_data_7));
    Odrv4 I__4309 (
            .O(N__20470),
            .I(uart_pc_data_7));
    Odrv12 I__4308 (
            .O(N__20467),
            .I(uart_pc_data_7));
    LocalMux I__4307 (
            .O(N__20464),
            .I(uart_pc_data_7));
    LocalMux I__4306 (
            .O(N__20461),
            .I(uart_pc_data_7));
    CascadeMux I__4305 (
            .O(N__20450),
            .I(N__20447));
    InMux I__4304 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__4303 (
            .O(N__20444),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNO_2 ));
    InMux I__4302 (
            .O(N__20441),
            .I(N__20436));
    CascadeMux I__4301 (
            .O(N__20440),
            .I(N__20433));
    InMux I__4300 (
            .O(N__20439),
            .I(N__20429));
    LocalMux I__4299 (
            .O(N__20436),
            .I(N__20426));
    InMux I__4298 (
            .O(N__20433),
            .I(N__20421));
    InMux I__4297 (
            .O(N__20432),
            .I(N__20421));
    LocalMux I__4296 (
            .O(N__20429),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__4295 (
            .O(N__20426),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__4294 (
            .O(N__20421),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__4293 (
            .O(N__20414),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__4292 (
            .O(N__20411),
            .I(N__20408));
    InMux I__4291 (
            .O(N__20408),
            .I(N__20402));
    InMux I__4290 (
            .O(N__20407),
            .I(N__20402));
    LocalMux I__4289 (
            .O(N__20402),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ));
    CascadeMux I__4288 (
            .O(N__20399),
            .I(N__20396));
    InMux I__4287 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__4286 (
            .O(N__20393),
            .I(N__20390));
    Span4Mux_h I__4285 (
            .O(N__20390),
            .I(N__20386));
    InMux I__4284 (
            .O(N__20389),
            .I(N__20383));
    Span4Mux_v I__4283 (
            .O(N__20386),
            .I(N__20380));
    LocalMux I__4282 (
            .O(N__20383),
            .I(N__20377));
    Span4Mux_v I__4281 (
            .O(N__20380),
            .I(N__20374));
    Span4Mux_v I__4280 (
            .O(N__20377),
            .I(N__20371));
    Odrv4 I__4279 (
            .O(N__20374),
            .I(scaler_4_data_7));
    Odrv4 I__4278 (
            .O(N__20371),
            .I(scaler_4_data_7));
    InMux I__4277 (
            .O(N__20366),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    CascadeMux I__4276 (
            .O(N__20363),
            .I(N__20360));
    InMux I__4275 (
            .O(N__20360),
            .I(N__20354));
    InMux I__4274 (
            .O(N__20359),
            .I(N__20354));
    LocalMux I__4273 (
            .O(N__20354),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ));
    InMux I__4272 (
            .O(N__20351),
            .I(N__20348));
    LocalMux I__4271 (
            .O(N__20348),
            .I(N__20344));
    InMux I__4270 (
            .O(N__20347),
            .I(N__20341));
    Span4Mux_v I__4269 (
            .O(N__20344),
            .I(N__20336));
    LocalMux I__4268 (
            .O(N__20341),
            .I(N__20336));
    Span4Mux_v I__4267 (
            .O(N__20336),
            .I(N__20333));
    Odrv4 I__4266 (
            .O(N__20333),
            .I(scaler_4_data_8));
    InMux I__4265 (
            .O(N__20330),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    CascadeMux I__4264 (
            .O(N__20327),
            .I(N__20324));
    InMux I__4263 (
            .O(N__20324),
            .I(N__20318));
    InMux I__4262 (
            .O(N__20323),
            .I(N__20318));
    LocalMux I__4261 (
            .O(N__20318),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNI15MI ));
    InMux I__4260 (
            .O(N__20315),
            .I(N__20312));
    LocalMux I__4259 (
            .O(N__20312),
            .I(N__20308));
    InMux I__4258 (
            .O(N__20311),
            .I(N__20305));
    Span4Mux_v I__4257 (
            .O(N__20308),
            .I(N__20300));
    LocalMux I__4256 (
            .O(N__20305),
            .I(N__20300));
    Span4Mux_v I__4255 (
            .O(N__20300),
            .I(N__20297));
    Odrv4 I__4254 (
            .O(N__20297),
            .I(scaler_4_data_9));
    InMux I__4253 (
            .O(N__20294),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__4252 (
            .O(N__20291),
            .I(N__20288));
    InMux I__4251 (
            .O(N__20288),
            .I(N__20282));
    InMux I__4250 (
            .O(N__20287),
            .I(N__20282));
    LocalMux I__4249 (
            .O(N__20282),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNI49NI ));
    InMux I__4248 (
            .O(N__20279),
            .I(N__20275));
    InMux I__4247 (
            .O(N__20278),
            .I(N__20272));
    LocalMux I__4246 (
            .O(N__20275),
            .I(N__20269));
    LocalMux I__4245 (
            .O(N__20272),
            .I(N__20266));
    Span12Mux_h I__4244 (
            .O(N__20269),
            .I(N__20263));
    Span4Mux_v I__4243 (
            .O(N__20266),
            .I(N__20260));
    Odrv12 I__4242 (
            .O(N__20263),
            .I(scaler_4_data_10));
    Odrv4 I__4241 (
            .O(N__20260),
            .I(scaler_4_data_10));
    InMux I__4240 (
            .O(N__20255),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__4239 (
            .O(N__20252),
            .I(N__20249));
    InMux I__4238 (
            .O(N__20249),
            .I(N__20243));
    InMux I__4237 (
            .O(N__20248),
            .I(N__20243));
    LocalMux I__4236 (
            .O(N__20243),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ));
    InMux I__4235 (
            .O(N__20240),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__4234 (
            .O(N__20237),
            .I(N__20234));
    InMux I__4233 (
            .O(N__20234),
            .I(N__20228));
    InMux I__4232 (
            .O(N__20233),
            .I(N__20228));
    LocalMux I__4231 (
            .O(N__20228),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ));
    InMux I__4230 (
            .O(N__20225),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__4229 (
            .O(N__20222),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__4228 (
            .O(N__20219),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__4227 (
            .O(N__20216),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__4226 (
            .O(N__20213),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__4225 (
            .O(N__20210),
            .I(bfn_11_30_0_));
    InMux I__4224 (
            .O(N__20207),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__4223 (
            .O(N__20204),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__4222 (
            .O(N__20201),
            .I(N__20192));
    SRMux I__4221 (
            .O(N__20200),
            .I(N__20192));
    SRMux I__4220 (
            .O(N__20199),
            .I(N__20192));
    GlobalMux I__4219 (
            .O(N__20192),
            .I(N__20189));
    gio2CtrlBuf I__4218 (
            .O(N__20189),
            .I(\ppm_encoder_1.N_228_g ));
    InMux I__4217 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__4216 (
            .O(N__20183),
            .I(N__20180));
    Span4Mux_s1_v I__4215 (
            .O(N__20180),
            .I(N__20177));
    Span4Mux_h I__4214 (
            .O(N__20177),
            .I(N__20173));
    CascadeMux I__4213 (
            .O(N__20176),
            .I(N__20170));
    Sp12to4 I__4212 (
            .O(N__20173),
            .I(N__20162));
    InMux I__4211 (
            .O(N__20170),
            .I(N__20153));
    InMux I__4210 (
            .O(N__20169),
            .I(N__20153));
    InMux I__4209 (
            .O(N__20168),
            .I(N__20153));
    InMux I__4208 (
            .O(N__20167),
            .I(N__20153));
    InMux I__4207 (
            .O(N__20166),
            .I(N__20148));
    InMux I__4206 (
            .O(N__20165),
            .I(N__20148));
    Span12Mux_s10_v I__4205 (
            .O(N__20162),
            .I(N__20145));
    LocalMux I__4204 (
            .O(N__20153),
            .I(pc_frame_decoder_dv));
    LocalMux I__4203 (
            .O(N__20148),
            .I(pc_frame_decoder_dv));
    Odrv12 I__4202 (
            .O(N__20145),
            .I(pc_frame_decoder_dv));
    IoInMux I__4201 (
            .O(N__20138),
            .I(N__20135));
    LocalMux I__4200 (
            .O(N__20135),
            .I(pc_frame_decoder_dv_0));
    CascadeMux I__4199 (
            .O(N__20132),
            .I(N__20129));
    InMux I__4198 (
            .O(N__20129),
            .I(N__20126));
    LocalMux I__4197 (
            .O(N__20126),
            .I(frame_decoder_OFF4data_4));
    CEMux I__4196 (
            .O(N__20123),
            .I(N__20120));
    LocalMux I__4195 (
            .O(N__20120),
            .I(N__20116));
    CEMux I__4194 (
            .O(N__20119),
            .I(N__20113));
    Span4Mux_h I__4193 (
            .O(N__20116),
            .I(N__20110));
    LocalMux I__4192 (
            .O(N__20113),
            .I(N__20107));
    Odrv4 I__4191 (
            .O(N__20110),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    Odrv4 I__4190 (
            .O(N__20107),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    CascadeMux I__4189 (
            .O(N__20102),
            .I(N__20097));
    InMux I__4188 (
            .O(N__20101),
            .I(N__20093));
    InMux I__4187 (
            .O(N__20100),
            .I(N__20088));
    InMux I__4186 (
            .O(N__20097),
            .I(N__20088));
    InMux I__4185 (
            .O(N__20096),
            .I(N__20085));
    LocalMux I__4184 (
            .O(N__20093),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__4183 (
            .O(N__20088),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__4182 (
            .O(N__20085),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__4181 (
            .O(N__20078),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__4180 (
            .O(N__20075),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__4179 (
            .O(N__20072),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__4178 (
            .O(N__20069),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__4177 (
            .O(N__20066),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__4176 (
            .O(N__20063),
            .I(bfn_11_29_0_));
    InMux I__4175 (
            .O(N__20060),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__4174 (
            .O(N__20057),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__4173 (
            .O(N__20054),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    CascadeMux I__4172 (
            .O(N__20051),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_ ));
    CascadeMux I__4171 (
            .O(N__20048),
            .I(N__20045));
    InMux I__4170 (
            .O(N__20045),
            .I(N__20042));
    LocalMux I__4169 (
            .O(N__20042),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__4168 (
            .O(N__20039),
            .I(N__20036));
    LocalMux I__4167 (
            .O(N__20036),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__4166 (
            .O(N__20033),
            .I(N__20030));
    LocalMux I__4165 (
            .O(N__20030),
            .I(N__20027));
    Span4Mux_v I__4164 (
            .O(N__20027),
            .I(N__20021));
    InMux I__4163 (
            .O(N__20026),
            .I(N__20014));
    InMux I__4162 (
            .O(N__20025),
            .I(N__20014));
    InMux I__4161 (
            .O(N__20024),
            .I(N__20014));
    Odrv4 I__4160 (
            .O(N__20021),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    LocalMux I__4159 (
            .O(N__20014),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__4158 (
            .O(N__20009),
            .I(N__20006));
    LocalMux I__4157 (
            .O(N__20006),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__4156 (
            .O(N__20003),
            .I(N__19999));
    InMux I__4155 (
            .O(N__20002),
            .I(N__19996));
    LocalMux I__4154 (
            .O(N__19999),
            .I(N__19990));
    LocalMux I__4153 (
            .O(N__19996),
            .I(N__19990));
    InMux I__4152 (
            .O(N__19995),
            .I(N__19985));
    Span4Mux_h I__4151 (
            .O(N__19990),
            .I(N__19982));
    InMux I__4150 (
            .O(N__19989),
            .I(N__19977));
    InMux I__4149 (
            .O(N__19988),
            .I(N__19977));
    LocalMux I__4148 (
            .O(N__19985),
            .I(N__19974));
    Odrv4 I__4147 (
            .O(N__19982),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    LocalMux I__4146 (
            .O(N__19977),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__4145 (
            .O(N__19974),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    CascadeMux I__4144 (
            .O(N__19967),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_ ));
    CascadeMux I__4143 (
            .O(N__19964),
            .I(N__19961));
    InMux I__4142 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__4141 (
            .O(N__19958),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    CascadeMux I__4140 (
            .O(N__19955),
            .I(N__19951));
    InMux I__4139 (
            .O(N__19954),
            .I(N__19948));
    InMux I__4138 (
            .O(N__19951),
            .I(N__19945));
    LocalMux I__4137 (
            .O(N__19948),
            .I(N__19940));
    LocalMux I__4136 (
            .O(N__19945),
            .I(N__19940));
    Span12Mux_s8_v I__4135 (
            .O(N__19940),
            .I(N__19937));
    Odrv12 I__4134 (
            .O(N__19937),
            .I(\ppm_encoder_1.N_614_i ));
    CascadeMux I__4133 (
            .O(N__19934),
            .I(N__19929));
    InMux I__4132 (
            .O(N__19933),
            .I(N__19926));
    InMux I__4131 (
            .O(N__19932),
            .I(N__19922));
    InMux I__4130 (
            .O(N__19929),
            .I(N__19919));
    LocalMux I__4129 (
            .O(N__19926),
            .I(N__19916));
    InMux I__4128 (
            .O(N__19925),
            .I(N__19913));
    LocalMux I__4127 (
            .O(N__19922),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__4126 (
            .O(N__19919),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__4125 (
            .O(N__19916),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__4124 (
            .O(N__19913),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__4123 (
            .O(N__19904),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__4122 (
            .O(N__19901),
            .I(N__19895));
    InMux I__4121 (
            .O(N__19900),
            .I(N__19890));
    InMux I__4120 (
            .O(N__19899),
            .I(N__19890));
    InMux I__4119 (
            .O(N__19898),
            .I(N__19887));
    LocalMux I__4118 (
            .O(N__19895),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__4117 (
            .O(N__19890),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__4116 (
            .O(N__19887),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__4115 (
            .O(N__19880),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    CascadeMux I__4114 (
            .O(N__19877),
            .I(N__19874));
    InMux I__4113 (
            .O(N__19874),
            .I(N__19870));
    InMux I__4112 (
            .O(N__19873),
            .I(N__19867));
    LocalMux I__4111 (
            .O(N__19870),
            .I(N__19864));
    LocalMux I__4110 (
            .O(N__19867),
            .I(N__19861));
    Span12Mux_s10_v I__4109 (
            .O(N__19864),
            .I(N__19858));
    Span12Mux_v I__4108 (
            .O(N__19861),
            .I(N__19855));
    Odrv12 I__4107 (
            .O(N__19858),
            .I(scaler_2_data_12));
    Odrv12 I__4106 (
            .O(N__19855),
            .I(scaler_2_data_12));
    InMux I__4105 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__4104 (
            .O(N__19847),
            .I(N__19844));
    Span4Mux_h I__4103 (
            .O(N__19844),
            .I(N__19841));
    Odrv4 I__4102 (
            .O(N__19841),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__4101 (
            .O(N__19838),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__4100 (
            .O(N__19835),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__4099 (
            .O(N__19832),
            .I(N__19829));
    LocalMux I__4098 (
            .O(N__19829),
            .I(N__19826));
    Span4Mux_v I__4097 (
            .O(N__19826),
            .I(N__19823));
    Span4Mux_v I__4096 (
            .O(N__19823),
            .I(N__19820));
    Span4Mux_v I__4095 (
            .O(N__19820),
            .I(N__19817));
    Odrv4 I__4094 (
            .O(N__19817),
            .I(scaler_2_data_14));
    InMux I__4093 (
            .O(N__19814),
            .I(bfn_11_25_0_));
    InMux I__4092 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__4091 (
            .O(N__19808),
            .I(N__19805));
    Span4Mux_v I__4090 (
            .O(N__19805),
            .I(N__19802));
    Span4Mux_h I__4089 (
            .O(N__19802),
            .I(N__19799));
    Odrv4 I__4088 (
            .O(N__19799),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__4087 (
            .O(N__19796),
            .I(N__19793));
    LocalMux I__4086 (
            .O(N__19793),
            .I(N__19790));
    Span4Mux_v I__4085 (
            .O(N__19790),
            .I(N__19787));
    Odrv4 I__4084 (
            .O(N__19787),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__4083 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__4082 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__4081 (
            .O(N__19778),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__4080 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__4079 (
            .O(N__19772),
            .I(N__19769));
    Span4Mux_h I__4078 (
            .O(N__19769),
            .I(N__19766));
    Odrv4 I__4077 (
            .O(N__19766),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    CascadeMux I__4076 (
            .O(N__19763),
            .I(N__19760));
    InMux I__4075 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__4074 (
            .O(N__19757),
            .I(N__19754));
    Span4Mux_s3_v I__4073 (
            .O(N__19754),
            .I(N__19751));
    Odrv4 I__4072 (
            .O(N__19751),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__4071 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__4070 (
            .O(N__19745),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    CascadeMux I__4069 (
            .O(N__19742),
            .I(N__19739));
    InMux I__4068 (
            .O(N__19739),
            .I(N__19736));
    LocalMux I__4067 (
            .O(N__19736),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__4066 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__4065 (
            .O(N__19730),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__4064 (
            .O(N__19727),
            .I(N__19724));
    LocalMux I__4063 (
            .O(N__19724),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__4062 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__4061 (
            .O(N__19718),
            .I(N__19715));
    Span4Mux_h I__4060 (
            .O(N__19715),
            .I(N__19712));
    Span4Mux_h I__4059 (
            .O(N__19712),
            .I(N__19709));
    Odrv4 I__4058 (
            .O(N__19709),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    CascadeMux I__4057 (
            .O(N__19706),
            .I(N__19696));
    InMux I__4056 (
            .O(N__19705),
            .I(N__19687));
    InMux I__4055 (
            .O(N__19704),
            .I(N__19687));
    InMux I__4054 (
            .O(N__19703),
            .I(N__19684));
    CascadeMux I__4053 (
            .O(N__19702),
            .I(N__19681));
    InMux I__4052 (
            .O(N__19701),
            .I(N__19678));
    InMux I__4051 (
            .O(N__19700),
            .I(N__19673));
    InMux I__4050 (
            .O(N__19699),
            .I(N__19673));
    InMux I__4049 (
            .O(N__19696),
            .I(N__19663));
    InMux I__4048 (
            .O(N__19695),
            .I(N__19658));
    InMux I__4047 (
            .O(N__19694),
            .I(N__19658));
    InMux I__4046 (
            .O(N__19693),
            .I(N__19653));
    InMux I__4045 (
            .O(N__19692),
            .I(N__19653));
    LocalMux I__4044 (
            .O(N__19687),
            .I(N__19648));
    LocalMux I__4043 (
            .O(N__19684),
            .I(N__19648));
    InMux I__4042 (
            .O(N__19681),
            .I(N__19645));
    LocalMux I__4041 (
            .O(N__19678),
            .I(N__19642));
    LocalMux I__4040 (
            .O(N__19673),
            .I(N__19639));
    InMux I__4039 (
            .O(N__19672),
            .I(N__19634));
    InMux I__4038 (
            .O(N__19671),
            .I(N__19634));
    InMux I__4037 (
            .O(N__19670),
            .I(N__19629));
    InMux I__4036 (
            .O(N__19669),
            .I(N__19629));
    InMux I__4035 (
            .O(N__19668),
            .I(N__19622));
    InMux I__4034 (
            .O(N__19667),
            .I(N__19622));
    InMux I__4033 (
            .O(N__19666),
            .I(N__19622));
    LocalMux I__4032 (
            .O(N__19663),
            .I(N__19613));
    LocalMux I__4031 (
            .O(N__19658),
            .I(N__19613));
    LocalMux I__4030 (
            .O(N__19653),
            .I(N__19613));
    Span4Mux_h I__4029 (
            .O(N__19648),
            .I(N__19613));
    LocalMux I__4028 (
            .O(N__19645),
            .I(N__19606));
    Span4Mux_v I__4027 (
            .O(N__19642),
            .I(N__19606));
    Span4Mux_h I__4026 (
            .O(N__19639),
            .I(N__19606));
    LocalMux I__4025 (
            .O(N__19634),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__4024 (
            .O(N__19629),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__4023 (
            .O(N__19622),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__4022 (
            .O(N__19613),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__4021 (
            .O(N__19606),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__4020 (
            .O(N__19595),
            .I(N__19592));
    LocalMux I__4019 (
            .O(N__19592),
            .I(N__19589));
    Span4Mux_h I__4018 (
            .O(N__19589),
            .I(N__19586));
    Odrv4 I__4017 (
            .O(N__19586),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    CascadeMux I__4016 (
            .O(N__19583),
            .I(N__19577));
    CascadeMux I__4015 (
            .O(N__19582),
            .I(N__19572));
    CascadeMux I__4014 (
            .O(N__19581),
            .I(N__19569));
    CascadeMux I__4013 (
            .O(N__19580),
            .I(N__19563));
    InMux I__4012 (
            .O(N__19577),
            .I(N__19558));
    InMux I__4011 (
            .O(N__19576),
            .I(N__19553));
    InMux I__4010 (
            .O(N__19575),
            .I(N__19553));
    InMux I__4009 (
            .O(N__19572),
            .I(N__19544));
    InMux I__4008 (
            .O(N__19569),
            .I(N__19544));
    CascadeMux I__4007 (
            .O(N__19568),
            .I(N__19541));
    CascadeMux I__4006 (
            .O(N__19567),
            .I(N__19538));
    CascadeMux I__4005 (
            .O(N__19566),
            .I(N__19535));
    InMux I__4004 (
            .O(N__19563),
            .I(N__19532));
    InMux I__4003 (
            .O(N__19562),
            .I(N__19527));
    InMux I__4002 (
            .O(N__19561),
            .I(N__19527));
    LocalMux I__4001 (
            .O(N__19558),
            .I(N__19522));
    LocalMux I__4000 (
            .O(N__19553),
            .I(N__19522));
    CascadeMux I__3999 (
            .O(N__19552),
            .I(N__19519));
    CascadeMux I__3998 (
            .O(N__19551),
            .I(N__19516));
    InMux I__3997 (
            .O(N__19550),
            .I(N__19512));
    CascadeMux I__3996 (
            .O(N__19549),
            .I(N__19509));
    LocalMux I__3995 (
            .O(N__19544),
            .I(N__19506));
    InMux I__3994 (
            .O(N__19541),
            .I(N__19501));
    InMux I__3993 (
            .O(N__19538),
            .I(N__19501));
    InMux I__3992 (
            .O(N__19535),
            .I(N__19498));
    LocalMux I__3991 (
            .O(N__19532),
            .I(N__19491));
    LocalMux I__3990 (
            .O(N__19527),
            .I(N__19491));
    Span4Mux_v I__3989 (
            .O(N__19522),
            .I(N__19488));
    InMux I__3988 (
            .O(N__19519),
            .I(N__19483));
    InMux I__3987 (
            .O(N__19516),
            .I(N__19483));
    InMux I__3986 (
            .O(N__19515),
            .I(N__19480));
    LocalMux I__3985 (
            .O(N__19512),
            .I(N__19477));
    InMux I__3984 (
            .O(N__19509),
            .I(N__19474));
    Span4Mux_v I__3983 (
            .O(N__19506),
            .I(N__19470));
    LocalMux I__3982 (
            .O(N__19501),
            .I(N__19465));
    LocalMux I__3981 (
            .O(N__19498),
            .I(N__19465));
    InMux I__3980 (
            .O(N__19497),
            .I(N__19460));
    InMux I__3979 (
            .O(N__19496),
            .I(N__19460));
    Span4Mux_v I__3978 (
            .O(N__19491),
            .I(N__19451));
    Span4Mux_h I__3977 (
            .O(N__19488),
            .I(N__19451));
    LocalMux I__3976 (
            .O(N__19483),
            .I(N__19451));
    LocalMux I__3975 (
            .O(N__19480),
            .I(N__19451));
    Span4Mux_h I__3974 (
            .O(N__19477),
            .I(N__19446));
    LocalMux I__3973 (
            .O(N__19474),
            .I(N__19446));
    InMux I__3972 (
            .O(N__19473),
            .I(N__19443));
    Odrv4 I__3971 (
            .O(N__19470),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv12 I__3970 (
            .O(N__19465),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__3969 (
            .O(N__19460),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__3968 (
            .O(N__19451),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__3967 (
            .O(N__19446),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__3966 (
            .O(N__19443),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__3965 (
            .O(N__19430),
            .I(N__19427));
    LocalMux I__3964 (
            .O(N__19427),
            .I(N__19424));
    Span4Mux_h I__3963 (
            .O(N__19424),
            .I(N__19421));
    Odrv4 I__3962 (
            .O(N__19421),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__3961 (
            .O(N__19418),
            .I(N__19412));
    InMux I__3960 (
            .O(N__19417),
            .I(N__19412));
    LocalMux I__3959 (
            .O(N__19412),
            .I(N__19408));
    InMux I__3958 (
            .O(N__19411),
            .I(N__19405));
    Span4Mux_h I__3957 (
            .O(N__19408),
            .I(N__19402));
    LocalMux I__3956 (
            .O(N__19405),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__3955 (
            .O(N__19402),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__3954 (
            .O(N__19397),
            .I(N__19393));
    InMux I__3953 (
            .O(N__19396),
            .I(N__19390));
    LocalMux I__3952 (
            .O(N__19393),
            .I(N__19387));
    LocalMux I__3951 (
            .O(N__19390),
            .I(N__19384));
    Span4Mux_v I__3950 (
            .O(N__19387),
            .I(N__19381));
    Span4Mux_v I__3949 (
            .O(N__19384),
            .I(N__19378));
    Span4Mux_v I__3948 (
            .O(N__19381),
            .I(N__19375));
    Span4Mux_v I__3947 (
            .O(N__19378),
            .I(N__19372));
    Span4Mux_v I__3946 (
            .O(N__19375),
            .I(N__19369));
    Odrv4 I__3945 (
            .O(N__19372),
            .I(scaler_2_data_6));
    Odrv4 I__3944 (
            .O(N__19369),
            .I(scaler_2_data_6));
    CascadeMux I__3943 (
            .O(N__19364),
            .I(N__19361));
    InMux I__3942 (
            .O(N__19361),
            .I(N__19357));
    InMux I__3941 (
            .O(N__19360),
            .I(N__19354));
    LocalMux I__3940 (
            .O(N__19357),
            .I(N__19351));
    LocalMux I__3939 (
            .O(N__19354),
            .I(N__19348));
    Span4Mux_v I__3938 (
            .O(N__19351),
            .I(N__19343));
    Span4Mux_v I__3937 (
            .O(N__19348),
            .I(N__19343));
    Span4Mux_v I__3936 (
            .O(N__19343),
            .I(N__19340));
    Odrv4 I__3935 (
            .O(N__19340),
            .I(scaler_2_data_7));
    InMux I__3934 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__3933 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__3932 (
            .O(N__19331),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__3931 (
            .O(N__19328),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__3930 (
            .O(N__19325),
            .I(N__19321));
    InMux I__3929 (
            .O(N__19324),
            .I(N__19318));
    LocalMux I__3928 (
            .O(N__19321),
            .I(N__19315));
    LocalMux I__3927 (
            .O(N__19318),
            .I(N__19312));
    Sp12to4 I__3926 (
            .O(N__19315),
            .I(N__19307));
    Span12Mux_h I__3925 (
            .O(N__19312),
            .I(N__19307));
    Odrv12 I__3924 (
            .O(N__19307),
            .I(scaler_2_data_8));
    InMux I__3923 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__3922 (
            .O(N__19301),
            .I(N__19298));
    Span4Mux_h I__3921 (
            .O(N__19298),
            .I(N__19295));
    Span4Mux_v I__3920 (
            .O(N__19295),
            .I(N__19292));
    Odrv4 I__3919 (
            .O(N__19292),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__3918 (
            .O(N__19289),
            .I(\ppm_encoder_1.un1_aileron_cry_7 ));
    InMux I__3917 (
            .O(N__19286),
            .I(N__19282));
    InMux I__3916 (
            .O(N__19285),
            .I(N__19279));
    LocalMux I__3915 (
            .O(N__19282),
            .I(N__19276));
    LocalMux I__3914 (
            .O(N__19279),
            .I(N__19271));
    Span4Mux_v I__3913 (
            .O(N__19276),
            .I(N__19271));
    Span4Mux_v I__3912 (
            .O(N__19271),
            .I(N__19268));
    Odrv4 I__3911 (
            .O(N__19268),
            .I(scaler_2_data_9));
    InMux I__3910 (
            .O(N__19265),
            .I(N__19262));
    LocalMux I__3909 (
            .O(N__19262),
            .I(N__19259));
    Span4Mux_v I__3908 (
            .O(N__19259),
            .I(N__19256));
    Odrv4 I__3907 (
            .O(N__19256),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__3906 (
            .O(N__19253),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    CascadeMux I__3905 (
            .O(N__19250),
            .I(N__19247));
    InMux I__3904 (
            .O(N__19247),
            .I(N__19243));
    InMux I__3903 (
            .O(N__19246),
            .I(N__19240));
    LocalMux I__3902 (
            .O(N__19243),
            .I(N__19235));
    LocalMux I__3901 (
            .O(N__19240),
            .I(N__19235));
    Span4Mux_v I__3900 (
            .O(N__19235),
            .I(N__19232));
    Span4Mux_v I__3899 (
            .O(N__19232),
            .I(N__19229));
    Odrv4 I__3898 (
            .O(N__19229),
            .I(scaler_2_data_10));
    InMux I__3897 (
            .O(N__19226),
            .I(N__19223));
    LocalMux I__3896 (
            .O(N__19223),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__3895 (
            .O(N__19220),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    CascadeMux I__3894 (
            .O(N__19217),
            .I(N__19214));
    InMux I__3893 (
            .O(N__19214),
            .I(N__19210));
    InMux I__3892 (
            .O(N__19213),
            .I(N__19207));
    LocalMux I__3891 (
            .O(N__19210),
            .I(N__19204));
    LocalMux I__3890 (
            .O(N__19207),
            .I(N__19201));
    Span4Mux_h I__3889 (
            .O(N__19204),
            .I(N__19196));
    Span4Mux_v I__3888 (
            .O(N__19201),
            .I(N__19196));
    Span4Mux_v I__3887 (
            .O(N__19196),
            .I(N__19193));
    Odrv4 I__3886 (
            .O(N__19193),
            .I(scaler_2_data_11));
    InMux I__3885 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__3884 (
            .O(N__19187),
            .I(N__19184));
    Span4Mux_h I__3883 (
            .O(N__19184),
            .I(N__19181));
    Odrv4 I__3882 (
            .O(N__19181),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__3881 (
            .O(N__19178),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    CascadeMux I__3880 (
            .O(N__19175),
            .I(N__19171));
    InMux I__3879 (
            .O(N__19174),
            .I(N__19168));
    InMux I__3878 (
            .O(N__19171),
            .I(N__19165));
    LocalMux I__3877 (
            .O(N__19168),
            .I(N__19162));
    LocalMux I__3876 (
            .O(N__19165),
            .I(N__19159));
    Odrv4 I__3875 (
            .O(N__19162),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    Odrv4 I__3874 (
            .O(N__19159),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    InMux I__3873 (
            .O(N__19154),
            .I(N__19151));
    LocalMux I__3872 (
            .O(N__19151),
            .I(N__19148));
    Span4Mux_h I__3871 (
            .O(N__19148),
            .I(N__19143));
    InMux I__3870 (
            .O(N__19147),
            .I(N__19138));
    InMux I__3869 (
            .O(N__19146),
            .I(N__19138));
    Odrv4 I__3868 (
            .O(N__19143),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    LocalMux I__3867 (
            .O(N__19138),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__3866 (
            .O(N__19133),
            .I(N__19128));
    InMux I__3865 (
            .O(N__19132),
            .I(N__19125));
    InMux I__3864 (
            .O(N__19131),
            .I(N__19122));
    LocalMux I__3863 (
            .O(N__19128),
            .I(N__19119));
    LocalMux I__3862 (
            .O(N__19125),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    LocalMux I__3861 (
            .O(N__19122),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__3860 (
            .O(N__19119),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__3859 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__3858 (
            .O(N__19109),
            .I(N__19106));
    Span4Mux_h I__3857 (
            .O(N__19106),
            .I(N__19103));
    Odrv4 I__3856 (
            .O(N__19103),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ));
    CascadeMux I__3855 (
            .O(N__19100),
            .I(N__19097));
    InMux I__3854 (
            .O(N__19097),
            .I(N__19094));
    LocalMux I__3853 (
            .O(N__19094),
            .I(N__19089));
    InMux I__3852 (
            .O(N__19093),
            .I(N__19084));
    InMux I__3851 (
            .O(N__19092),
            .I(N__19084));
    Odrv4 I__3850 (
            .O(N__19089),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    LocalMux I__3849 (
            .O(N__19084),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    InMux I__3848 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__3847 (
            .O(N__19076),
            .I(N__19073));
    Span12Mux_v I__3846 (
            .O(N__19073),
            .I(N__19068));
    InMux I__3845 (
            .O(N__19072),
            .I(N__19063));
    InMux I__3844 (
            .O(N__19071),
            .I(N__19063));
    Odrv12 I__3843 (
            .O(N__19068),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    LocalMux I__3842 (
            .O(N__19063),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__3841 (
            .O(N__19058),
            .I(N__19055));
    LocalMux I__3840 (
            .O(N__19055),
            .I(N__19051));
    InMux I__3839 (
            .O(N__19054),
            .I(N__19048));
    Span4Mux_h I__3838 (
            .O(N__19051),
            .I(N__19043));
    LocalMux I__3837 (
            .O(N__19048),
            .I(N__19043));
    Span4Mux_h I__3836 (
            .O(N__19043),
            .I(N__19040));
    Odrv4 I__3835 (
            .O(N__19040),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    CascadeMux I__3834 (
            .O(N__19037),
            .I(N__19033));
    InMux I__3833 (
            .O(N__19036),
            .I(N__19029));
    InMux I__3832 (
            .O(N__19033),
            .I(N__19026));
    CascadeMux I__3831 (
            .O(N__19032),
            .I(N__19023));
    LocalMux I__3830 (
            .O(N__19029),
            .I(N__19020));
    LocalMux I__3829 (
            .O(N__19026),
            .I(N__19017));
    InMux I__3828 (
            .O(N__19023),
            .I(N__19014));
    Span4Mux_v I__3827 (
            .O(N__19020),
            .I(N__19011));
    Span4Mux_h I__3826 (
            .O(N__19017),
            .I(N__19008));
    LocalMux I__3825 (
            .O(N__19014),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__3824 (
            .O(N__19011),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__3823 (
            .O(N__19008),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    CascadeMux I__3822 (
            .O(N__19001),
            .I(N__18998));
    InMux I__3821 (
            .O(N__18998),
            .I(N__18995));
    LocalMux I__3820 (
            .O(N__18995),
            .I(N__18992));
    Span4Mux_h I__3819 (
            .O(N__18992),
            .I(N__18989));
    Span4Mux_h I__3818 (
            .O(N__18989),
            .I(N__18984));
    InMux I__3817 (
            .O(N__18988),
            .I(N__18979));
    InMux I__3816 (
            .O(N__18987),
            .I(N__18979));
    Odrv4 I__3815 (
            .O(N__18984),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    LocalMux I__3814 (
            .O(N__18979),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__3813 (
            .O(N__18974),
            .I(N__18971));
    LocalMux I__3812 (
            .O(N__18971),
            .I(N__18968));
    Odrv4 I__3811 (
            .O(N__18968),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__3810 (
            .O(N__18965),
            .I(N__18962));
    LocalMux I__3809 (
            .O(N__18962),
            .I(N__18959));
    Span4Mux_h I__3808 (
            .O(N__18959),
            .I(N__18956));
    Odrv4 I__3807 (
            .O(N__18956),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__3806 (
            .O(N__18953),
            .I(N__18950));
    LocalMux I__3805 (
            .O(N__18950),
            .I(N__18947));
    Span4Mux_h I__3804 (
            .O(N__18947),
            .I(N__18944));
    Odrv4 I__3803 (
            .O(N__18944),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__3802 (
            .O(N__18941),
            .I(N__18938));
    LocalMux I__3801 (
            .O(N__18938),
            .I(N__18935));
    Span4Mux_v I__3800 (
            .O(N__18935),
            .I(N__18932));
    Odrv4 I__3799 (
            .O(N__18932),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__3798 (
            .O(N__18929),
            .I(N__18926));
    LocalMux I__3797 (
            .O(N__18926),
            .I(N__18923));
    Span4Mux_h I__3796 (
            .O(N__18923),
            .I(N__18920));
    Odrv4 I__3795 (
            .O(N__18920),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__3794 (
            .O(N__18917),
            .I(N__18913));
    InMux I__3793 (
            .O(N__18916),
            .I(N__18910));
    LocalMux I__3792 (
            .O(N__18913),
            .I(N__18907));
    LocalMux I__3791 (
            .O(N__18910),
            .I(N__18904));
    Span4Mux_v I__3790 (
            .O(N__18907),
            .I(N__18901));
    Odrv12 I__3789 (
            .O(N__18904),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    Odrv4 I__3788 (
            .O(N__18901),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__3787 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__3786 (
            .O(N__18893),
            .I(N__18889));
    InMux I__3785 (
            .O(N__18892),
            .I(N__18886));
    Span4Mux_v I__3784 (
            .O(N__18889),
            .I(N__18883));
    LocalMux I__3783 (
            .O(N__18886),
            .I(N__18880));
    Odrv4 I__3782 (
            .O(N__18883),
            .I(scaler_3_data_12));
    Odrv12 I__3781 (
            .O(N__18880),
            .I(scaler_3_data_12));
    InMux I__3780 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__3779 (
            .O(N__18872),
            .I(N__18869));
    Odrv4 I__3778 (
            .O(N__18869),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__3777 (
            .O(N__18866),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    CascadeMux I__3776 (
            .O(N__18863),
            .I(N__18860));
    InMux I__3775 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__3774 (
            .O(N__18857),
            .I(N__18853));
    CascadeMux I__3773 (
            .O(N__18856),
            .I(N__18850));
    Sp12to4 I__3772 (
            .O(N__18853),
            .I(N__18847));
    InMux I__3771 (
            .O(N__18850),
            .I(N__18844));
    Span12Mux_s6_v I__3770 (
            .O(N__18847),
            .I(N__18839));
    LocalMux I__3769 (
            .O(N__18844),
            .I(N__18839));
    Odrv12 I__3768 (
            .O(N__18839),
            .I(scaler_3_data_13));
    InMux I__3767 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__3766 (
            .O(N__18833),
            .I(N__18830));
    Sp12to4 I__3765 (
            .O(N__18830),
            .I(N__18827));
    Odrv12 I__3764 (
            .O(N__18827),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__3763 (
            .O(N__18824),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__3762 (
            .O(N__18821),
            .I(N__18818));
    LocalMux I__3761 (
            .O(N__18818),
            .I(N__18815));
    Span4Mux_v I__3760 (
            .O(N__18815),
            .I(N__18812));
    Odrv4 I__3759 (
            .O(N__18812),
            .I(scaler_3_data_14));
    InMux I__3758 (
            .O(N__18809),
            .I(bfn_11_20_0_));
    InMux I__3757 (
            .O(N__18806),
            .I(N__18803));
    LocalMux I__3756 (
            .O(N__18803),
            .I(N__18800));
    Odrv12 I__3755 (
            .O(N__18800),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    CascadeMux I__3754 (
            .O(N__18797),
            .I(N__18794));
    InMux I__3753 (
            .O(N__18794),
            .I(N__18791));
    LocalMux I__3752 (
            .O(N__18791),
            .I(N__18788));
    Odrv12 I__3751 (
            .O(N__18788),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    CascadeMux I__3750 (
            .O(N__18785),
            .I(N__18782));
    InMux I__3749 (
            .O(N__18782),
            .I(N__18777));
    CascadeMux I__3748 (
            .O(N__18781),
            .I(N__18774));
    CascadeMux I__3747 (
            .O(N__18780),
            .I(N__18770));
    LocalMux I__3746 (
            .O(N__18777),
            .I(N__18762));
    InMux I__3745 (
            .O(N__18774),
            .I(N__18759));
    CascadeMux I__3744 (
            .O(N__18773),
            .I(N__18756));
    InMux I__3743 (
            .O(N__18770),
            .I(N__18753));
    InMux I__3742 (
            .O(N__18769),
            .I(N__18750));
    CascadeMux I__3741 (
            .O(N__18768),
            .I(N__18747));
    CascadeMux I__3740 (
            .O(N__18767),
            .I(N__18743));
    CascadeMux I__3739 (
            .O(N__18766),
            .I(N__18740));
    CascadeMux I__3738 (
            .O(N__18765),
            .I(N__18737));
    Span4Mux_h I__3737 (
            .O(N__18762),
            .I(N__18732));
    LocalMux I__3736 (
            .O(N__18759),
            .I(N__18732));
    InMux I__3735 (
            .O(N__18756),
            .I(N__18729));
    LocalMux I__3734 (
            .O(N__18753),
            .I(N__18726));
    LocalMux I__3733 (
            .O(N__18750),
            .I(N__18723));
    InMux I__3732 (
            .O(N__18747),
            .I(N__18718));
    InMux I__3731 (
            .O(N__18746),
            .I(N__18718));
    InMux I__3730 (
            .O(N__18743),
            .I(N__18715));
    InMux I__3729 (
            .O(N__18740),
            .I(N__18712));
    InMux I__3728 (
            .O(N__18737),
            .I(N__18709));
    Odrv4 I__3727 (
            .O(N__18732),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__3726 (
            .O(N__18729),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__3725 (
            .O(N__18726),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__3724 (
            .O(N__18723),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__3723 (
            .O(N__18718),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__3722 (
            .O(N__18715),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__3721 (
            .O(N__18712),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__3720 (
            .O(N__18709),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    InMux I__3719 (
            .O(N__18692),
            .I(N__18684));
    InMux I__3718 (
            .O(N__18691),
            .I(N__18681));
    InMux I__3717 (
            .O(N__18690),
            .I(N__18678));
    CascadeMux I__3716 (
            .O(N__18689),
            .I(N__18675));
    InMux I__3715 (
            .O(N__18688),
            .I(N__18669));
    InMux I__3714 (
            .O(N__18687),
            .I(N__18666));
    LocalMux I__3713 (
            .O(N__18684),
            .I(N__18660));
    LocalMux I__3712 (
            .O(N__18681),
            .I(N__18660));
    LocalMux I__3711 (
            .O(N__18678),
            .I(N__18657));
    InMux I__3710 (
            .O(N__18675),
            .I(N__18653));
    InMux I__3709 (
            .O(N__18674),
            .I(N__18648));
    InMux I__3708 (
            .O(N__18673),
            .I(N__18648));
    InMux I__3707 (
            .O(N__18672),
            .I(N__18645));
    LocalMux I__3706 (
            .O(N__18669),
            .I(N__18638));
    LocalMux I__3705 (
            .O(N__18666),
            .I(N__18638));
    CascadeMux I__3704 (
            .O(N__18665),
            .I(N__18634));
    Span4Mux_v I__3703 (
            .O(N__18660),
            .I(N__18631));
    Span4Mux_h I__3702 (
            .O(N__18657),
            .I(N__18628));
    InMux I__3701 (
            .O(N__18656),
            .I(N__18625));
    LocalMux I__3700 (
            .O(N__18653),
            .I(N__18620));
    LocalMux I__3699 (
            .O(N__18648),
            .I(N__18620));
    LocalMux I__3698 (
            .O(N__18645),
            .I(N__18617));
    InMux I__3697 (
            .O(N__18644),
            .I(N__18614));
    InMux I__3696 (
            .O(N__18643),
            .I(N__18611));
    Span4Mux_h I__3695 (
            .O(N__18638),
            .I(N__18608));
    InMux I__3694 (
            .O(N__18637),
            .I(N__18603));
    InMux I__3693 (
            .O(N__18634),
            .I(N__18603));
    Odrv4 I__3692 (
            .O(N__18631),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3691 (
            .O(N__18628),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3690 (
            .O(N__18625),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3689 (
            .O(N__18620),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3688 (
            .O(N__18617),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3687 (
            .O(N__18614),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3686 (
            .O(N__18611),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__3685 (
            .O(N__18608),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__3684 (
            .O(N__18603),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    InMux I__3683 (
            .O(N__18584),
            .I(N__18581));
    LocalMux I__3682 (
            .O(N__18581),
            .I(N__18578));
    Span4Mux_v I__3681 (
            .O(N__18578),
            .I(N__18574));
    InMux I__3680 (
            .O(N__18577),
            .I(N__18571));
    Odrv4 I__3679 (
            .O(N__18574),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    LocalMux I__3678 (
            .O(N__18571),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    CascadeMux I__3677 (
            .O(N__18566),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ));
    CascadeMux I__3676 (
            .O(N__18563),
            .I(N__18560));
    InMux I__3675 (
            .O(N__18560),
            .I(N__18557));
    LocalMux I__3674 (
            .O(N__18557),
            .I(N__18554));
    Span4Mux_v I__3673 (
            .O(N__18554),
            .I(N__18551));
    Odrv4 I__3672 (
            .O(N__18551),
            .I(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ));
    CascadeMux I__3671 (
            .O(N__18548),
            .I(N__18545));
    InMux I__3670 (
            .O(N__18545),
            .I(N__18540));
    CascadeMux I__3669 (
            .O(N__18544),
            .I(N__18537));
    CascadeMux I__3668 (
            .O(N__18543),
            .I(N__18532));
    LocalMux I__3667 (
            .O(N__18540),
            .I(N__18527));
    InMux I__3666 (
            .O(N__18537),
            .I(N__18524));
    CascadeMux I__3665 (
            .O(N__18536),
            .I(N__18521));
    InMux I__3664 (
            .O(N__18535),
            .I(N__18518));
    InMux I__3663 (
            .O(N__18532),
            .I(N__18514));
    CascadeMux I__3662 (
            .O(N__18531),
            .I(N__18509));
    CascadeMux I__3661 (
            .O(N__18530),
            .I(N__18506));
    Span4Mux_v I__3660 (
            .O(N__18527),
            .I(N__18500));
    LocalMux I__3659 (
            .O(N__18524),
            .I(N__18500));
    InMux I__3658 (
            .O(N__18521),
            .I(N__18497));
    LocalMux I__3657 (
            .O(N__18518),
            .I(N__18494));
    InMux I__3656 (
            .O(N__18517),
            .I(N__18491));
    LocalMux I__3655 (
            .O(N__18514),
            .I(N__18488));
    InMux I__3654 (
            .O(N__18513),
            .I(N__18483));
    InMux I__3653 (
            .O(N__18512),
            .I(N__18483));
    InMux I__3652 (
            .O(N__18509),
            .I(N__18480));
    InMux I__3651 (
            .O(N__18506),
            .I(N__18477));
    InMux I__3650 (
            .O(N__18505),
            .I(N__18474));
    Odrv4 I__3649 (
            .O(N__18500),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3648 (
            .O(N__18497),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__3647 (
            .O(N__18494),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3646 (
            .O(N__18491),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__3645 (
            .O(N__18488),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3644 (
            .O(N__18483),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3643 (
            .O(N__18480),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3642 (
            .O(N__18477),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__3641 (
            .O(N__18474),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    InMux I__3640 (
            .O(N__18455),
            .I(N__18448));
    InMux I__3639 (
            .O(N__18454),
            .I(N__18445));
    InMux I__3638 (
            .O(N__18453),
            .I(N__18441));
    InMux I__3637 (
            .O(N__18452),
            .I(N__18437));
    CascadeMux I__3636 (
            .O(N__18451),
            .I(N__18432));
    LocalMux I__3635 (
            .O(N__18448),
            .I(N__18424));
    LocalMux I__3634 (
            .O(N__18445),
            .I(N__18424));
    InMux I__3633 (
            .O(N__18444),
            .I(N__18421));
    LocalMux I__3632 (
            .O(N__18441),
            .I(N__18418));
    InMux I__3631 (
            .O(N__18440),
            .I(N__18415));
    LocalMux I__3630 (
            .O(N__18437),
            .I(N__18412));
    InMux I__3629 (
            .O(N__18436),
            .I(N__18409));
    InMux I__3628 (
            .O(N__18435),
            .I(N__18404));
    InMux I__3627 (
            .O(N__18432),
            .I(N__18404));
    InMux I__3626 (
            .O(N__18431),
            .I(N__18401));
    InMux I__3625 (
            .O(N__18430),
            .I(N__18398));
    InMux I__3624 (
            .O(N__18429),
            .I(N__18395));
    Odrv4 I__3623 (
            .O(N__18424),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3622 (
            .O(N__18421),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__3621 (
            .O(N__18418),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3620 (
            .O(N__18415),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__3619 (
            .O(N__18412),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3618 (
            .O(N__18409),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3617 (
            .O(N__18404),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3616 (
            .O(N__18401),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3615 (
            .O(N__18398),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__3614 (
            .O(N__18395),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__3613 (
            .O(N__18374),
            .I(N__18371));
    LocalMux I__3612 (
            .O(N__18371),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    InMux I__3611 (
            .O(N__18368),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__3610 (
            .O(N__18365),
            .I(bfn_11_18_0_));
    InMux I__3609 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__3608 (
            .O(N__18359),
            .I(N__18355));
    InMux I__3607 (
            .O(N__18358),
            .I(N__18352));
    Span4Mux_v I__3606 (
            .O(N__18355),
            .I(N__18347));
    LocalMux I__3605 (
            .O(N__18352),
            .I(N__18347));
    Span4Mux_v I__3604 (
            .O(N__18347),
            .I(N__18344));
    Odrv4 I__3603 (
            .O(N__18344),
            .I(scaler_3_data_6));
    InMux I__3602 (
            .O(N__18341),
            .I(N__18338));
    LocalMux I__3601 (
            .O(N__18338),
            .I(N__18334));
    InMux I__3600 (
            .O(N__18337),
            .I(N__18331));
    Span4Mux_v I__3599 (
            .O(N__18334),
            .I(N__18328));
    LocalMux I__3598 (
            .O(N__18331),
            .I(N__18325));
    Odrv4 I__3597 (
            .O(N__18328),
            .I(scaler_3_data_7));
    Odrv12 I__3596 (
            .O(N__18325),
            .I(scaler_3_data_7));
    CascadeMux I__3595 (
            .O(N__18320),
            .I(N__18317));
    InMux I__3594 (
            .O(N__18317),
            .I(N__18314));
    LocalMux I__3593 (
            .O(N__18314),
            .I(N__18311));
    Span4Mux_v I__3592 (
            .O(N__18311),
            .I(N__18308));
    Odrv4 I__3591 (
            .O(N__18308),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__3590 (
            .O(N__18305),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__3589 (
            .O(N__18302),
            .I(N__18298));
    InMux I__3588 (
            .O(N__18301),
            .I(N__18295));
    LocalMux I__3587 (
            .O(N__18298),
            .I(N__18290));
    LocalMux I__3586 (
            .O(N__18295),
            .I(N__18290));
    Span4Mux_v I__3585 (
            .O(N__18290),
            .I(N__18287));
    Odrv4 I__3584 (
            .O(N__18287),
            .I(scaler_3_data_8));
    InMux I__3583 (
            .O(N__18284),
            .I(N__18281));
    LocalMux I__3582 (
            .O(N__18281),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__3581 (
            .O(N__18278),
            .I(\ppm_encoder_1.un1_elevator_cry_7 ));
    InMux I__3580 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__3579 (
            .O(N__18272),
            .I(N__18269));
    Span4Mux_h I__3578 (
            .O(N__18269),
            .I(N__18265));
    InMux I__3577 (
            .O(N__18268),
            .I(N__18262));
    Span4Mux_v I__3576 (
            .O(N__18265),
            .I(N__18259));
    LocalMux I__3575 (
            .O(N__18262),
            .I(N__18256));
    Odrv4 I__3574 (
            .O(N__18259),
            .I(scaler_3_data_9));
    Odrv12 I__3573 (
            .O(N__18256),
            .I(scaler_3_data_9));
    InMux I__3572 (
            .O(N__18251),
            .I(N__18248));
    LocalMux I__3571 (
            .O(N__18248),
            .I(N__18245));
    Span4Mux_v I__3570 (
            .O(N__18245),
            .I(N__18242));
    Odrv4 I__3569 (
            .O(N__18242),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__3568 (
            .O(N__18239),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__3567 (
            .O(N__18236),
            .I(N__18233));
    LocalMux I__3566 (
            .O(N__18233),
            .I(N__18230));
    Span4Mux_v I__3565 (
            .O(N__18230),
            .I(N__18226));
    InMux I__3564 (
            .O(N__18229),
            .I(N__18223));
    Span4Mux_v I__3563 (
            .O(N__18226),
            .I(N__18220));
    LocalMux I__3562 (
            .O(N__18223),
            .I(N__18217));
    Odrv4 I__3561 (
            .O(N__18220),
            .I(scaler_3_data_10));
    Odrv12 I__3560 (
            .O(N__18217),
            .I(scaler_3_data_10));
    InMux I__3559 (
            .O(N__18212),
            .I(N__18209));
    LocalMux I__3558 (
            .O(N__18209),
            .I(N__18206));
    Span4Mux_v I__3557 (
            .O(N__18206),
            .I(N__18203));
    Odrv4 I__3556 (
            .O(N__18203),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__3555 (
            .O(N__18200),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__3554 (
            .O(N__18197),
            .I(N__18193));
    CascadeMux I__3553 (
            .O(N__18196),
            .I(N__18190));
    LocalMux I__3552 (
            .O(N__18193),
            .I(N__18187));
    InMux I__3551 (
            .O(N__18190),
            .I(N__18184));
    Sp12to4 I__3550 (
            .O(N__18187),
            .I(N__18179));
    LocalMux I__3549 (
            .O(N__18184),
            .I(N__18179));
    Odrv12 I__3548 (
            .O(N__18179),
            .I(scaler_3_data_11));
    InMux I__3547 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__3546 (
            .O(N__18173),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__3545 (
            .O(N__18170),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__3544 (
            .O(N__18167),
            .I(N__18163));
    InMux I__3543 (
            .O(N__18166),
            .I(N__18160));
    LocalMux I__3542 (
            .O(N__18163),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ));
    LocalMux I__3541 (
            .O(N__18160),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ));
    CascadeMux I__3540 (
            .O(N__18155),
            .I(N__18152));
    InMux I__3539 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__3538 (
            .O(N__18149),
            .I(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ));
    InMux I__3537 (
            .O(N__18146),
            .I(bfn_11_16_0_));
    InMux I__3536 (
            .O(N__18143),
            .I(\scaler_3.un2_source_data_0_cry_9 ));
    InMux I__3535 (
            .O(N__18140),
            .I(N__18137));
    LocalMux I__3534 (
            .O(N__18137),
            .I(N__18134));
    Span4Mux_v I__3533 (
            .O(N__18134),
            .I(N__18131));
    Odrv4 I__3532 (
            .O(N__18131),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__3531 (
            .O(N__18128),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__3530 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__3529 (
            .O(N__18122),
            .I(N__18119));
    Odrv4 I__3528 (
            .O(N__18119),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__3527 (
            .O(N__18116),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__3526 (
            .O(N__18113),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__3525 (
            .O(N__18110),
            .I(N__18107));
    LocalMux I__3524 (
            .O(N__18107),
            .I(N__18104));
    Span4Mux_v I__3523 (
            .O(N__18104),
            .I(N__18101));
    Odrv4 I__3522 (
            .O(N__18101),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    InMux I__3521 (
            .O(N__18098),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__3520 (
            .O(N__18095),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__3519 (
            .O(N__18092),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    CascadeMux I__3518 (
            .O(N__18089),
            .I(N__18086));
    InMux I__3517 (
            .O(N__18086),
            .I(N__18083));
    LocalMux I__3516 (
            .O(N__18083),
            .I(N__18080));
    Span4Mux_h I__3515 (
            .O(N__18080),
            .I(N__18077));
    Odrv4 I__3514 (
            .O(N__18077),
            .I(\scaler_3.un2_source_data_0_cry_1_c_RNO_1 ));
    InMux I__3513 (
            .O(N__18074),
            .I(N__18070));
    CascadeMux I__3512 (
            .O(N__18073),
            .I(N__18066));
    LocalMux I__3511 (
            .O(N__18070),
            .I(N__18062));
    InMux I__3510 (
            .O(N__18069),
            .I(N__18059));
    InMux I__3509 (
            .O(N__18066),
            .I(N__18054));
    InMux I__3508 (
            .O(N__18065),
            .I(N__18054));
    Odrv4 I__3507 (
            .O(N__18062),
            .I(\scaler_3.un2_source_data_0 ));
    LocalMux I__3506 (
            .O(N__18059),
            .I(\scaler_3.un2_source_data_0 ));
    LocalMux I__3505 (
            .O(N__18054),
            .I(\scaler_3.un2_source_data_0 ));
    InMux I__3504 (
            .O(N__18047),
            .I(\scaler_3.un2_source_data_0_cry_1 ));
    CascadeMux I__3503 (
            .O(N__18044),
            .I(N__18041));
    InMux I__3502 (
            .O(N__18041),
            .I(N__18035));
    InMux I__3501 (
            .O(N__18040),
            .I(N__18035));
    LocalMux I__3500 (
            .O(N__18035),
            .I(\scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ));
    InMux I__3499 (
            .O(N__18032),
            .I(\scaler_3.un2_source_data_0_cry_2 ));
    CascadeMux I__3498 (
            .O(N__18029),
            .I(N__18026));
    InMux I__3497 (
            .O(N__18026),
            .I(N__18020));
    InMux I__3496 (
            .O(N__18025),
            .I(N__18020));
    LocalMux I__3495 (
            .O(N__18020),
            .I(\scaler_3.un3_source_data_0_cry_2_c_RNIR08I ));
    InMux I__3494 (
            .O(N__18017),
            .I(\scaler_3.un2_source_data_0_cry_3 ));
    CascadeMux I__3493 (
            .O(N__18014),
            .I(N__18011));
    InMux I__3492 (
            .O(N__18011),
            .I(N__18005));
    InMux I__3491 (
            .O(N__18010),
            .I(N__18005));
    LocalMux I__3490 (
            .O(N__18005),
            .I(\scaler_3.un3_source_data_0_cry_3_c_RNIU49I ));
    InMux I__3489 (
            .O(N__18002),
            .I(\scaler_3.un2_source_data_0_cry_4 ));
    CascadeMux I__3488 (
            .O(N__17999),
            .I(N__17996));
    InMux I__3487 (
            .O(N__17996),
            .I(N__17990));
    InMux I__3486 (
            .O(N__17995),
            .I(N__17990));
    LocalMux I__3485 (
            .O(N__17990),
            .I(\scaler_3.un3_source_data_0_cry_4_c_RNI19AI ));
    InMux I__3484 (
            .O(N__17987),
            .I(\scaler_3.un2_source_data_0_cry_5 ));
    CascadeMux I__3483 (
            .O(N__17984),
            .I(N__17981));
    InMux I__3482 (
            .O(N__17981),
            .I(N__17975));
    InMux I__3481 (
            .O(N__17980),
            .I(N__17975));
    LocalMux I__3480 (
            .O(N__17975),
            .I(\scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ));
    InMux I__3479 (
            .O(N__17972),
            .I(\scaler_3.un2_source_data_0_cry_6 ));
    CascadeMux I__3478 (
            .O(N__17969),
            .I(N__17966));
    InMux I__3477 (
            .O(N__17966),
            .I(N__17960));
    InMux I__3476 (
            .O(N__17965),
            .I(N__17960));
    LocalMux I__3475 (
            .O(N__17960),
            .I(\scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ));
    InMux I__3474 (
            .O(N__17957),
            .I(\scaler_3.un2_source_data_0_cry_7 ));
    InMux I__3473 (
            .O(N__17954),
            .I(bfn_11_13_0_));
    InMux I__3472 (
            .O(N__17951),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CEMux I__3471 (
            .O(N__17948),
            .I(N__17945));
    LocalMux I__3470 (
            .O(N__17945),
            .I(N__17942));
    Sp12to4 I__3469 (
            .O(N__17942),
            .I(N__17939));
    Odrv12 I__3468 (
            .O(N__17939),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__3467 (
            .O(N__17936),
            .I(N__17932));
    InMux I__3466 (
            .O(N__17935),
            .I(N__17929));
    LocalMux I__3465 (
            .O(N__17932),
            .I(N__17926));
    LocalMux I__3464 (
            .O(N__17929),
            .I(N__17922));
    Span4Mux_h I__3463 (
            .O(N__17926),
            .I(N__17919));
    InMux I__3462 (
            .O(N__17925),
            .I(N__17916));
    Span4Mux_v I__3461 (
            .O(N__17922),
            .I(N__17908));
    Span4Mux_v I__3460 (
            .O(N__17919),
            .I(N__17908));
    LocalMux I__3459 (
            .O(N__17916),
            .I(N__17908));
    InMux I__3458 (
            .O(N__17915),
            .I(N__17905));
    Odrv4 I__3457 (
            .O(N__17908),
            .I(frame_decoder_CH4data_0));
    LocalMux I__3456 (
            .O(N__17905),
            .I(frame_decoder_CH4data_0));
    InMux I__3455 (
            .O(N__17900),
            .I(N__17897));
    LocalMux I__3454 (
            .O(N__17897),
            .I(N__17892));
    InMux I__3453 (
            .O(N__17896),
            .I(N__17889));
    CascadeMux I__3452 (
            .O(N__17895),
            .I(N__17885));
    Span4Mux_v I__3451 (
            .O(N__17892),
            .I(N__17880));
    LocalMux I__3450 (
            .O(N__17889),
            .I(N__17880));
    InMux I__3449 (
            .O(N__17888),
            .I(N__17877));
    InMux I__3448 (
            .O(N__17885),
            .I(N__17874));
    Odrv4 I__3447 (
            .O(N__17880),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__3446 (
            .O(N__17877),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__3445 (
            .O(N__17874),
            .I(frame_decoder_OFF4data_0));
    InMux I__3444 (
            .O(N__17867),
            .I(N__17864));
    LocalMux I__3443 (
            .O(N__17864),
            .I(\scaler_4.N_544_i_l_ofxZ0 ));
    InMux I__3442 (
            .O(N__17861),
            .I(N__17857));
    InMux I__3441 (
            .O(N__17860),
            .I(N__17854));
    LocalMux I__3440 (
            .O(N__17857),
            .I(N__17851));
    LocalMux I__3439 (
            .O(N__17854),
            .I(frame_decoder_OFF2data_7));
    Odrv4 I__3438 (
            .O(N__17851),
            .I(frame_decoder_OFF2data_7));
    InMux I__3437 (
            .O(N__17846),
            .I(N__17843));
    LocalMux I__3436 (
            .O(N__17843),
            .I(N__17840));
    Odrv4 I__3435 (
            .O(N__17840),
            .I(\scaler_2.un3_source_data_0_axb_7 ));
    InMux I__3434 (
            .O(N__17837),
            .I(N__17834));
    LocalMux I__3433 (
            .O(N__17834),
            .I(N__17831));
    Span4Mux_h I__3432 (
            .O(N__17831),
            .I(N__17827));
    InMux I__3431 (
            .O(N__17830),
            .I(N__17824));
    Odrv4 I__3430 (
            .O(N__17827),
            .I(frame_decoder_CH2data_7));
    LocalMux I__3429 (
            .O(N__17824),
            .I(frame_decoder_CH2data_7));
    CEMux I__3428 (
            .O(N__17819),
            .I(N__17816));
    LocalMux I__3427 (
            .O(N__17816),
            .I(N__17812));
    CEMux I__3426 (
            .O(N__17815),
            .I(N__17809));
    Span4Mux_h I__3425 (
            .O(N__17812),
            .I(N__17806));
    LocalMux I__3424 (
            .O(N__17809),
            .I(N__17803));
    Odrv4 I__3423 (
            .O(N__17806),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    Odrv12 I__3422 (
            .O(N__17803),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__3421 (
            .O(N__17798),
            .I(N__17795));
    LocalMux I__3420 (
            .O(N__17795),
            .I(N__17791));
    InMux I__3419 (
            .O(N__17794),
            .I(N__17788));
    Span4Mux_h I__3418 (
            .O(N__17791),
            .I(N__17785));
    LocalMux I__3417 (
            .O(N__17788),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    Odrv4 I__3416 (
            .O(N__17785),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    InMux I__3415 (
            .O(N__17780),
            .I(N__17777));
    LocalMux I__3414 (
            .O(N__17777),
            .I(N__17774));
    Span4Mux_v I__3413 (
            .O(N__17774),
            .I(N__17770));
    InMux I__3412 (
            .O(N__17773),
            .I(N__17767));
    Odrv4 I__3411 (
            .O(N__17770),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa ));
    LocalMux I__3410 (
            .O(N__17767),
            .I(\uart_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__3409 (
            .O(N__17762),
            .I(N__17758));
    InMux I__3408 (
            .O(N__17761),
            .I(N__17755));
    LocalMux I__3407 (
            .O(N__17758),
            .I(N__17752));
    LocalMux I__3406 (
            .O(N__17755),
            .I(frame_decoder_OFF4data_7));
    Odrv4 I__3405 (
            .O(N__17752),
            .I(frame_decoder_OFF4data_7));
    InMux I__3404 (
            .O(N__17747),
            .I(N__17743));
    InMux I__3403 (
            .O(N__17746),
            .I(N__17740));
    LocalMux I__3402 (
            .O(N__17743),
            .I(N__17735));
    LocalMux I__3401 (
            .O(N__17740),
            .I(N__17735));
    Odrv4 I__3400 (
            .O(N__17735),
            .I(frame_decoder_CH4data_7));
    InMux I__3399 (
            .O(N__17732),
            .I(N__17729));
    LocalMux I__3398 (
            .O(N__17729),
            .I(N__17726));
    Odrv4 I__3397 (
            .O(N__17726),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__3396 (
            .O(N__17723),
            .I(N__17720));
    LocalMux I__3395 (
            .O(N__17720),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__3394 (
            .O(N__17717),
            .I(N__17714));
    InMux I__3393 (
            .O(N__17714),
            .I(N__17711));
    LocalMux I__3392 (
            .O(N__17711),
            .I(frame_decoder_OFF4data_1));
    InMux I__3391 (
            .O(N__17708),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__3390 (
            .O(N__17705),
            .I(N__17702));
    LocalMux I__3389 (
            .O(N__17702),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__3388 (
            .O(N__17699),
            .I(N__17696));
    InMux I__3387 (
            .O(N__17696),
            .I(N__17693));
    LocalMux I__3386 (
            .O(N__17693),
            .I(frame_decoder_OFF4data_2));
    InMux I__3385 (
            .O(N__17690),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__3384 (
            .O(N__17687),
            .I(N__17684));
    LocalMux I__3383 (
            .O(N__17684),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__3382 (
            .O(N__17681),
            .I(N__17678));
    InMux I__3381 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__3380 (
            .O(N__17675),
            .I(frame_decoder_OFF4data_3));
    InMux I__3379 (
            .O(N__17672),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__3378 (
            .O(N__17669),
            .I(N__17666));
    LocalMux I__3377 (
            .O(N__17666),
            .I(frame_decoder_CH4data_4));
    InMux I__3376 (
            .O(N__17663),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__3375 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__3374 (
            .O(N__17657),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__3373 (
            .O(N__17654),
            .I(N__17651));
    InMux I__3372 (
            .O(N__17651),
            .I(N__17648));
    LocalMux I__3371 (
            .O(N__17648),
            .I(frame_decoder_OFF4data_5));
    InMux I__3370 (
            .O(N__17645),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__3369 (
            .O(N__17642),
            .I(N__17639));
    LocalMux I__3368 (
            .O(N__17639),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__3367 (
            .O(N__17636),
            .I(N__17633));
    InMux I__3366 (
            .O(N__17633),
            .I(N__17630));
    LocalMux I__3365 (
            .O(N__17630),
            .I(frame_decoder_OFF4data_6));
    InMux I__3364 (
            .O(N__17627),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__3363 (
            .O(N__17624),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__3362 (
            .O(N__17621),
            .I(N__17618));
    LocalMux I__3361 (
            .O(N__17618),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__3360 (
            .O(N__17615),
            .I(N__17612));
    LocalMux I__3359 (
            .O(N__17612),
            .I(N__17609));
    Odrv4 I__3358 (
            .O(N__17609),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__3357 (
            .O(N__17606),
            .I(N__17603));
    LocalMux I__3356 (
            .O(N__17603),
            .I(N__17600));
    Span4Mux_s3_v I__3355 (
            .O(N__17600),
            .I(N__17597));
    Span4Mux_v I__3354 (
            .O(N__17597),
            .I(N__17594));
    Odrv4 I__3353 (
            .O(N__17594),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    CascadeMux I__3352 (
            .O(N__17591),
            .I(N__17588));
    InMux I__3351 (
            .O(N__17588),
            .I(N__17585));
    LocalMux I__3350 (
            .O(N__17585),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__3349 (
            .O(N__17582),
            .I(N__17579));
    LocalMux I__3348 (
            .O(N__17579),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__3347 (
            .O(N__17576),
            .I(N__17573));
    LocalMux I__3346 (
            .O(N__17573),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__3345 (
            .O(N__17570),
            .I(N__17567));
    LocalMux I__3344 (
            .O(N__17567),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__3343 (
            .O(N__17564),
            .I(N__17560));
    InMux I__3342 (
            .O(N__17563),
            .I(N__17557));
    LocalMux I__3341 (
            .O(N__17560),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    LocalMux I__3340 (
            .O(N__17557),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    CascadeMux I__3339 (
            .O(N__17552),
            .I(N__17548));
    InMux I__3338 (
            .O(N__17551),
            .I(N__17545));
    InMux I__3337 (
            .O(N__17548),
            .I(N__17542));
    LocalMux I__3336 (
            .O(N__17545),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    LocalMux I__3335 (
            .O(N__17542),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__3334 (
            .O(N__17537),
            .I(N__17534));
    LocalMux I__3333 (
            .O(N__17534),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__3332 (
            .O(N__17531),
            .I(N__17527));
    InMux I__3331 (
            .O(N__17530),
            .I(N__17524));
    LocalMux I__3330 (
            .O(N__17527),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    LocalMux I__3329 (
            .O(N__17524),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    CascadeMux I__3328 (
            .O(N__17519),
            .I(N__17516));
    InMux I__3327 (
            .O(N__17516),
            .I(N__17513));
    LocalMux I__3326 (
            .O(N__17513),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__3325 (
            .O(N__17510),
            .I(N__17507));
    LocalMux I__3324 (
            .O(N__17507),
            .I(N__17504));
    Span4Mux_s2_v I__3323 (
            .O(N__17504),
            .I(N__17501));
    Span4Mux_v I__3322 (
            .O(N__17501),
            .I(N__17498));
    Odrv4 I__3321 (
            .O(N__17498),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__3320 (
            .O(N__17495),
            .I(N__17492));
    LocalMux I__3319 (
            .O(N__17492),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    InMux I__3318 (
            .O(N__17489),
            .I(N__17486));
    LocalMux I__3317 (
            .O(N__17486),
            .I(N__17483));
    Span4Mux_s3_v I__3316 (
            .O(N__17483),
            .I(N__17480));
    Odrv4 I__3315 (
            .O(N__17480),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__3314 (
            .O(N__17477),
            .I(N__17474));
    LocalMux I__3313 (
            .O(N__17474),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__3312 (
            .O(N__17471),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__3311 (
            .O(N__17468),
            .I(N__17465));
    LocalMux I__3310 (
            .O(N__17465),
            .I(N__17462));
    Span4Mux_s3_v I__3309 (
            .O(N__17462),
            .I(N__17459));
    Span4Mux_v I__3308 (
            .O(N__17459),
            .I(N__17456));
    Odrv4 I__3307 (
            .O(N__17456),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__3306 (
            .O(N__17453),
            .I(N__17450));
    InMux I__3305 (
            .O(N__17450),
            .I(N__17447));
    LocalMux I__3304 (
            .O(N__17447),
            .I(N__17444));
    Odrv12 I__3303 (
            .O(N__17444),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__3302 (
            .O(N__17441),
            .I(N__17438));
    LocalMux I__3301 (
            .O(N__17438),
            .I(N__17435));
    Span4Mux_v I__3300 (
            .O(N__17435),
            .I(N__17432));
    Odrv4 I__3299 (
            .O(N__17432),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__3298 (
            .O(N__17429),
            .I(N__17426));
    LocalMux I__3297 (
            .O(N__17426),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__3296 (
            .O(N__17423),
            .I(N__17420));
    LocalMux I__3295 (
            .O(N__17420),
            .I(N__17416));
    InMux I__3294 (
            .O(N__17419),
            .I(N__17413));
    Sp12to4 I__3293 (
            .O(N__17416),
            .I(N__17410));
    LocalMux I__3292 (
            .O(N__17413),
            .I(N__17407));
    Odrv12 I__3291 (
            .O(N__17410),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    Odrv4 I__3290 (
            .O(N__17407),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    InMux I__3289 (
            .O(N__17402),
            .I(N__17399));
    LocalMux I__3288 (
            .O(N__17399),
            .I(N__17396));
    Span4Mux_h I__3287 (
            .O(N__17396),
            .I(N__17393));
    Odrv4 I__3286 (
            .O(N__17393),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__3285 (
            .O(N__17390),
            .I(N__17387));
    LocalMux I__3284 (
            .O(N__17387),
            .I(N__17384));
    Span4Mux_v I__3283 (
            .O(N__17384),
            .I(N__17381));
    Odrv4 I__3282 (
            .O(N__17381),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__3281 (
            .O(N__17378),
            .I(N__17375));
    LocalMux I__3280 (
            .O(N__17375),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__3279 (
            .O(N__17372),
            .I(N__17369));
    LocalMux I__3278 (
            .O(N__17369),
            .I(N__17366));
    Span4Mux_v I__3277 (
            .O(N__17366),
            .I(N__17362));
    InMux I__3276 (
            .O(N__17365),
            .I(N__17359));
    Odrv4 I__3275 (
            .O(N__17362),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    LocalMux I__3274 (
            .O(N__17359),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    InMux I__3273 (
            .O(N__17354),
            .I(N__17351));
    LocalMux I__3272 (
            .O(N__17351),
            .I(N__17348));
    Span4Mux_h I__3271 (
            .O(N__17348),
            .I(N__17345));
    Odrv4 I__3270 (
            .O(N__17345),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    CascadeMux I__3269 (
            .O(N__17342),
            .I(\ppm_encoder_1.N_305_cascade_ ));
    InMux I__3268 (
            .O(N__17339),
            .I(N__17330));
    InMux I__3267 (
            .O(N__17338),
            .I(N__17330));
    InMux I__3266 (
            .O(N__17337),
            .I(N__17330));
    LocalMux I__3265 (
            .O(N__17330),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__3264 (
            .O(N__17327),
            .I(N__17318));
    InMux I__3263 (
            .O(N__17326),
            .I(N__17318));
    InMux I__3262 (
            .O(N__17325),
            .I(N__17318));
    LocalMux I__3261 (
            .O(N__17318),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__3260 (
            .O(N__17315),
            .I(N__17311));
    InMux I__3259 (
            .O(N__17314),
            .I(N__17308));
    LocalMux I__3258 (
            .O(N__17311),
            .I(N__17303));
    LocalMux I__3257 (
            .O(N__17308),
            .I(N__17303));
    Odrv12 I__3256 (
            .O(N__17303),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    CascadeMux I__3255 (
            .O(N__17300),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ));
    CascadeMux I__3254 (
            .O(N__17297),
            .I(N__17294));
    InMux I__3253 (
            .O(N__17294),
            .I(N__17291));
    LocalMux I__3252 (
            .O(N__17291),
            .I(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ));
    InMux I__3251 (
            .O(N__17288),
            .I(N__17285));
    LocalMux I__3250 (
            .O(N__17285),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13 ));
    CascadeMux I__3249 (
            .O(N__17282),
            .I(\ppm_encoder_1.N_308_cascade_ ));
    InMux I__3248 (
            .O(N__17279),
            .I(N__17270));
    InMux I__3247 (
            .O(N__17278),
            .I(N__17270));
    InMux I__3246 (
            .O(N__17277),
            .I(N__17270));
    LocalMux I__3245 (
            .O(N__17270),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__3244 (
            .O(N__17267),
            .I(N__17258));
    InMux I__3243 (
            .O(N__17266),
            .I(N__17258));
    InMux I__3242 (
            .O(N__17265),
            .I(N__17258));
    LocalMux I__3241 (
            .O(N__17258),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    InMux I__3240 (
            .O(N__17255),
            .I(N__17252));
    LocalMux I__3239 (
            .O(N__17252),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    InMux I__3238 (
            .O(N__17249),
            .I(N__17240));
    InMux I__3237 (
            .O(N__17248),
            .I(N__17240));
    InMux I__3236 (
            .O(N__17247),
            .I(N__17240));
    LocalMux I__3235 (
            .O(N__17240),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__3234 (
            .O(N__17237),
            .I(N__17228));
    InMux I__3233 (
            .O(N__17236),
            .I(N__17228));
    InMux I__3232 (
            .O(N__17235),
            .I(N__17228));
    LocalMux I__3231 (
            .O(N__17228),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    InMux I__3230 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__3229 (
            .O(N__17222),
            .I(N__17218));
    InMux I__3228 (
            .O(N__17221),
            .I(N__17215));
    Span4Mux_h I__3227 (
            .O(N__17218),
            .I(N__17210));
    LocalMux I__3226 (
            .O(N__17215),
            .I(N__17210));
    Odrv4 I__3225 (
            .O(N__17210),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    CascadeMux I__3224 (
            .O(N__17207),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ));
    CascadeMux I__3223 (
            .O(N__17204),
            .I(N__17201));
    InMux I__3222 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__3221 (
            .O(N__17198),
            .I(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ));
    InMux I__3220 (
            .O(N__17195),
            .I(N__17192));
    LocalMux I__3219 (
            .O(N__17192),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10 ));
    InMux I__3218 (
            .O(N__17189),
            .I(N__17185));
    CascadeMux I__3217 (
            .O(N__17188),
            .I(N__17182));
    LocalMux I__3216 (
            .O(N__17185),
            .I(N__17179));
    InMux I__3215 (
            .O(N__17182),
            .I(N__17176));
    Span4Mux_v I__3214 (
            .O(N__17179),
            .I(N__17171));
    LocalMux I__3213 (
            .O(N__17176),
            .I(N__17171));
    Span4Mux_h I__3212 (
            .O(N__17171),
            .I(N__17168));
    Odrv4 I__3211 (
            .O(N__17168),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    CascadeMux I__3210 (
            .O(N__17165),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    InMux I__3209 (
            .O(N__17162),
            .I(N__17159));
    LocalMux I__3208 (
            .O(N__17159),
            .I(N__17156));
    Odrv4 I__3207 (
            .O(N__17156),
            .I(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ));
    InMux I__3206 (
            .O(N__17153),
            .I(N__17150));
    LocalMux I__3205 (
            .O(N__17150),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    CascadeMux I__3204 (
            .O(N__17147),
            .I(N__17142));
    InMux I__3203 (
            .O(N__17146),
            .I(N__17137));
    InMux I__3202 (
            .O(N__17145),
            .I(N__17137));
    InMux I__3201 (
            .O(N__17142),
            .I(N__17134));
    LocalMux I__3200 (
            .O(N__17137),
            .I(N__17131));
    LocalMux I__3199 (
            .O(N__17134),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    Odrv4 I__3198 (
            .O(N__17131),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__3197 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__3196 (
            .O(N__17123),
            .I(N__17120));
    Odrv4 I__3195 (
            .O(N__17120),
            .I(\ppm_encoder_1.N_302 ));
    InMux I__3194 (
            .O(N__17117),
            .I(N__17112));
    InMux I__3193 (
            .O(N__17116),
            .I(N__17107));
    InMux I__3192 (
            .O(N__17115),
            .I(N__17107));
    LocalMux I__3191 (
            .O(N__17112),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    LocalMux I__3190 (
            .O(N__17107),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__3189 (
            .O(N__17102),
            .I(N__17099));
    LocalMux I__3188 (
            .O(N__17099),
            .I(N__17094));
    InMux I__3187 (
            .O(N__17098),
            .I(N__17089));
    InMux I__3186 (
            .O(N__17097),
            .I(N__17089));
    Odrv4 I__3185 (
            .O(N__17094),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    LocalMux I__3184 (
            .O(N__17089),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__3183 (
            .O(N__17084),
            .I(N__17080));
    InMux I__3182 (
            .O(N__17083),
            .I(N__17077));
    LocalMux I__3181 (
            .O(N__17080),
            .I(N__17074));
    LocalMux I__3180 (
            .O(N__17077),
            .I(N__17071));
    Span4Mux_v I__3179 (
            .O(N__17074),
            .I(N__17068));
    Span4Mux_h I__3178 (
            .O(N__17071),
            .I(N__17065));
    Odrv4 I__3177 (
            .O(N__17068),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    Odrv4 I__3176 (
            .O(N__17065),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    CascadeMux I__3175 (
            .O(N__17060),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    CascadeMux I__3174 (
            .O(N__17057),
            .I(N__17054));
    InMux I__3173 (
            .O(N__17054),
            .I(N__17051));
    LocalMux I__3172 (
            .O(N__17051),
            .I(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ));
    CascadeMux I__3171 (
            .O(N__17048),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__3170 (
            .O(N__17045),
            .I(N__17042));
    LocalMux I__3169 (
            .O(N__17042),
            .I(N__17039));
    Span4Mux_h I__3168 (
            .O(N__17039),
            .I(N__17035));
    InMux I__3167 (
            .O(N__17038),
            .I(N__17032));
    Odrv4 I__3166 (
            .O(N__17035),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    LocalMux I__3165 (
            .O(N__17032),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    CascadeMux I__3164 (
            .O(N__17027),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    CascadeMux I__3163 (
            .O(N__17024),
            .I(N__17021));
    InMux I__3162 (
            .O(N__17021),
            .I(N__17018));
    LocalMux I__3161 (
            .O(N__17018),
            .I(N__17015));
    Span4Mux_v I__3160 (
            .O(N__17015),
            .I(N__17012));
    Odrv4 I__3159 (
            .O(N__17012),
            .I(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ));
    InMux I__3158 (
            .O(N__17009),
            .I(N__17006));
    LocalMux I__3157 (
            .O(N__17006),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    InMux I__3156 (
            .O(N__17003),
            .I(N__17000));
    LocalMux I__3155 (
            .O(N__17000),
            .I(N__16997));
    Odrv4 I__3154 (
            .O(N__16997),
            .I(\ppm_encoder_1.N_307 ));
    InMux I__3153 (
            .O(N__16994),
            .I(N__16985));
    InMux I__3152 (
            .O(N__16993),
            .I(N__16985));
    InMux I__3151 (
            .O(N__16992),
            .I(N__16985));
    LocalMux I__3150 (
            .O(N__16985),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__3149 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__3148 (
            .O(N__16979),
            .I(N__16976));
    Span4Mux_h I__3147 (
            .O(N__16976),
            .I(N__16971));
    InMux I__3146 (
            .O(N__16975),
            .I(N__16966));
    InMux I__3145 (
            .O(N__16974),
            .I(N__16966));
    Odrv4 I__3144 (
            .O(N__16971),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    LocalMux I__3143 (
            .O(N__16966),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    CascadeMux I__3142 (
            .O(N__16961),
            .I(N__16957));
    InMux I__3141 (
            .O(N__16960),
            .I(N__16954));
    InMux I__3140 (
            .O(N__16957),
            .I(N__16950));
    LocalMux I__3139 (
            .O(N__16954),
            .I(N__16947));
    InMux I__3138 (
            .O(N__16953),
            .I(N__16944));
    LocalMux I__3137 (
            .O(N__16950),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__3136 (
            .O(N__16947),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    LocalMux I__3135 (
            .O(N__16944),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    InMux I__3134 (
            .O(N__16937),
            .I(N__16930));
    InMux I__3133 (
            .O(N__16936),
            .I(N__16930));
    InMux I__3132 (
            .O(N__16935),
            .I(N__16927));
    LocalMux I__3131 (
            .O(N__16930),
            .I(N__16924));
    LocalMux I__3130 (
            .O(N__16927),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__3129 (
            .O(N__16924),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__3128 (
            .O(N__16919),
            .I(N__16914));
    InMux I__3127 (
            .O(N__16918),
            .I(N__16909));
    InMux I__3126 (
            .O(N__16917),
            .I(N__16909));
    LocalMux I__3125 (
            .O(N__16914),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__3124 (
            .O(N__16909),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    CascadeMux I__3123 (
            .O(N__16904),
            .I(N__16900));
    InMux I__3122 (
            .O(N__16903),
            .I(N__16896));
    InMux I__3121 (
            .O(N__16900),
            .I(N__16893));
    InMux I__3120 (
            .O(N__16899),
            .I(N__16890));
    LocalMux I__3119 (
            .O(N__16896),
            .I(N__16887));
    LocalMux I__3118 (
            .O(N__16893),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__3117 (
            .O(N__16890),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__3116 (
            .O(N__16887),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__3115 (
            .O(N__16880),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ));
    CascadeMux I__3114 (
            .O(N__16877),
            .I(N__16873));
    InMux I__3113 (
            .O(N__16876),
            .I(N__16869));
    InMux I__3112 (
            .O(N__16873),
            .I(N__16866));
    InMux I__3111 (
            .O(N__16872),
            .I(N__16863));
    LocalMux I__3110 (
            .O(N__16869),
            .I(N__16860));
    LocalMux I__3109 (
            .O(N__16866),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    LocalMux I__3108 (
            .O(N__16863),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__3107 (
            .O(N__16860),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    CascadeMux I__3106 (
            .O(N__16853),
            .I(\ppm_encoder_1.N_303_cascade_ ));
    CascadeMux I__3105 (
            .O(N__16850),
            .I(N__16846));
    InMux I__3104 (
            .O(N__16849),
            .I(N__16842));
    InMux I__3103 (
            .O(N__16846),
            .I(N__16839));
    InMux I__3102 (
            .O(N__16845),
            .I(N__16836));
    LocalMux I__3101 (
            .O(N__16842),
            .I(N__16833));
    LocalMux I__3100 (
            .O(N__16839),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__3099 (
            .O(N__16836),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    Odrv4 I__3098 (
            .O(N__16833),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__3097 (
            .O(N__16826),
            .I(N__16823));
    InMux I__3096 (
            .O(N__16823),
            .I(N__16817));
    InMux I__3095 (
            .O(N__16822),
            .I(N__16817));
    LocalMux I__3094 (
            .O(N__16817),
            .I(N__16814));
    Odrv4 I__3093 (
            .O(N__16814),
            .I(\scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ));
    InMux I__3092 (
            .O(N__16811),
            .I(\scaler_1.un2_source_data_0_cry_3 ));
    CascadeMux I__3091 (
            .O(N__16808),
            .I(N__16805));
    InMux I__3090 (
            .O(N__16805),
            .I(N__16799));
    InMux I__3089 (
            .O(N__16804),
            .I(N__16799));
    LocalMux I__3088 (
            .O(N__16799),
            .I(N__16796));
    Odrv4 I__3087 (
            .O(N__16796),
            .I(\scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ));
    InMux I__3086 (
            .O(N__16793),
            .I(\scaler_1.un2_source_data_0_cry_4 ));
    CascadeMux I__3085 (
            .O(N__16790),
            .I(N__16787));
    InMux I__3084 (
            .O(N__16787),
            .I(N__16781));
    InMux I__3083 (
            .O(N__16786),
            .I(N__16781));
    LocalMux I__3082 (
            .O(N__16781),
            .I(N__16778));
    Odrv12 I__3081 (
            .O(N__16778),
            .I(\scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ));
    InMux I__3080 (
            .O(N__16775),
            .I(\scaler_1.un2_source_data_0_cry_5 ));
    CascadeMux I__3079 (
            .O(N__16772),
            .I(N__16769));
    InMux I__3078 (
            .O(N__16769),
            .I(N__16763));
    InMux I__3077 (
            .O(N__16768),
            .I(N__16763));
    LocalMux I__3076 (
            .O(N__16763),
            .I(N__16760));
    Odrv12 I__3075 (
            .O(N__16760),
            .I(\scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ));
    InMux I__3074 (
            .O(N__16757),
            .I(\scaler_1.un2_source_data_0_cry_6 ));
    CascadeMux I__3073 (
            .O(N__16754),
            .I(N__16751));
    InMux I__3072 (
            .O(N__16751),
            .I(N__16745));
    InMux I__3071 (
            .O(N__16750),
            .I(N__16745));
    LocalMux I__3070 (
            .O(N__16745),
            .I(N__16742));
    Odrv12 I__3069 (
            .O(N__16742),
            .I(\scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ));
    InMux I__3068 (
            .O(N__16739),
            .I(\scaler_1.un2_source_data_0_cry_7 ));
    InMux I__3067 (
            .O(N__16736),
            .I(N__16732));
    InMux I__3066 (
            .O(N__16735),
            .I(N__16729));
    LocalMux I__3065 (
            .O(N__16732),
            .I(N__16724));
    LocalMux I__3064 (
            .O(N__16729),
            .I(N__16724));
    Span4Mux_v I__3063 (
            .O(N__16724),
            .I(N__16721));
    Odrv4 I__3062 (
            .O(N__16721),
            .I(\scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ));
    CascadeMux I__3061 (
            .O(N__16718),
            .I(N__16715));
    InMux I__3060 (
            .O(N__16715),
            .I(N__16712));
    LocalMux I__3059 (
            .O(N__16712),
            .I(N__16709));
    Odrv4 I__3058 (
            .O(N__16709),
            .I(\scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ));
    InMux I__3057 (
            .O(N__16706),
            .I(bfn_10_18_0_));
    InMux I__3056 (
            .O(N__16703),
            .I(\scaler_1.un2_source_data_0_cry_9 ));
    InMux I__3055 (
            .O(N__16700),
            .I(bfn_10_16_0_));
    InMux I__3054 (
            .O(N__16697),
            .I(\scaler_3.un3_source_data_0_cry_8 ));
    InMux I__3053 (
            .O(N__16694),
            .I(N__16691));
    LocalMux I__3052 (
            .O(N__16691),
            .I(N__16687));
    InMux I__3051 (
            .O(N__16690),
            .I(N__16684));
    Span4Mux_h I__3050 (
            .O(N__16687),
            .I(N__16681));
    LocalMux I__3049 (
            .O(N__16684),
            .I(\uart_frame_decoder.count8_0_i ));
    Odrv4 I__3048 (
            .O(N__16681),
            .I(\uart_frame_decoder.count8_0_i ));
    InMux I__3047 (
            .O(N__16676),
            .I(N__16673));
    LocalMux I__3046 (
            .O(N__16673),
            .I(N__16670));
    Span4Mux_h I__3045 (
            .O(N__16670),
            .I(N__16666));
    InMux I__3044 (
            .O(N__16669),
            .I(N__16663));
    Odrv4 I__3043 (
            .O(N__16666),
            .I(frame_decoder_OFF3data_7));
    LocalMux I__3042 (
            .O(N__16663),
            .I(frame_decoder_OFF3data_7));
    InMux I__3041 (
            .O(N__16658),
            .I(N__16655));
    LocalMux I__3040 (
            .O(N__16655),
            .I(\scaler_3.N_532_i_l_ofxZ0 ));
    InMux I__3039 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__3038 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_v I__3037 (
            .O(N__16646),
            .I(N__16643));
    Odrv4 I__3036 (
            .O(N__16643),
            .I(\uart_frame_decoder.state_1_RNINMHJZ0Z_10 ));
    InMux I__3035 (
            .O(N__16640),
            .I(N__16637));
    LocalMux I__3034 (
            .O(N__16637),
            .I(N__16632));
    InMux I__3033 (
            .O(N__16636),
            .I(N__16627));
    InMux I__3032 (
            .O(N__16635),
            .I(N__16627));
    Odrv4 I__3031 (
            .O(N__16632),
            .I(\uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61 ));
    LocalMux I__3030 (
            .O(N__16627),
            .I(\uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61 ));
    InMux I__3029 (
            .O(N__16622),
            .I(N__16619));
    LocalMux I__3028 (
            .O(N__16619),
            .I(N__16615));
    InMux I__3027 (
            .O(N__16618),
            .I(N__16612));
    Span4Mux_h I__3026 (
            .O(N__16615),
            .I(N__16607));
    LocalMux I__3025 (
            .O(N__16612),
            .I(N__16604));
    InMux I__3024 (
            .O(N__16611),
            .I(N__16599));
    InMux I__3023 (
            .O(N__16610),
            .I(N__16599));
    Odrv4 I__3022 (
            .O(N__16607),
            .I(\uart_frame_decoder.count8_0 ));
    Odrv4 I__3021 (
            .O(N__16604),
            .I(\uart_frame_decoder.count8_0 ));
    LocalMux I__3020 (
            .O(N__16599),
            .I(\uart_frame_decoder.count8_0 ));
    InMux I__3019 (
            .O(N__16592),
            .I(N__16588));
    InMux I__3018 (
            .O(N__16591),
            .I(N__16584));
    LocalMux I__3017 (
            .O(N__16588),
            .I(N__16580));
    InMux I__3016 (
            .O(N__16587),
            .I(N__16577));
    LocalMux I__3015 (
            .O(N__16584),
            .I(N__16574));
    CascadeMux I__3014 (
            .O(N__16583),
            .I(N__16571));
    Span4Mux_v I__3013 (
            .O(N__16580),
            .I(N__16564));
    LocalMux I__3012 (
            .O(N__16577),
            .I(N__16564));
    Span4Mux_v I__3011 (
            .O(N__16574),
            .I(N__16564));
    InMux I__3010 (
            .O(N__16571),
            .I(N__16561));
    Odrv4 I__3009 (
            .O(N__16564),
            .I(frame_decoder_OFF1data_0));
    LocalMux I__3008 (
            .O(N__16561),
            .I(frame_decoder_OFF1data_0));
    InMux I__3007 (
            .O(N__16556),
            .I(N__16551));
    InMux I__3006 (
            .O(N__16555),
            .I(N__16548));
    InMux I__3005 (
            .O(N__16554),
            .I(N__16545));
    LocalMux I__3004 (
            .O(N__16551),
            .I(N__16542));
    LocalMux I__3003 (
            .O(N__16548),
            .I(N__16537));
    LocalMux I__3002 (
            .O(N__16545),
            .I(N__16537));
    Span4Mux_v I__3001 (
            .O(N__16542),
            .I(N__16533));
    Span4Mux_h I__3000 (
            .O(N__16537),
            .I(N__16530));
    InMux I__2999 (
            .O(N__16536),
            .I(N__16527));
    Odrv4 I__2998 (
            .O(N__16533),
            .I(frame_decoder_CH1data_0));
    Odrv4 I__2997 (
            .O(N__16530),
            .I(frame_decoder_CH1data_0));
    LocalMux I__2996 (
            .O(N__16527),
            .I(frame_decoder_CH1data_0));
    CascadeMux I__2995 (
            .O(N__16520),
            .I(N__16517));
    InMux I__2994 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__2993 (
            .O(N__16514),
            .I(\scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__2992 (
            .O(N__16511),
            .I(N__16507));
    CascadeMux I__2991 (
            .O(N__16510),
            .I(N__16504));
    LocalMux I__2990 (
            .O(N__16507),
            .I(N__16499));
    InMux I__2989 (
            .O(N__16504),
            .I(N__16494));
    InMux I__2988 (
            .O(N__16503),
            .I(N__16494));
    InMux I__2987 (
            .O(N__16502),
            .I(N__16491));
    Span4Mux_v I__2986 (
            .O(N__16499),
            .I(N__16486));
    LocalMux I__2985 (
            .O(N__16494),
            .I(N__16486));
    LocalMux I__2984 (
            .O(N__16491),
            .I(\scaler_1.un2_source_data_0 ));
    Odrv4 I__2983 (
            .O(N__16486),
            .I(\scaler_1.un2_source_data_0 ));
    InMux I__2982 (
            .O(N__16481),
            .I(\scaler_1.un2_source_data_0_cry_1 ));
    CascadeMux I__2981 (
            .O(N__16478),
            .I(N__16475));
    InMux I__2980 (
            .O(N__16475),
            .I(N__16469));
    InMux I__2979 (
            .O(N__16474),
            .I(N__16469));
    LocalMux I__2978 (
            .O(N__16469),
            .I(N__16466));
    Odrv4 I__2977 (
            .O(N__16466),
            .I(\scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ));
    InMux I__2976 (
            .O(N__16463),
            .I(\scaler_1.un2_source_data_0_cry_2 ));
    CascadeMux I__2975 (
            .O(N__16460),
            .I(N__16456));
    CascadeMux I__2974 (
            .O(N__16459),
            .I(N__16452));
    InMux I__2973 (
            .O(N__16456),
            .I(N__16446));
    InMux I__2972 (
            .O(N__16455),
            .I(N__16446));
    InMux I__2971 (
            .O(N__16452),
            .I(N__16443));
    InMux I__2970 (
            .O(N__16451),
            .I(N__16440));
    LocalMux I__2969 (
            .O(N__16446),
            .I(N__16437));
    LocalMux I__2968 (
            .O(N__16443),
            .I(N__16434));
    LocalMux I__2967 (
            .O(N__16440),
            .I(frame_decoder_OFF3data_0));
    Odrv4 I__2966 (
            .O(N__16437),
            .I(frame_decoder_OFF3data_0));
    Odrv4 I__2965 (
            .O(N__16434),
            .I(frame_decoder_OFF3data_0));
    CascadeMux I__2964 (
            .O(N__16427),
            .I(N__16424));
    InMux I__2963 (
            .O(N__16424),
            .I(N__16421));
    LocalMux I__2962 (
            .O(N__16421),
            .I(N__16418));
    Odrv4 I__2961 (
            .O(N__16418),
            .I(frame_decoder_OFF3data_1));
    InMux I__2960 (
            .O(N__16415),
            .I(\scaler_3.un3_source_data_0_cry_0 ));
    CascadeMux I__2959 (
            .O(N__16412),
            .I(N__16409));
    InMux I__2958 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2957 (
            .O(N__16406),
            .I(N__16403));
    Odrv4 I__2956 (
            .O(N__16403),
            .I(frame_decoder_OFF3data_2));
    InMux I__2955 (
            .O(N__16400),
            .I(\scaler_3.un3_source_data_0_cry_1 ));
    InMux I__2954 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__2953 (
            .O(N__16394),
            .I(N__16391));
    Odrv4 I__2952 (
            .O(N__16391),
            .I(frame_decoder_OFF3data_3));
    InMux I__2951 (
            .O(N__16388),
            .I(\scaler_3.un3_source_data_0_cry_2 ));
    InMux I__2950 (
            .O(N__16385),
            .I(N__16382));
    LocalMux I__2949 (
            .O(N__16382),
            .I(N__16379));
    Odrv4 I__2948 (
            .O(N__16379),
            .I(frame_decoder_OFF3data_4));
    InMux I__2947 (
            .O(N__16376),
            .I(\scaler_3.un3_source_data_0_cry_3 ));
    CascadeMux I__2946 (
            .O(N__16373),
            .I(N__16370));
    InMux I__2945 (
            .O(N__16370),
            .I(N__16367));
    LocalMux I__2944 (
            .O(N__16367),
            .I(N__16364));
    Span4Mux_h I__2943 (
            .O(N__16364),
            .I(N__16361));
    Odrv4 I__2942 (
            .O(N__16361),
            .I(frame_decoder_OFF3data_5));
    InMux I__2941 (
            .O(N__16358),
            .I(\scaler_3.un3_source_data_0_cry_4 ));
    InMux I__2940 (
            .O(N__16355),
            .I(N__16352));
    LocalMux I__2939 (
            .O(N__16352),
            .I(N__16349));
    Odrv4 I__2938 (
            .O(N__16349),
            .I(frame_decoder_OFF3data_6));
    InMux I__2937 (
            .O(N__16346),
            .I(\scaler_3.un3_source_data_0_cry_5 ));
    InMux I__2936 (
            .O(N__16343),
            .I(N__16340));
    LocalMux I__2935 (
            .O(N__16340),
            .I(\scaler_3.un3_source_data_0_axb_7 ));
    InMux I__2934 (
            .O(N__16337),
            .I(\scaler_3.un3_source_data_0_cry_6 ));
    InMux I__2933 (
            .O(N__16334),
            .I(\scaler_2.un2_source_data_0_cry_2 ));
    CascadeMux I__2932 (
            .O(N__16331),
            .I(N__16328));
    InMux I__2931 (
            .O(N__16328),
            .I(N__16322));
    InMux I__2930 (
            .O(N__16327),
            .I(N__16322));
    LocalMux I__2929 (
            .O(N__16322),
            .I(\scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ));
    InMux I__2928 (
            .O(N__16319),
            .I(\scaler_2.un2_source_data_0_cry_3 ));
    CascadeMux I__2927 (
            .O(N__16316),
            .I(N__16313));
    InMux I__2926 (
            .O(N__16313),
            .I(N__16307));
    InMux I__2925 (
            .O(N__16312),
            .I(N__16307));
    LocalMux I__2924 (
            .O(N__16307),
            .I(\scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ));
    InMux I__2923 (
            .O(N__16304),
            .I(\scaler_2.un2_source_data_0_cry_4 ));
    CascadeMux I__2922 (
            .O(N__16301),
            .I(N__16298));
    InMux I__2921 (
            .O(N__16298),
            .I(N__16292));
    InMux I__2920 (
            .O(N__16297),
            .I(N__16292));
    LocalMux I__2919 (
            .O(N__16292),
            .I(\scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ));
    InMux I__2918 (
            .O(N__16289),
            .I(\scaler_2.un2_source_data_0_cry_5 ));
    CascadeMux I__2917 (
            .O(N__16286),
            .I(N__16283));
    InMux I__2916 (
            .O(N__16283),
            .I(N__16277));
    InMux I__2915 (
            .O(N__16282),
            .I(N__16277));
    LocalMux I__2914 (
            .O(N__16277),
            .I(\scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ));
    InMux I__2913 (
            .O(N__16274),
            .I(\scaler_2.un2_source_data_0_cry_6 ));
    CascadeMux I__2912 (
            .O(N__16271),
            .I(N__16268));
    InMux I__2911 (
            .O(N__16268),
            .I(N__16262));
    InMux I__2910 (
            .O(N__16267),
            .I(N__16262));
    LocalMux I__2909 (
            .O(N__16262),
            .I(\scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ));
    InMux I__2908 (
            .O(N__16259),
            .I(\scaler_2.un2_source_data_0_cry_7 ));
    InMux I__2907 (
            .O(N__16256),
            .I(N__16252));
    InMux I__2906 (
            .O(N__16255),
            .I(N__16249));
    LocalMux I__2905 (
            .O(N__16252),
            .I(N__16246));
    LocalMux I__2904 (
            .O(N__16249),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ));
    Odrv4 I__2903 (
            .O(N__16246),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ));
    CascadeMux I__2902 (
            .O(N__16241),
            .I(N__16238));
    InMux I__2901 (
            .O(N__16238),
            .I(N__16235));
    LocalMux I__2900 (
            .O(N__16235),
            .I(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ));
    InMux I__2899 (
            .O(N__16232),
            .I(bfn_10_14_0_));
    InMux I__2898 (
            .O(N__16229),
            .I(\scaler_2.un2_source_data_0_cry_9 ));
    InMux I__2897 (
            .O(N__16226),
            .I(N__16223));
    LocalMux I__2896 (
            .O(N__16223),
            .I(N__16220));
    Span4Mux_h I__2895 (
            .O(N__16220),
            .I(N__16217));
    Span4Mux_v I__2894 (
            .O(N__16217),
            .I(N__16214));
    Odrv4 I__2893 (
            .O(N__16214),
            .I(scaler_4_data_5));
    CascadeMux I__2892 (
            .O(N__16211),
            .I(N__16208));
    InMux I__2891 (
            .O(N__16208),
            .I(N__16205));
    LocalMux I__2890 (
            .O(N__16205),
            .I(\scaler_2.un2_source_data_0_cry_1_c_RNO_0 ));
    InMux I__2889 (
            .O(N__16202),
            .I(N__16197));
    InMux I__2888 (
            .O(N__16201),
            .I(N__16194));
    CascadeMux I__2887 (
            .O(N__16200),
            .I(N__16191));
    LocalMux I__2886 (
            .O(N__16197),
            .I(N__16187));
    LocalMux I__2885 (
            .O(N__16194),
            .I(N__16184));
    InMux I__2884 (
            .O(N__16191),
            .I(N__16179));
    InMux I__2883 (
            .O(N__16190),
            .I(N__16179));
    Odrv4 I__2882 (
            .O(N__16187),
            .I(\scaler_2.un2_source_data_0 ));
    Odrv4 I__2881 (
            .O(N__16184),
            .I(\scaler_2.un2_source_data_0 ));
    LocalMux I__2880 (
            .O(N__16179),
            .I(\scaler_2.un2_source_data_0 ));
    InMux I__2879 (
            .O(N__16172),
            .I(\scaler_2.un2_source_data_0_cry_1 ));
    CascadeMux I__2878 (
            .O(N__16169),
            .I(N__16166));
    InMux I__2877 (
            .O(N__16166),
            .I(N__16160));
    InMux I__2876 (
            .O(N__16165),
            .I(N__16160));
    LocalMux I__2875 (
            .O(N__16160),
            .I(\scaler_2.un3_source_data_0_cry_1_c_RNILSPH ));
    InMux I__2874 (
            .O(N__16157),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__2873 (
            .O(N__16154),
            .I(N__16151));
    LocalMux I__2872 (
            .O(N__16151),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__2871 (
            .O(N__16148),
            .I(N__16143));
    CascadeMux I__2870 (
            .O(N__16147),
            .I(N__16140));
    InMux I__2869 (
            .O(N__16146),
            .I(N__16136));
    LocalMux I__2868 (
            .O(N__16143),
            .I(N__16133));
    InMux I__2867 (
            .O(N__16140),
            .I(N__16128));
    InMux I__2866 (
            .O(N__16139),
            .I(N__16128));
    LocalMux I__2865 (
            .O(N__16136),
            .I(N__16120));
    Span4Mux_h I__2864 (
            .O(N__16133),
            .I(N__16115));
    LocalMux I__2863 (
            .O(N__16128),
            .I(N__16115));
    InMux I__2862 (
            .O(N__16127),
            .I(N__16108));
    InMux I__2861 (
            .O(N__16126),
            .I(N__16108));
    InMux I__2860 (
            .O(N__16125),
            .I(N__16108));
    InMux I__2859 (
            .O(N__16124),
            .I(N__16103));
    InMux I__2858 (
            .O(N__16123),
            .I(N__16103));
    Odrv4 I__2857 (
            .O(N__16120),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    Odrv4 I__2856 (
            .O(N__16115),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__2855 (
            .O(N__16108),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__2854 (
            .O(N__16103),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    InMux I__2853 (
            .O(N__16094),
            .I(N__16091));
    LocalMux I__2852 (
            .O(N__16091),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__2851 (
            .O(N__16088),
            .I(N__16085));
    LocalMux I__2850 (
            .O(N__16085),
            .I(N__16082));
    Span4Mux_v I__2849 (
            .O(N__16082),
            .I(N__16079));
    Odrv4 I__2848 (
            .O(N__16079),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ));
    CascadeMux I__2847 (
            .O(N__16076),
            .I(N__16073));
    InMux I__2846 (
            .O(N__16073),
            .I(N__16068));
    InMux I__2845 (
            .O(N__16072),
            .I(N__16065));
    InMux I__2844 (
            .O(N__16071),
            .I(N__16062));
    LocalMux I__2843 (
            .O(N__16068),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__2842 (
            .O(N__16065),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__2841 (
            .O(N__16062),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    InMux I__2840 (
            .O(N__16055),
            .I(N__16052));
    LocalMux I__2839 (
            .O(N__16052),
            .I(N__16047));
    InMux I__2838 (
            .O(N__16051),
            .I(N__16042));
    InMux I__2837 (
            .O(N__16050),
            .I(N__16042));
    Odrv4 I__2836 (
            .O(N__16047),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__2835 (
            .O(N__16042),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    CascadeMux I__2834 (
            .O(N__16037),
            .I(N__16034));
    InMux I__2833 (
            .O(N__16034),
            .I(N__16030));
    InMux I__2832 (
            .O(N__16033),
            .I(N__16027));
    LocalMux I__2831 (
            .O(N__16030),
            .I(N__16024));
    LocalMux I__2830 (
            .O(N__16027),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    Odrv4 I__2829 (
            .O(N__16024),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    CascadeMux I__2828 (
            .O(N__16019),
            .I(N__16013));
    CascadeMux I__2827 (
            .O(N__16018),
            .I(N__16010));
    InMux I__2826 (
            .O(N__16017),
            .I(N__16001));
    InMux I__2825 (
            .O(N__16016),
            .I(N__16001));
    InMux I__2824 (
            .O(N__16013),
            .I(N__16001));
    InMux I__2823 (
            .O(N__16010),
            .I(N__16001));
    LocalMux I__2822 (
            .O(N__16001),
            .I(N__15998));
    Span12Mux_s8_v I__2821 (
            .O(N__15998),
            .I(N__15994));
    InMux I__2820 (
            .O(N__15997),
            .I(N__15991));
    Odrv12 I__2819 (
            .O(N__15994),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_162_d ));
    LocalMux I__2818 (
            .O(N__15991),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_162_d ));
    CascadeMux I__2817 (
            .O(N__15986),
            .I(N__15982));
    InMux I__2816 (
            .O(N__15985),
            .I(N__15979));
    InMux I__2815 (
            .O(N__15982),
            .I(N__15975));
    LocalMux I__2814 (
            .O(N__15979),
            .I(N__15972));
    CascadeMux I__2813 (
            .O(N__15978),
            .I(N__15969));
    LocalMux I__2812 (
            .O(N__15975),
            .I(N__15964));
    Span4Mux_h I__2811 (
            .O(N__15972),
            .I(N__15964));
    InMux I__2810 (
            .O(N__15969),
            .I(N__15961));
    Odrv4 I__2809 (
            .O(N__15964),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__2808 (
            .O(N__15961),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__2807 (
            .O(N__15956),
            .I(N__15951));
    InMux I__2806 (
            .O(N__15955),
            .I(N__15946));
    InMux I__2805 (
            .O(N__15954),
            .I(N__15946));
    LocalMux I__2804 (
            .O(N__15951),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__2803 (
            .O(N__15946),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__2802 (
            .O(N__15941),
            .I(N__15938));
    LocalMux I__2801 (
            .O(N__15938),
            .I(N__15935));
    Odrv4 I__2800 (
            .O(N__15935),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__2799 (
            .O(N__15932),
            .I(N__15929));
    LocalMux I__2798 (
            .O(N__15929),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__2797 (
            .O(N__15926),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__2796 (
            .O(N__15923),
            .I(N__15920));
    LocalMux I__2795 (
            .O(N__15920),
            .I(N__15916));
    InMux I__2794 (
            .O(N__15919),
            .I(N__15913));
    Span4Mux_v I__2793 (
            .O(N__15916),
            .I(N__15910));
    LocalMux I__2792 (
            .O(N__15913),
            .I(N__15907));
    Odrv4 I__2791 (
            .O(N__15910),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    Odrv4 I__2790 (
            .O(N__15907),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    CascadeMux I__2789 (
            .O(N__15902),
            .I(N__15899));
    InMux I__2788 (
            .O(N__15899),
            .I(N__15896));
    LocalMux I__2787 (
            .O(N__15896),
            .I(N__15893));
    Odrv12 I__2786 (
            .O(N__15893),
            .I(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ));
    InMux I__2785 (
            .O(N__15890),
            .I(N__15887));
    LocalMux I__2784 (
            .O(N__15887),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__2783 (
            .O(N__15884),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__2782 (
            .O(N__15881),
            .I(N__15878));
    LocalMux I__2781 (
            .O(N__15878),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__2780 (
            .O(N__15875),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__2779 (
            .O(N__15872),
            .I(N__15869));
    LocalMux I__2778 (
            .O(N__15869),
            .I(N__15866));
    Span4Mux_h I__2777 (
            .O(N__15866),
            .I(N__15863));
    Odrv4 I__2776 (
            .O(N__15863),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__2775 (
            .O(N__15860),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__2774 (
            .O(N__15857),
            .I(N__15854));
    LocalMux I__2773 (
            .O(N__15854),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__2772 (
            .O(N__15851),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__2771 (
            .O(N__15848),
            .I(N__15845));
    LocalMux I__2770 (
            .O(N__15845),
            .I(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ));
    CascadeMux I__2769 (
            .O(N__15842),
            .I(N__15839));
    InMux I__2768 (
            .O(N__15839),
            .I(N__15836));
    LocalMux I__2767 (
            .O(N__15836),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ));
    InMux I__2766 (
            .O(N__15833),
            .I(N__15830));
    LocalMux I__2765 (
            .O(N__15830),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__2764 (
            .O(N__15827),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__2763 (
            .O(N__15824),
            .I(N__15821));
    LocalMux I__2762 (
            .O(N__15821),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__2761 (
            .O(N__15818),
            .I(bfn_9_26_0_));
    InMux I__2760 (
            .O(N__15815),
            .I(N__15812));
    LocalMux I__2759 (
            .O(N__15812),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    CascadeMux I__2758 (
            .O(N__15809),
            .I(N__15806));
    InMux I__2757 (
            .O(N__15806),
            .I(N__15803));
    LocalMux I__2756 (
            .O(N__15803),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__2755 (
            .O(N__15800),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__2754 (
            .O(N__15797),
            .I(N__15794));
    LocalMux I__2753 (
            .O(N__15794),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    CascadeMux I__2752 (
            .O(N__15791),
            .I(N__15788));
    InMux I__2751 (
            .O(N__15788),
            .I(N__15785));
    LocalMux I__2750 (
            .O(N__15785),
            .I(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ));
    CascadeMux I__2749 (
            .O(N__15782),
            .I(N__15779));
    InMux I__2748 (
            .O(N__15779),
            .I(N__15776));
    LocalMux I__2747 (
            .O(N__15776),
            .I(N__15773));
    Odrv4 I__2746 (
            .O(N__15773),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__2745 (
            .O(N__15770),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__2744 (
            .O(N__15767),
            .I(N__15764));
    LocalMux I__2743 (
            .O(N__15764),
            .I(N__15760));
    InMux I__2742 (
            .O(N__15763),
            .I(N__15757));
    Odrv4 I__2741 (
            .O(N__15760),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    LocalMux I__2740 (
            .O(N__15757),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    CascadeMux I__2739 (
            .O(N__15752),
            .I(N__15749));
    InMux I__2738 (
            .O(N__15749),
            .I(N__15746));
    LocalMux I__2737 (
            .O(N__15746),
            .I(N__15743));
    Odrv4 I__2736 (
            .O(N__15743),
            .I(\ppm_encoder_1.init_pulses_RNI60223Z0Z_3 ));
    InMux I__2735 (
            .O(N__15740),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__2734 (
            .O(N__15737),
            .I(N__15733));
    InMux I__2733 (
            .O(N__15736),
            .I(N__15730));
    LocalMux I__2732 (
            .O(N__15733),
            .I(N__15727));
    LocalMux I__2731 (
            .O(N__15730),
            .I(N__15724));
    Span4Mux_v I__2730 (
            .O(N__15727),
            .I(N__15721));
    Span4Mux_h I__2729 (
            .O(N__15724),
            .I(N__15718));
    Odrv4 I__2728 (
            .O(N__15721),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    Odrv4 I__2727 (
            .O(N__15718),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    CascadeMux I__2726 (
            .O(N__15713),
            .I(N__15710));
    InMux I__2725 (
            .O(N__15710),
            .I(N__15707));
    LocalMux I__2724 (
            .O(N__15707),
            .I(N__15704));
    Odrv4 I__2723 (
            .O(N__15704),
            .I(\ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4 ));
    InMux I__2722 (
            .O(N__15701),
            .I(N__15698));
    LocalMux I__2721 (
            .O(N__15698),
            .I(N__15695));
    Span4Mux_h I__2720 (
            .O(N__15695),
            .I(N__15692));
    Odrv4 I__2719 (
            .O(N__15692),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__2718 (
            .O(N__15689),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    CascadeMux I__2717 (
            .O(N__15686),
            .I(N__15683));
    InMux I__2716 (
            .O(N__15683),
            .I(N__15680));
    LocalMux I__2715 (
            .O(N__15680),
            .I(\ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5 ));
    InMux I__2714 (
            .O(N__15677),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__2713 (
            .O(N__15674),
            .I(N__15671));
    LocalMux I__2712 (
            .O(N__15671),
            .I(N__15668));
    Span4Mux_h I__2711 (
            .O(N__15668),
            .I(N__15665));
    Odrv4 I__2710 (
            .O(N__15665),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__2709 (
            .O(N__15662),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__2708 (
            .O(N__15659),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    CascadeMux I__2707 (
            .O(N__15656),
            .I(N__15653));
    InMux I__2706 (
            .O(N__15653),
            .I(N__15650));
    LocalMux I__2705 (
            .O(N__15650),
            .I(N__15647));
    Odrv12 I__2704 (
            .O(N__15647),
            .I(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ));
    InMux I__2703 (
            .O(N__15644),
            .I(bfn_9_25_0_));
    CascadeMux I__2702 (
            .O(N__15641),
            .I(N__15638));
    InMux I__2701 (
            .O(N__15638),
            .I(N__15635));
    LocalMux I__2700 (
            .O(N__15635),
            .I(N__15632));
    Odrv12 I__2699 (
            .O(N__15632),
            .I(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ));
    InMux I__2698 (
            .O(N__15629),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__2697 (
            .O(N__15626),
            .I(N__15621));
    CascadeMux I__2696 (
            .O(N__15625),
            .I(N__15618));
    InMux I__2695 (
            .O(N__15624),
            .I(N__15612));
    LocalMux I__2694 (
            .O(N__15621),
            .I(N__15609));
    InMux I__2693 (
            .O(N__15618),
            .I(N__15604));
    InMux I__2692 (
            .O(N__15617),
            .I(N__15604));
    InMux I__2691 (
            .O(N__15616),
            .I(N__15599));
    InMux I__2690 (
            .O(N__15615),
            .I(N__15599));
    LocalMux I__2689 (
            .O(N__15612),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv12 I__2688 (
            .O(N__15609),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__2687 (
            .O(N__15604),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__2686 (
            .O(N__15599),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__2685 (
            .O(N__15590),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ));
    InMux I__2684 (
            .O(N__15587),
            .I(N__15584));
    LocalMux I__2683 (
            .O(N__15584),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5 ));
    InMux I__2682 (
            .O(N__15581),
            .I(N__15575));
    InMux I__2681 (
            .O(N__15580),
            .I(N__15575));
    LocalMux I__2680 (
            .O(N__15575),
            .I(N__15572));
    Odrv4 I__2679 (
            .O(N__15572),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    InMux I__2678 (
            .O(N__15569),
            .I(N__15563));
    InMux I__2677 (
            .O(N__15568),
            .I(N__15563));
    LocalMux I__2676 (
            .O(N__15563),
            .I(N__15560));
    Odrv4 I__2675 (
            .O(N__15560),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__2674 (
            .O(N__15557),
            .I(\ppm_encoder_1.N_300_cascade_ ));
    InMux I__2673 (
            .O(N__15554),
            .I(N__15551));
    LocalMux I__2672 (
            .O(N__15551),
            .I(N__15548));
    Odrv12 I__2671 (
            .O(N__15548),
            .I(scaler_2_data_5));
    CascadeMux I__2670 (
            .O(N__15545),
            .I(N__15541));
    InMux I__2669 (
            .O(N__15544),
            .I(N__15538));
    InMux I__2668 (
            .O(N__15541),
            .I(N__15535));
    LocalMux I__2667 (
            .O(N__15538),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    LocalMux I__2666 (
            .O(N__15535),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__2665 (
            .O(N__15530),
            .I(N__15526));
    InMux I__2664 (
            .O(N__15529),
            .I(N__15523));
    LocalMux I__2663 (
            .O(N__15526),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    LocalMux I__2662 (
            .O(N__15523),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    InMux I__2661 (
            .O(N__15518),
            .I(N__15515));
    LocalMux I__2660 (
            .O(N__15515),
            .I(N__15511));
    InMux I__2659 (
            .O(N__15514),
            .I(N__15508));
    Odrv12 I__2658 (
            .O(N__15511),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    LocalMux I__2657 (
            .O(N__15508),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    CascadeMux I__2656 (
            .O(N__15503),
            .I(N__15500));
    InMux I__2655 (
            .O(N__15500),
            .I(N__15497));
    LocalMux I__2654 (
            .O(N__15497),
            .I(N__15494));
    Odrv4 I__2653 (
            .O(N__15494),
            .I(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ));
    InMux I__2652 (
            .O(N__15491),
            .I(N__15488));
    LocalMux I__2651 (
            .O(N__15488),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__2650 (
            .O(N__15485),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__2649 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__2648 (
            .O(N__15479),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9 ));
    InMux I__2647 (
            .O(N__15476),
            .I(N__15471));
    InMux I__2646 (
            .O(N__15475),
            .I(N__15468));
    InMux I__2645 (
            .O(N__15474),
            .I(N__15465));
    LocalMux I__2644 (
            .O(N__15471),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__2643 (
            .O(N__15468),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__2642 (
            .O(N__15465),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__2641 (
            .O(N__15458),
            .I(N__15453));
    InMux I__2640 (
            .O(N__15457),
            .I(N__15450));
    InMux I__2639 (
            .O(N__15456),
            .I(N__15447));
    InMux I__2638 (
            .O(N__15453),
            .I(N__15444));
    LocalMux I__2637 (
            .O(N__15450),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__2636 (
            .O(N__15447),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__2635 (
            .O(N__15444),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    InMux I__2634 (
            .O(N__15437),
            .I(N__15433));
    InMux I__2633 (
            .O(N__15436),
            .I(N__15430));
    LocalMux I__2632 (
            .O(N__15433),
            .I(N__15425));
    LocalMux I__2631 (
            .O(N__15430),
            .I(N__15425));
    Odrv4 I__2630 (
            .O(N__15425),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__2629 (
            .O(N__15422),
            .I(N__15418));
    InMux I__2628 (
            .O(N__15421),
            .I(N__15415));
    LocalMux I__2627 (
            .O(N__15418),
            .I(N__15412));
    LocalMux I__2626 (
            .O(N__15415),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    Odrv4 I__2625 (
            .O(N__15412),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    CascadeMux I__2624 (
            .O(N__15407),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ));
    InMux I__2623 (
            .O(N__15404),
            .I(N__15400));
    InMux I__2622 (
            .O(N__15403),
            .I(N__15397));
    LocalMux I__2621 (
            .O(N__15400),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    LocalMux I__2620 (
            .O(N__15397),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    InMux I__2619 (
            .O(N__15392),
            .I(N__15388));
    InMux I__2618 (
            .O(N__15391),
            .I(N__15385));
    LocalMux I__2617 (
            .O(N__15388),
            .I(N__15380));
    LocalMux I__2616 (
            .O(N__15385),
            .I(N__15380));
    Span4Mux_v I__2615 (
            .O(N__15380),
            .I(N__15377));
    Odrv4 I__2614 (
            .O(N__15377),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    CascadeMux I__2613 (
            .O(N__15374),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    CascadeMux I__2612 (
            .O(N__15371),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ));
    InMux I__2611 (
            .O(N__15368),
            .I(N__15365));
    LocalMux I__2610 (
            .O(N__15365),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4 ));
    InMux I__2609 (
            .O(N__15362),
            .I(N__15359));
    LocalMux I__2608 (
            .O(N__15359),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    CascadeMux I__2607 (
            .O(N__15356),
            .I(\ppm_encoder_1.N_306_cascade_ ));
    InMux I__2606 (
            .O(N__15353),
            .I(N__15344));
    InMux I__2605 (
            .O(N__15352),
            .I(N__15344));
    InMux I__2604 (
            .O(N__15351),
            .I(N__15344));
    LocalMux I__2603 (
            .O(N__15344),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    CascadeMux I__2602 (
            .O(N__15341),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ));
    InMux I__2601 (
            .O(N__15338),
            .I(N__15335));
    LocalMux I__2600 (
            .O(N__15335),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8 ));
    CascadeMux I__2599 (
            .O(N__15332),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ));
    InMux I__2598 (
            .O(N__15329),
            .I(N__15322));
    InMux I__2597 (
            .O(N__15328),
            .I(N__15322));
    InMux I__2596 (
            .O(N__15327),
            .I(N__15319));
    LocalMux I__2595 (
            .O(N__15322),
            .I(N__15310));
    LocalMux I__2594 (
            .O(N__15319),
            .I(N__15310));
    InMux I__2593 (
            .O(N__15318),
            .I(N__15306));
    InMux I__2592 (
            .O(N__15317),
            .I(N__15301));
    InMux I__2591 (
            .O(N__15316),
            .I(N__15301));
    InMux I__2590 (
            .O(N__15315),
            .I(N__15298));
    Span4Mux_v I__2589 (
            .O(N__15310),
            .I(N__15295));
    InMux I__2588 (
            .O(N__15309),
            .I(N__15292));
    LocalMux I__2587 (
            .O(N__15306),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__2586 (
            .O(N__15301),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__2585 (
            .O(N__15298),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    Odrv4 I__2584 (
            .O(N__15295),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__2583 (
            .O(N__15292),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    InMux I__2582 (
            .O(N__15281),
            .I(N__15275));
    InMux I__2581 (
            .O(N__15280),
            .I(N__15275));
    LocalMux I__2580 (
            .O(N__15275),
            .I(\uart_frame_decoder.count8_THRU_CO ));
    CascadeMux I__2579 (
            .O(N__15272),
            .I(N__15263));
    CascadeMux I__2578 (
            .O(N__15271),
            .I(N__15260));
    CascadeMux I__2577 (
            .O(N__15270),
            .I(N__15257));
    CascadeMux I__2576 (
            .O(N__15269),
            .I(N__15254));
    InMux I__2575 (
            .O(N__15268),
            .I(N__15248));
    InMux I__2574 (
            .O(N__15267),
            .I(N__15243));
    InMux I__2573 (
            .O(N__15266),
            .I(N__15240));
    InMux I__2572 (
            .O(N__15263),
            .I(N__15225));
    InMux I__2571 (
            .O(N__15260),
            .I(N__15225));
    InMux I__2570 (
            .O(N__15257),
            .I(N__15225));
    InMux I__2569 (
            .O(N__15254),
            .I(N__15225));
    InMux I__2568 (
            .O(N__15253),
            .I(N__15225));
    InMux I__2567 (
            .O(N__15252),
            .I(N__15225));
    InMux I__2566 (
            .O(N__15251),
            .I(N__15225));
    LocalMux I__2565 (
            .O(N__15248),
            .I(N__15222));
    InMux I__2564 (
            .O(N__15247),
            .I(N__15218));
    InMux I__2563 (
            .O(N__15246),
            .I(N__15215));
    LocalMux I__2562 (
            .O(N__15243),
            .I(N__15212));
    LocalMux I__2561 (
            .O(N__15240),
            .I(N__15209));
    LocalMux I__2560 (
            .O(N__15225),
            .I(N__15206));
    Span4Mux_v I__2559 (
            .O(N__15222),
            .I(N__15203));
    InMux I__2558 (
            .O(N__15221),
            .I(N__15200));
    LocalMux I__2557 (
            .O(N__15218),
            .I(N__15193));
    LocalMux I__2556 (
            .O(N__15215),
            .I(N__15193));
    Sp12to4 I__2555 (
            .O(N__15212),
            .I(N__15193));
    Span4Mux_h I__2554 (
            .O(N__15209),
            .I(N__15190));
    Span4Mux_v I__2553 (
            .O(N__15206),
            .I(N__15187));
    Span4Mux_v I__2552 (
            .O(N__15203),
            .I(N__15184));
    LocalMux I__2551 (
            .O(N__15200),
            .I(N__15181));
    Span12Mux_v I__2550 (
            .O(N__15193),
            .I(N__15178));
    Odrv4 I__2549 (
            .O(N__15190),
            .I(uart_input_pc_sync));
    Odrv4 I__2548 (
            .O(N__15187),
            .I(uart_input_pc_sync));
    Odrv4 I__2547 (
            .O(N__15184),
            .I(uart_input_pc_sync));
    Odrv4 I__2546 (
            .O(N__15181),
            .I(uart_input_pc_sync));
    Odrv12 I__2545 (
            .O(N__15178),
            .I(uart_input_pc_sync));
    InMux I__2544 (
            .O(N__15167),
            .I(N__15160));
    InMux I__2543 (
            .O(N__15166),
            .I(N__15160));
    InMux I__2542 (
            .O(N__15165),
            .I(N__15157));
    LocalMux I__2541 (
            .O(N__15160),
            .I(N__15154));
    LocalMux I__2540 (
            .O(N__15157),
            .I(N__15151));
    Span4Mux_h I__2539 (
            .O(N__15154),
            .I(N__15148));
    Span4Mux_h I__2538 (
            .O(N__15151),
            .I(N__15145));
    Span4Mux_v I__2537 (
            .O(N__15148),
            .I(N__15142));
    Odrv4 I__2536 (
            .O(N__15145),
            .I(\uart_pc.state_1_sqmuxa ));
    Odrv4 I__2535 (
            .O(N__15142),
            .I(\uart_pc.state_1_sqmuxa ));
    CascadeMux I__2534 (
            .O(N__15137),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ));
    InMux I__2533 (
            .O(N__15134),
            .I(N__15131));
    LocalMux I__2532 (
            .O(N__15131),
            .I(\scaler_2.N_520_i_l_ofxZ0 ));
    InMux I__2531 (
            .O(N__15128),
            .I(N__15125));
    LocalMux I__2530 (
            .O(N__15125),
            .I(N__15122));
    Span4Mux_v I__2529 (
            .O(N__15122),
            .I(N__15119));
    Odrv4 I__2528 (
            .O(N__15119),
            .I(scaler_1_data_5));
    InMux I__2527 (
            .O(N__15116),
            .I(N__15113));
    LocalMux I__2526 (
            .O(N__15113),
            .I(N__15110));
    Span4Mux_v I__2525 (
            .O(N__15110),
            .I(N__15107));
    Odrv4 I__2524 (
            .O(N__15107),
            .I(scaler_3_data_5));
    InMux I__2523 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__2522 (
            .O(N__15101),
            .I(N__15098));
    Span4Mux_v I__2521 (
            .O(N__15098),
            .I(N__15094));
    InMux I__2520 (
            .O(N__15097),
            .I(N__15091));
    Odrv4 I__2519 (
            .O(N__15094),
            .I(scaler_1_data_4));
    LocalMux I__2518 (
            .O(N__15091),
            .I(scaler_1_data_4));
    InMux I__2517 (
            .O(N__15086),
            .I(N__15082));
    CascadeMux I__2516 (
            .O(N__15085),
            .I(N__15077));
    LocalMux I__2515 (
            .O(N__15082),
            .I(N__15074));
    InMux I__2514 (
            .O(N__15081),
            .I(N__15071));
    InMux I__2513 (
            .O(N__15080),
            .I(N__15068));
    InMux I__2512 (
            .O(N__15077),
            .I(N__15065));
    Span4Mux_v I__2511 (
            .O(N__15074),
            .I(N__15060));
    LocalMux I__2510 (
            .O(N__15071),
            .I(N__15060));
    LocalMux I__2509 (
            .O(N__15068),
            .I(N__15057));
    LocalMux I__2508 (
            .O(N__15065),
            .I(N__15054));
    Odrv4 I__2507 (
            .O(N__15060),
            .I(frame_decoder_OFF2data_0));
    Odrv4 I__2506 (
            .O(N__15057),
            .I(frame_decoder_OFF2data_0));
    Odrv4 I__2505 (
            .O(N__15054),
            .I(frame_decoder_OFF2data_0));
    InMux I__2504 (
            .O(N__15047),
            .I(N__15043));
    InMux I__2503 (
            .O(N__15046),
            .I(N__15040));
    LocalMux I__2502 (
            .O(N__15043),
            .I(N__15033));
    LocalMux I__2501 (
            .O(N__15040),
            .I(N__15033));
    InMux I__2500 (
            .O(N__15039),
            .I(N__15030));
    InMux I__2499 (
            .O(N__15038),
            .I(N__15027));
    Odrv12 I__2498 (
            .O(N__15033),
            .I(frame_decoder_CH2data_0));
    LocalMux I__2497 (
            .O(N__15030),
            .I(frame_decoder_CH2data_0));
    LocalMux I__2496 (
            .O(N__15027),
            .I(frame_decoder_CH2data_0));
    InMux I__2495 (
            .O(N__15020),
            .I(N__15017));
    LocalMux I__2494 (
            .O(N__15017),
            .I(N__15013));
    CascadeMux I__2493 (
            .O(N__15016),
            .I(N__15010));
    Span4Mux_h I__2492 (
            .O(N__15013),
            .I(N__15007));
    InMux I__2491 (
            .O(N__15010),
            .I(N__15004));
    Odrv4 I__2490 (
            .O(N__15007),
            .I(scaler_2_data_4));
    LocalMux I__2489 (
            .O(N__15004),
            .I(scaler_2_data_4));
    InMux I__2488 (
            .O(N__14999),
            .I(N__14995));
    InMux I__2487 (
            .O(N__14998),
            .I(N__14992));
    LocalMux I__2486 (
            .O(N__14995),
            .I(N__14989));
    LocalMux I__2485 (
            .O(N__14992),
            .I(N__14986));
    Odrv4 I__2484 (
            .O(N__14989),
            .I(scaler_3_data_4));
    Odrv4 I__2483 (
            .O(N__14986),
            .I(scaler_3_data_4));
    InMux I__2482 (
            .O(N__14981),
            .I(N__14978));
    LocalMux I__2481 (
            .O(N__14978),
            .I(N__14974));
    CascadeMux I__2480 (
            .O(N__14977),
            .I(N__14971));
    Span4Mux_v I__2479 (
            .O(N__14974),
            .I(N__14968));
    InMux I__2478 (
            .O(N__14971),
            .I(N__14965));
    Odrv4 I__2477 (
            .O(N__14968),
            .I(scaler_4_data_4));
    LocalMux I__2476 (
            .O(N__14965),
            .I(scaler_4_data_4));
    InMux I__2475 (
            .O(N__14960),
            .I(N__14957));
    LocalMux I__2474 (
            .O(N__14957),
            .I(frame_decoder_CH2data_4));
    CascadeMux I__2473 (
            .O(N__14954),
            .I(N__14951));
    InMux I__2472 (
            .O(N__14951),
            .I(N__14948));
    LocalMux I__2471 (
            .O(N__14948),
            .I(frame_decoder_OFF2data_4));
    InMux I__2470 (
            .O(N__14945),
            .I(\scaler_2.un3_source_data_0_cry_3 ));
    InMux I__2469 (
            .O(N__14942),
            .I(N__14939));
    LocalMux I__2468 (
            .O(N__14939),
            .I(frame_decoder_CH2data_5));
    CascadeMux I__2467 (
            .O(N__14936),
            .I(N__14933));
    InMux I__2466 (
            .O(N__14933),
            .I(N__14930));
    LocalMux I__2465 (
            .O(N__14930),
            .I(frame_decoder_OFF2data_5));
    InMux I__2464 (
            .O(N__14927),
            .I(\scaler_2.un3_source_data_0_cry_4 ));
    InMux I__2463 (
            .O(N__14924),
            .I(N__14921));
    LocalMux I__2462 (
            .O(N__14921),
            .I(frame_decoder_CH2data_6));
    CascadeMux I__2461 (
            .O(N__14918),
            .I(N__14915));
    InMux I__2460 (
            .O(N__14915),
            .I(N__14912));
    LocalMux I__2459 (
            .O(N__14912),
            .I(frame_decoder_OFF2data_6));
    InMux I__2458 (
            .O(N__14909),
            .I(\scaler_2.un3_source_data_0_cry_5 ));
    InMux I__2457 (
            .O(N__14906),
            .I(\scaler_2.un3_source_data_0_cry_6 ));
    InMux I__2456 (
            .O(N__14903),
            .I(bfn_9_15_0_));
    InMux I__2455 (
            .O(N__14900),
            .I(\scaler_2.un3_source_data_0_cry_8 ));
    InMux I__2454 (
            .O(N__14897),
            .I(N__14894));
    LocalMux I__2453 (
            .O(N__14894),
            .I(N__14890));
    InMux I__2452 (
            .O(N__14893),
            .I(N__14887));
    Span4Mux_v I__2451 (
            .O(N__14890),
            .I(N__14884));
    LocalMux I__2450 (
            .O(N__14887),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    Odrv4 I__2449 (
            .O(N__14884),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    InMux I__2448 (
            .O(N__14879),
            .I(N__14876));
    LocalMux I__2447 (
            .O(N__14876),
            .I(N__14873));
    Sp12to4 I__2446 (
            .O(N__14873),
            .I(N__14870));
    Odrv12 I__2445 (
            .O(N__14870),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__2444 (
            .O(N__14867),
            .I(\uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ));
    InMux I__2443 (
            .O(N__14864),
            .I(N__14861));
    LocalMux I__2442 (
            .O(N__14861),
            .I(frame_decoder_CH2data_1));
    CascadeMux I__2441 (
            .O(N__14858),
            .I(N__14855));
    InMux I__2440 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__2439 (
            .O(N__14852),
            .I(frame_decoder_OFF2data_1));
    InMux I__2438 (
            .O(N__14849),
            .I(\scaler_2.un3_source_data_0_cry_0 ));
    InMux I__2437 (
            .O(N__14846),
            .I(N__14843));
    LocalMux I__2436 (
            .O(N__14843),
            .I(frame_decoder_CH2data_2));
    CascadeMux I__2435 (
            .O(N__14840),
            .I(N__14837));
    InMux I__2434 (
            .O(N__14837),
            .I(N__14834));
    LocalMux I__2433 (
            .O(N__14834),
            .I(frame_decoder_OFF2data_2));
    InMux I__2432 (
            .O(N__14831),
            .I(\scaler_2.un3_source_data_0_cry_1 ));
    InMux I__2431 (
            .O(N__14828),
            .I(N__14825));
    LocalMux I__2430 (
            .O(N__14825),
            .I(frame_decoder_CH2data_3));
    CascadeMux I__2429 (
            .O(N__14822),
            .I(N__14819));
    InMux I__2428 (
            .O(N__14819),
            .I(N__14816));
    LocalMux I__2427 (
            .O(N__14816),
            .I(frame_decoder_OFF2data_3));
    InMux I__2426 (
            .O(N__14813),
            .I(\scaler_2.un3_source_data_0_cry_2 ));
    SRMux I__2425 (
            .O(N__14810),
            .I(N__14805));
    SRMux I__2424 (
            .O(N__14809),
            .I(N__14802));
    SRMux I__2423 (
            .O(N__14808),
            .I(N__14799));
    LocalMux I__2422 (
            .O(N__14805),
            .I(N__14796));
    LocalMux I__2421 (
            .O(N__14802),
            .I(N__14791));
    LocalMux I__2420 (
            .O(N__14799),
            .I(N__14791));
    Odrv4 I__2419 (
            .O(N__14796),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__2418 (
            .O(N__14791),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    InMux I__2417 (
            .O(N__14786),
            .I(N__14783));
    LocalMux I__2416 (
            .O(N__14783),
            .I(\uart_frame_decoder.state_1_ns_i_i_0_0 ));
    CascadeMux I__2415 (
            .O(N__14780),
            .I(N__14777));
    InMux I__2414 (
            .O(N__14777),
            .I(N__14774));
    LocalMux I__2413 (
            .O(N__14774),
            .I(\uart_frame_decoder.N_39_i_1 ));
    CascadeMux I__2412 (
            .O(N__14771),
            .I(N__14766));
    InMux I__2411 (
            .O(N__14770),
            .I(N__14763));
    InMux I__2410 (
            .O(N__14769),
            .I(N__14758));
    InMux I__2409 (
            .O(N__14766),
            .I(N__14758));
    LocalMux I__2408 (
            .O(N__14763),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    LocalMux I__2407 (
            .O(N__14758),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    InMux I__2406 (
            .O(N__14753),
            .I(N__14749));
    InMux I__2405 (
            .O(N__14752),
            .I(N__14746));
    LocalMux I__2404 (
            .O(N__14749),
            .I(\uart_frame_decoder.state_1Z0Z_9 ));
    LocalMux I__2403 (
            .O(N__14746),
            .I(\uart_frame_decoder.state_1Z0Z_9 ));
    CascadeMux I__2402 (
            .O(N__14741),
            .I(N__14738));
    InMux I__2401 (
            .O(N__14738),
            .I(N__14735));
    LocalMux I__2400 (
            .O(N__14735),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa ));
    CascadeMux I__2399 (
            .O(N__14732),
            .I(\uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ));
    InMux I__2398 (
            .O(N__14729),
            .I(N__14726));
    LocalMux I__2397 (
            .O(N__14726),
            .I(N__14722));
    InMux I__2396 (
            .O(N__14725),
            .I(N__14718));
    Span4Mux_v I__2395 (
            .O(N__14722),
            .I(N__14715));
    InMux I__2394 (
            .O(N__14721),
            .I(N__14712));
    LocalMux I__2393 (
            .O(N__14718),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    Odrv4 I__2392 (
            .O(N__14715),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    LocalMux I__2391 (
            .O(N__14712),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    InMux I__2390 (
            .O(N__14705),
            .I(N__14701));
    CascadeMux I__2389 (
            .O(N__14704),
            .I(N__14698));
    LocalMux I__2388 (
            .O(N__14701),
            .I(N__14694));
    InMux I__2387 (
            .O(N__14698),
            .I(N__14688));
    InMux I__2386 (
            .O(N__14697),
            .I(N__14688));
    Span4Mux_v I__2385 (
            .O(N__14694),
            .I(N__14685));
    InMux I__2384 (
            .O(N__14693),
            .I(N__14682));
    LocalMux I__2383 (
            .O(N__14688),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    Odrv4 I__2382 (
            .O(N__14685),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    LocalMux I__2381 (
            .O(N__14682),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    CascadeMux I__2380 (
            .O(N__14675),
            .I(\uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_ ));
    InMux I__2379 (
            .O(N__14672),
            .I(N__14666));
    InMux I__2378 (
            .O(N__14671),
            .I(N__14666));
    LocalMux I__2377 (
            .O(N__14666),
            .I(\uart_frame_decoder.state_1_ns_0_i_o2_0_10 ));
    CascadeMux I__2376 (
            .O(N__14663),
            .I(N__14660));
    InMux I__2375 (
            .O(N__14660),
            .I(N__14657));
    LocalMux I__2374 (
            .O(N__14657),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    CascadeMux I__2373 (
            .O(N__14654),
            .I(N__14651));
    InMux I__2372 (
            .O(N__14651),
            .I(N__14648));
    LocalMux I__2371 (
            .O(N__14648),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__2370 (
            .O(N__14645),
            .I(N__14642));
    LocalMux I__2369 (
            .O(N__14642),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__2368 (
            .O(N__14639),
            .I(N__14636));
    LocalMux I__2367 (
            .O(N__14636),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__2366 (
            .O(N__14633),
            .I(N__14630));
    LocalMux I__2365 (
            .O(N__14630),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__2364 (
            .O(N__14627),
            .I(N__14624));
    LocalMux I__2363 (
            .O(N__14624),
            .I(N__14620));
    CascadeMux I__2362 (
            .O(N__14623),
            .I(N__14617));
    Span4Mux_h I__2361 (
            .O(N__14620),
            .I(N__14614));
    InMux I__2360 (
            .O(N__14617),
            .I(N__14611));
    Odrv4 I__2359 (
            .O(N__14614),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__2358 (
            .O(N__14611),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    CEMux I__2357 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__2356 (
            .O(N__14603),
            .I(N__14598));
    CEMux I__2355 (
            .O(N__14602),
            .I(N__14595));
    CEMux I__2354 (
            .O(N__14601),
            .I(N__14592));
    Span4Mux_h I__2353 (
            .O(N__14598),
            .I(N__14589));
    LocalMux I__2352 (
            .O(N__14595),
            .I(N__14586));
    LocalMux I__2351 (
            .O(N__14592),
            .I(N__14583));
    Odrv4 I__2350 (
            .O(N__14589),
            .I(\uart_pc.state_1_sqmuxa_0 ));
    Odrv4 I__2349 (
            .O(N__14586),
            .I(\uart_pc.state_1_sqmuxa_0 ));
    Odrv4 I__2348 (
            .O(N__14583),
            .I(\uart_pc.state_1_sqmuxa_0 ));
    InMux I__2347 (
            .O(N__14576),
            .I(N__14573));
    LocalMux I__2346 (
            .O(N__14573),
            .I(N__14570));
    Odrv4 I__2345 (
            .O(N__14570),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__2344 (
            .O(N__14567),
            .I(N__14564));
    LocalMux I__2343 (
            .O(N__14564),
            .I(N__14561));
    Odrv4 I__2342 (
            .O(N__14561),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__2341 (
            .O(N__14558),
            .I(N__14555));
    LocalMux I__2340 (
            .O(N__14555),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__2339 (
            .O(N__14552),
            .I(N__14549));
    LocalMux I__2338 (
            .O(N__14549),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__2337 (
            .O(N__14546),
            .I(N__14543));
    LocalMux I__2336 (
            .O(N__14543),
            .I(N__14540));
    Odrv4 I__2335 (
            .O(N__14540),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    CascadeMux I__2334 (
            .O(N__14537),
            .I(N__14534));
    InMux I__2333 (
            .O(N__14534),
            .I(N__14531));
    LocalMux I__2332 (
            .O(N__14531),
            .I(N__14528));
    Odrv4 I__2331 (
            .O(N__14528),
            .I(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ));
    CascadeMux I__2330 (
            .O(N__14525),
            .I(N__14521));
    InMux I__2329 (
            .O(N__14524),
            .I(N__14516));
    InMux I__2328 (
            .O(N__14521),
            .I(N__14516));
    LocalMux I__2327 (
            .O(N__14516),
            .I(N__14506));
    InMux I__2326 (
            .O(N__14515),
            .I(N__14499));
    InMux I__2325 (
            .O(N__14514),
            .I(N__14499));
    InMux I__2324 (
            .O(N__14513),
            .I(N__14499));
    InMux I__2323 (
            .O(N__14512),
            .I(N__14490));
    InMux I__2322 (
            .O(N__14511),
            .I(N__14490));
    InMux I__2321 (
            .O(N__14510),
            .I(N__14490));
    InMux I__2320 (
            .O(N__14509),
            .I(N__14490));
    Odrv4 I__2319 (
            .O(N__14506),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__2318 (
            .O(N__14499),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__2317 (
            .O(N__14490),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    InMux I__2316 (
            .O(N__14483),
            .I(N__14480));
    LocalMux I__2315 (
            .O(N__14480),
            .I(N__14477));
    Odrv4 I__2314 (
            .O(N__14477),
            .I(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ));
    InMux I__2313 (
            .O(N__14474),
            .I(N__14471));
    LocalMux I__2312 (
            .O(N__14471),
            .I(N__14468));
    Odrv4 I__2311 (
            .O(N__14468),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    CascadeMux I__2310 (
            .O(N__14465),
            .I(\ppm_encoder_1.un1_init_pulses_0_2_cascade_ ));
    InMux I__2309 (
            .O(N__14462),
            .I(N__14459));
    LocalMux I__2308 (
            .O(N__14459),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2 ));
    InMux I__2307 (
            .O(N__14456),
            .I(N__14453));
    LocalMux I__2306 (
            .O(N__14453),
            .I(N__14450));
    Odrv4 I__2305 (
            .O(N__14450),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__2304 (
            .O(N__14447),
            .I(N__14444));
    LocalMux I__2303 (
            .O(N__14444),
            .I(N__14441));
    Span4Mux_v I__2302 (
            .O(N__14441),
            .I(N__14438));
    Odrv4 I__2301 (
            .O(N__14438),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__2300 (
            .O(N__14435),
            .I(N__14432));
    LocalMux I__2299 (
            .O(N__14432),
            .I(N__14429));
    Odrv4 I__2298 (
            .O(N__14429),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    CascadeMux I__2297 (
            .O(N__14426),
            .I(N__14423));
    InMux I__2296 (
            .O(N__14423),
            .I(N__14420));
    LocalMux I__2295 (
            .O(N__14420),
            .I(N__14417));
    Odrv4 I__2294 (
            .O(N__14417),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    CascadeMux I__2293 (
            .O(N__14414),
            .I(\ppm_encoder_1.PPM_STATE_62_d_cascade_ ));
    CascadeMux I__2292 (
            .O(N__14411),
            .I(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ));
    InMux I__2291 (
            .O(N__14408),
            .I(N__14405));
    LocalMux I__2290 (
            .O(N__14405),
            .I(N__14402));
    Span4Mux_v I__2289 (
            .O(N__14402),
            .I(N__14399));
    Odrv4 I__2288 (
            .O(N__14399),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    CascadeMux I__2287 (
            .O(N__14396),
            .I(N__14392));
    CascadeMux I__2286 (
            .O(N__14395),
            .I(N__14389));
    InMux I__2285 (
            .O(N__14392),
            .I(N__14386));
    InMux I__2284 (
            .O(N__14389),
            .I(N__14383));
    LocalMux I__2283 (
            .O(N__14386),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    LocalMux I__2282 (
            .O(N__14383),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    InMux I__2281 (
            .O(N__14378),
            .I(N__14375));
    LocalMux I__2280 (
            .O(N__14375),
            .I(N__14372));
    Odrv4 I__2279 (
            .O(N__14372),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    CascadeMux I__2278 (
            .O(N__14369),
            .I(N__14364));
    InMux I__2277 (
            .O(N__14368),
            .I(N__14361));
    InMux I__2276 (
            .O(N__14367),
            .I(N__14356));
    InMux I__2275 (
            .O(N__14364),
            .I(N__14356));
    LocalMux I__2274 (
            .O(N__14361),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__2273 (
            .O(N__14356),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__2272 (
            .O(N__14351),
            .I(N__14345));
    InMux I__2271 (
            .O(N__14350),
            .I(N__14338));
    InMux I__2270 (
            .O(N__14349),
            .I(N__14338));
    InMux I__2269 (
            .O(N__14348),
            .I(N__14338));
    LocalMux I__2268 (
            .O(N__14345),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__2267 (
            .O(N__14338),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    CascadeMux I__2266 (
            .O(N__14333),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ));
    CascadeMux I__2265 (
            .O(N__14330),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    InMux I__2264 (
            .O(N__14327),
            .I(N__14324));
    LocalMux I__2263 (
            .O(N__14324),
            .I(N__14321));
    Span4Mux_h I__2262 (
            .O(N__14321),
            .I(N__14318));
    Odrv4 I__2261 (
            .O(N__14318),
            .I(\ppm_encoder_1.N_299 ));
    InMux I__2260 (
            .O(N__14315),
            .I(\uart_frame_decoder.count8 ));
    CEMux I__2259 (
            .O(N__14312),
            .I(N__14309));
    LocalMux I__2258 (
            .O(N__14309),
            .I(N__14305));
    CEMux I__2257 (
            .O(N__14308),
            .I(N__14302));
    Span4Mux_v I__2256 (
            .O(N__14305),
            .I(N__14297));
    LocalMux I__2255 (
            .O(N__14302),
            .I(N__14297));
    Span4Mux_h I__2254 (
            .O(N__14297),
            .I(N__14294));
    Odrv4 I__2253 (
            .O(N__14294),
            .I(\uart_frame_decoder.source_CH1data_1_sqmuxa_0 ));
    InMux I__2252 (
            .O(N__14291),
            .I(\scaler_1.un3_source_data_0_cry_8 ));
    InMux I__2251 (
            .O(N__14288),
            .I(N__14285));
    LocalMux I__2250 (
            .O(N__14285),
            .I(\scaler_1.un3_source_data_0_axb_7 ));
    InMux I__2249 (
            .O(N__14282),
            .I(N__14276));
    InMux I__2248 (
            .O(N__14281),
            .I(N__14276));
    LocalMux I__2247 (
            .O(N__14276),
            .I(frame_decoder_CH1data_7));
    CascadeMux I__2246 (
            .O(N__14273),
            .I(N__14270));
    InMux I__2245 (
            .O(N__14270),
            .I(N__14264));
    InMux I__2244 (
            .O(N__14269),
            .I(N__14264));
    LocalMux I__2243 (
            .O(N__14264),
            .I(frame_decoder_OFF1data_7));
    InMux I__2242 (
            .O(N__14261),
            .I(N__14258));
    LocalMux I__2241 (
            .O(N__14258),
            .I(\scaler_1.N_508_i_l_ofxZ0 ));
    InMux I__2240 (
            .O(N__14255),
            .I(N__14249));
    InMux I__2239 (
            .O(N__14254),
            .I(N__14249));
    LocalMux I__2238 (
            .O(N__14249),
            .I(N__14246));
    Odrv4 I__2237 (
            .O(N__14246),
            .I(\uart_frame_decoder.count_RNIHJ501Z0Z_0 ));
    InMux I__2236 (
            .O(N__14243),
            .I(N__14240));
    LocalMux I__2235 (
            .O(N__14240),
            .I(\uart_frame_decoder.count8_axb_1 ));
    InMux I__2234 (
            .O(N__14237),
            .I(N__14234));
    LocalMux I__2233 (
            .O(N__14234),
            .I(\uart_frame_decoder.count_i_2 ));
    InMux I__2232 (
            .O(N__14231),
            .I(N__14228));
    LocalMux I__2231 (
            .O(N__14228),
            .I(frame_decoder_CH1data_1));
    CascadeMux I__2230 (
            .O(N__14225),
            .I(N__14222));
    InMux I__2229 (
            .O(N__14222),
            .I(N__14219));
    LocalMux I__2228 (
            .O(N__14219),
            .I(frame_decoder_OFF1data_1));
    InMux I__2227 (
            .O(N__14216),
            .I(\scaler_1.un3_source_data_0_cry_0 ));
    InMux I__2226 (
            .O(N__14213),
            .I(N__14210));
    LocalMux I__2225 (
            .O(N__14210),
            .I(frame_decoder_CH1data_2));
    CascadeMux I__2224 (
            .O(N__14207),
            .I(N__14204));
    InMux I__2223 (
            .O(N__14204),
            .I(N__14201));
    LocalMux I__2222 (
            .O(N__14201),
            .I(frame_decoder_OFF1data_2));
    InMux I__2221 (
            .O(N__14198),
            .I(\scaler_1.un3_source_data_0_cry_1 ));
    InMux I__2220 (
            .O(N__14195),
            .I(N__14192));
    LocalMux I__2219 (
            .O(N__14192),
            .I(frame_decoder_CH1data_3));
    CascadeMux I__2218 (
            .O(N__14189),
            .I(N__14186));
    InMux I__2217 (
            .O(N__14186),
            .I(N__14183));
    LocalMux I__2216 (
            .O(N__14183),
            .I(frame_decoder_OFF1data_3));
    InMux I__2215 (
            .O(N__14180),
            .I(\scaler_1.un3_source_data_0_cry_2 ));
    InMux I__2214 (
            .O(N__14177),
            .I(N__14174));
    LocalMux I__2213 (
            .O(N__14174),
            .I(frame_decoder_CH1data_4));
    CascadeMux I__2212 (
            .O(N__14171),
            .I(N__14168));
    InMux I__2211 (
            .O(N__14168),
            .I(N__14165));
    LocalMux I__2210 (
            .O(N__14165),
            .I(frame_decoder_OFF1data_4));
    InMux I__2209 (
            .O(N__14162),
            .I(\scaler_1.un3_source_data_0_cry_3 ));
    InMux I__2208 (
            .O(N__14159),
            .I(N__14156));
    LocalMux I__2207 (
            .O(N__14156),
            .I(frame_decoder_CH1data_5));
    CascadeMux I__2206 (
            .O(N__14153),
            .I(N__14150));
    InMux I__2205 (
            .O(N__14150),
            .I(N__14147));
    LocalMux I__2204 (
            .O(N__14147),
            .I(frame_decoder_OFF1data_5));
    InMux I__2203 (
            .O(N__14144),
            .I(\scaler_1.un3_source_data_0_cry_4 ));
    InMux I__2202 (
            .O(N__14141),
            .I(N__14138));
    LocalMux I__2201 (
            .O(N__14138),
            .I(frame_decoder_CH1data_6));
    CascadeMux I__2200 (
            .O(N__14135),
            .I(N__14132));
    InMux I__2199 (
            .O(N__14132),
            .I(N__14129));
    LocalMux I__2198 (
            .O(N__14129),
            .I(frame_decoder_OFF1data_6));
    InMux I__2197 (
            .O(N__14126),
            .I(\scaler_1.un3_source_data_0_cry_5 ));
    InMux I__2196 (
            .O(N__14123),
            .I(\scaler_1.un3_source_data_0_cry_6 ));
    InMux I__2195 (
            .O(N__14120),
            .I(bfn_8_18_0_));
    CEMux I__2194 (
            .O(N__14117),
            .I(N__14114));
    LocalMux I__2193 (
            .O(N__14114),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    InMux I__2192 (
            .O(N__14111),
            .I(N__14107));
    InMux I__2191 (
            .O(N__14110),
            .I(N__14104));
    LocalMux I__2190 (
            .O(N__14107),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__2189 (
            .O(N__14104),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    InMux I__2188 (
            .O(N__14099),
            .I(N__14094));
    InMux I__2187 (
            .O(N__14098),
            .I(N__14089));
    InMux I__2186 (
            .O(N__14097),
            .I(N__14089));
    LocalMux I__2185 (
            .O(N__14094),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__2184 (
            .O(N__14089),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    InMux I__2183 (
            .O(N__14084),
            .I(N__14080));
    InMux I__2182 (
            .O(N__14083),
            .I(N__14077));
    LocalMux I__2181 (
            .O(N__14080),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__2180 (
            .O(N__14077),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    CascadeMux I__2179 (
            .O(N__14072),
            .I(N__14068));
    InMux I__2178 (
            .O(N__14071),
            .I(N__14065));
    InMux I__2177 (
            .O(N__14068),
            .I(N__14062));
    LocalMux I__2176 (
            .O(N__14065),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__2175 (
            .O(N__14062),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    InMux I__2174 (
            .O(N__14057),
            .I(N__14052));
    InMux I__2173 (
            .O(N__14056),
            .I(N__14047));
    InMux I__2172 (
            .O(N__14055),
            .I(N__14047));
    LocalMux I__2171 (
            .O(N__14052),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__2170 (
            .O(N__14047),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    InMux I__2169 (
            .O(N__14042),
            .I(N__14038));
    InMux I__2168 (
            .O(N__14041),
            .I(N__14035));
    LocalMux I__2167 (
            .O(N__14038),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__2166 (
            .O(N__14035),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    CascadeMux I__2165 (
            .O(N__14030),
            .I(\uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ));
    InMux I__2164 (
            .O(N__14027),
            .I(N__14024));
    LocalMux I__2163 (
            .O(N__14024),
            .I(\uart_frame_decoder.WDT8lto13_1 ));
    InMux I__2162 (
            .O(N__14021),
            .I(N__14018));
    LocalMux I__2161 (
            .O(N__14018),
            .I(N__14015));
    Odrv4 I__2160 (
            .O(N__14015),
            .I(\uart_frame_decoder.WDT8lt14_0 ));
    InMux I__2159 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__2158 (
            .O(N__14009),
            .I(N__14005));
    InMux I__2157 (
            .O(N__14008),
            .I(N__14001));
    Span4Mux_h I__2156 (
            .O(N__14005),
            .I(N__13998));
    InMux I__2155 (
            .O(N__14004),
            .I(N__13995));
    LocalMux I__2154 (
            .O(N__14001),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__2153 (
            .O(N__13998),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__2152 (
            .O(N__13995),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    CascadeMux I__2151 (
            .O(N__13988),
            .I(\uart_frame_decoder.WDT8lt14_0_cascade_ ));
    InMux I__2150 (
            .O(N__13985),
            .I(N__13982));
    LocalMux I__2149 (
            .O(N__13982),
            .I(N__13978));
    InMux I__2148 (
            .O(N__13981),
            .I(N__13974));
    Span4Mux_h I__2147 (
            .O(N__13978),
            .I(N__13971));
    InMux I__2146 (
            .O(N__13977),
            .I(N__13968));
    LocalMux I__2145 (
            .O(N__13974),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__2144 (
            .O(N__13971),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__2143 (
            .O(N__13968),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    CascadeMux I__2142 (
            .O(N__13961),
            .I(N__13957));
    InMux I__2141 (
            .O(N__13960),
            .I(N__13954));
    InMux I__2140 (
            .O(N__13957),
            .I(N__13951));
    LocalMux I__2139 (
            .O(N__13954),
            .I(\uart_frame_decoder.WDT8_0_i ));
    LocalMux I__2138 (
            .O(N__13951),
            .I(\uart_frame_decoder.WDT8_0_i ));
    InMux I__2137 (
            .O(N__13946),
            .I(N__13942));
    InMux I__2136 (
            .O(N__13945),
            .I(N__13939));
    LocalMux I__2135 (
            .O(N__13942),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__2134 (
            .O(N__13939),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    InMux I__2133 (
            .O(N__13934),
            .I(N__13930));
    InMux I__2132 (
            .O(N__13933),
            .I(N__13927));
    LocalMux I__2131 (
            .O(N__13930),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__2130 (
            .O(N__13927),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    CascadeMux I__2129 (
            .O(N__13922),
            .I(N__13918));
    InMux I__2128 (
            .O(N__13921),
            .I(N__13915));
    InMux I__2127 (
            .O(N__13918),
            .I(N__13912));
    LocalMux I__2126 (
            .O(N__13915),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__2125 (
            .O(N__13912),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    InMux I__2124 (
            .O(N__13907),
            .I(N__13903));
    InMux I__2123 (
            .O(N__13906),
            .I(N__13900));
    LocalMux I__2122 (
            .O(N__13903),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__2121 (
            .O(N__13900),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    InMux I__2120 (
            .O(N__13895),
            .I(N__13892));
    LocalMux I__2119 (
            .O(N__13892),
            .I(\uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ));
    SRMux I__2118 (
            .O(N__13889),
            .I(N__13886));
    LocalMux I__2117 (
            .O(N__13886),
            .I(N__13882));
    SRMux I__2116 (
            .O(N__13885),
            .I(N__13879));
    Span4Mux_h I__2115 (
            .O(N__13882),
            .I(N__13876));
    LocalMux I__2114 (
            .O(N__13879),
            .I(N__13873));
    Odrv4 I__2113 (
            .O(N__13876),
            .I(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ));
    Odrv4 I__2112 (
            .O(N__13873),
            .I(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ));
    CEMux I__2111 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__2110 (
            .O(N__13865),
            .I(N__13862));
    Span4Mux_h I__2109 (
            .O(N__13862),
            .I(N__13859));
    Span4Mux_h I__2108 (
            .O(N__13859),
            .I(N__13856));
    Odrv4 I__2107 (
            .O(N__13856),
            .I(\uart_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    InMux I__2106 (
            .O(N__13853),
            .I(N__13849));
    InMux I__2105 (
            .O(N__13852),
            .I(N__13846));
    LocalMux I__2104 (
            .O(N__13849),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    LocalMux I__2103 (
            .O(N__13846),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    InMux I__2102 (
            .O(N__13841),
            .I(N__13837));
    InMux I__2101 (
            .O(N__13840),
            .I(N__13834));
    LocalMux I__2100 (
            .O(N__13837),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa ));
    LocalMux I__2099 (
            .O(N__13834),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa ));
    InMux I__2098 (
            .O(N__13829),
            .I(N__13825));
    InMux I__2097 (
            .O(N__13828),
            .I(N__13822));
    LocalMux I__2096 (
            .O(N__13825),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    LocalMux I__2095 (
            .O(N__13822),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    InMux I__2094 (
            .O(N__13817),
            .I(N__13814));
    LocalMux I__2093 (
            .O(N__13814),
            .I(N__13811));
    Odrv4 I__2092 (
            .O(N__13811),
            .I(\uart_frame_decoder.source_offset2data_1_sqmuxa ));
    InMux I__2091 (
            .O(N__13808),
            .I(N__13804));
    InMux I__2090 (
            .O(N__13807),
            .I(N__13801));
    LocalMux I__2089 (
            .O(N__13804),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    LocalMux I__2088 (
            .O(N__13801),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    CascadeMux I__2087 (
            .O(N__13796),
            .I(N__13793));
    InMux I__2086 (
            .O(N__13793),
            .I(N__13789));
    InMux I__2085 (
            .O(N__13792),
            .I(N__13786));
    LocalMux I__2084 (
            .O(N__13789),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa ));
    LocalMux I__2083 (
            .O(N__13786),
            .I(\uart_frame_decoder.source_offset3data_1_sqmuxa ));
    InMux I__2082 (
            .O(N__13781),
            .I(N__13778));
    LocalMux I__2081 (
            .O(N__13778),
            .I(\uart_frame_decoder.N_138_4 ));
    CascadeMux I__2080 (
            .O(N__13775),
            .I(\uart_frame_decoder.N_138_4_cascade_ ));
    CascadeMux I__2079 (
            .O(N__13772),
            .I(N__13769));
    InMux I__2078 (
            .O(N__13769),
            .I(N__13766));
    LocalMux I__2077 (
            .O(N__13766),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ));
    InMux I__2076 (
            .O(N__13763),
            .I(N__13756));
    InMux I__2075 (
            .O(N__13762),
            .I(N__13749));
    InMux I__2074 (
            .O(N__13761),
            .I(N__13749));
    InMux I__2073 (
            .O(N__13760),
            .I(N__13749));
    InMux I__2072 (
            .O(N__13759),
            .I(N__13746));
    LocalMux I__2071 (
            .O(N__13756),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__2070 (
            .O(N__13749),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__2069 (
            .O(N__13746),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    InMux I__2068 (
            .O(N__13739),
            .I(N__13736));
    LocalMux I__2067 (
            .O(N__13736),
            .I(\uart_frame_decoder.state_1_RNO_2Z0Z_0 ));
    CascadeMux I__2066 (
            .O(N__13733),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ));
    CascadeMux I__2065 (
            .O(N__13730),
            .I(\uart_frame_decoder.N_85_cascade_ ));
    InMux I__2064 (
            .O(N__13727),
            .I(N__13724));
    LocalMux I__2063 (
            .O(N__13724),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__2062 (
            .O(N__13721),
            .I(N__13718));
    LocalMux I__2061 (
            .O(N__13718),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__2060 (
            .O(N__13715),
            .I(N__13712));
    LocalMux I__2059 (
            .O(N__13712),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__2058 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__2057 (
            .O(N__13706),
            .I(N__13703));
    Odrv12 I__2056 (
            .O(N__13703),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    CascadeMux I__2055 (
            .O(N__13700),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ));
    CascadeMux I__2054 (
            .O(N__13697),
            .I(\uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_ ));
    CascadeMux I__2053 (
            .O(N__13694),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ));
    InMux I__2052 (
            .O(N__13691),
            .I(N__13688));
    LocalMux I__2051 (
            .O(N__13688),
            .I(N__13685));
    Span4Mux_v I__2050 (
            .O(N__13685),
            .I(N__13682));
    Odrv4 I__2049 (
            .O(N__13682),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__2048 (
            .O(N__13679),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__2047 (
            .O(N__13676),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__2046 (
            .O(N__13673),
            .I(bfn_7_28_0_));
    InMux I__2045 (
            .O(N__13670),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__2044 (
            .O(N__13667),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__2043 (
            .O(N__13664),
            .I(N__13661));
    LocalMux I__2042 (
            .O(N__13661),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__2041 (
            .O(N__13658),
            .I(N__13655));
    LocalMux I__2040 (
            .O(N__13655),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__2039 (
            .O(N__13652),
            .I(N__13649));
    LocalMux I__2038 (
            .O(N__13649),
            .I(N__13646));
    Odrv4 I__2037 (
            .O(N__13646),
            .I(uart_input_pc_c));
    InMux I__2036 (
            .O(N__13643),
            .I(N__13640));
    LocalMux I__2035 (
            .O(N__13640),
            .I(N__13637));
    Odrv12 I__2034 (
            .O(N__13637),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ));
    CascadeMux I__2033 (
            .O(N__13634),
            .I(N__13631));
    InMux I__2032 (
            .O(N__13631),
            .I(N__13628));
    LocalMux I__2031 (
            .O(N__13628),
            .I(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ));
    CascadeMux I__2030 (
            .O(N__13625),
            .I(N__13622));
    InMux I__2029 (
            .O(N__13622),
            .I(N__13619));
    LocalMux I__2028 (
            .O(N__13619),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__2027 (
            .O(N__13616),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__2026 (
            .O(N__13613),
            .I(N__13610));
    LocalMux I__2025 (
            .O(N__13610),
            .I(N__13607));
    Odrv12 I__2024 (
            .O(N__13607),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__2023 (
            .O(N__13604),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__2022 (
            .O(N__13601),
            .I(bfn_7_27_0_));
    InMux I__2021 (
            .O(N__13598),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__2020 (
            .O(N__13595),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__2019 (
            .O(N__13592),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__2018 (
            .O(N__13589),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__2017 (
            .O(N__13586),
            .I(N__13583));
    LocalMux I__2016 (
            .O(N__13583),
            .I(N__13580));
    Odrv12 I__2015 (
            .O(N__13580),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ));
    CascadeMux I__2014 (
            .O(N__13577),
            .I(N__13574));
    InMux I__2013 (
            .O(N__13574),
            .I(N__13571));
    LocalMux I__2012 (
            .O(N__13571),
            .I(N__13568));
    Odrv4 I__2011 (
            .O(N__13568),
            .I(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ));
    InMux I__2010 (
            .O(N__13565),
            .I(N__13562));
    LocalMux I__2009 (
            .O(N__13562),
            .I(N__13559));
    Odrv4 I__2008 (
            .O(N__13559),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__2007 (
            .O(N__13556),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__2006 (
            .O(N__13553),
            .I(N__13550));
    LocalMux I__2005 (
            .O(N__13550),
            .I(N__13547));
    Odrv4 I__2004 (
            .O(N__13547),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ));
    InMux I__2003 (
            .O(N__13544),
            .I(N__13541));
    LocalMux I__2002 (
            .O(N__13541),
            .I(N__13538));
    Odrv12 I__2001 (
            .O(N__13538),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__2000 (
            .O(N__13535),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    CascadeMux I__1999 (
            .O(N__13532),
            .I(N__13529));
    InMux I__1998 (
            .O(N__13529),
            .I(N__13526));
    LocalMux I__1997 (
            .O(N__13526),
            .I(N__13523));
    Odrv4 I__1996 (
            .O(N__13523),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ));
    InMux I__1995 (
            .O(N__13520),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__1994 (
            .O(N__13517),
            .I(N__13514));
    LocalMux I__1993 (
            .O(N__13514),
            .I(N__13511));
    Odrv4 I__1992 (
            .O(N__13511),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__1991 (
            .O(N__13508),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__1990 (
            .O(N__13505),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__1989 (
            .O(N__13502),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    CascadeMux I__1988 (
            .O(N__13499),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    InMux I__1987 (
            .O(N__13496),
            .I(N__13487));
    InMux I__1986 (
            .O(N__13495),
            .I(N__13487));
    InMux I__1985 (
            .O(N__13494),
            .I(N__13487));
    LocalMux I__1984 (
            .O(N__13487),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    CascadeMux I__1983 (
            .O(N__13484),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ));
    CascadeMux I__1982 (
            .O(N__13481),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ));
    CascadeMux I__1981 (
            .O(N__13478),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ));
    CEMux I__1980 (
            .O(N__13475),
            .I(N__13472));
    LocalMux I__1979 (
            .O(N__13472),
            .I(N__13469));
    Span4Mux_v I__1978 (
            .O(N__13469),
            .I(N__13466));
    Odrv4 I__1977 (
            .O(N__13466),
            .I(\uart_frame_decoder.source_offset1data_1_sqmuxa_0 ));
    InMux I__1976 (
            .O(N__13463),
            .I(\uart_frame_decoder.un1_WDT_cry_10 ));
    InMux I__1975 (
            .O(N__13460),
            .I(\uart_frame_decoder.un1_WDT_cry_11 ));
    InMux I__1974 (
            .O(N__13457),
            .I(\uart_frame_decoder.un1_WDT_cry_12 ));
    InMux I__1973 (
            .O(N__13454),
            .I(\uart_frame_decoder.un1_WDT_cry_13 ));
    InMux I__1972 (
            .O(N__13451),
            .I(\uart_frame_decoder.un1_WDT_cry_14 ));
    InMux I__1971 (
            .O(N__13448),
            .I(\uart_frame_decoder.un1_WDT_cry_1 ));
    InMux I__1970 (
            .O(N__13445),
            .I(N__13442));
    LocalMux I__1969 (
            .O(N__13442),
            .I(\uart_frame_decoder.WDTZ0Z_3 ));
    InMux I__1968 (
            .O(N__13439),
            .I(\uart_frame_decoder.un1_WDT_cry_2 ));
    InMux I__1967 (
            .O(N__13436),
            .I(\uart_frame_decoder.un1_WDT_cry_3 ));
    InMux I__1966 (
            .O(N__13433),
            .I(\uart_frame_decoder.un1_WDT_cry_4 ));
    InMux I__1965 (
            .O(N__13430),
            .I(\uart_frame_decoder.un1_WDT_cry_5 ));
    InMux I__1964 (
            .O(N__13427),
            .I(\uart_frame_decoder.un1_WDT_cry_6 ));
    InMux I__1963 (
            .O(N__13424),
            .I(bfn_7_16_0_));
    InMux I__1962 (
            .O(N__13421),
            .I(\uart_frame_decoder.un1_WDT_cry_8 ));
    InMux I__1961 (
            .O(N__13418),
            .I(\uart_frame_decoder.un1_WDT_cry_9 ));
    CascadeMux I__1960 (
            .O(N__13415),
            .I(\uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ));
    InMux I__1959 (
            .O(N__13412),
            .I(N__13409));
    LocalMux I__1958 (
            .O(N__13409),
            .I(\uart_frame_decoder.WDTZ0Z_0 ));
    InMux I__1957 (
            .O(N__13406),
            .I(N__13403));
    LocalMux I__1956 (
            .O(N__13403),
            .I(\uart_frame_decoder.WDTZ0Z_1 ));
    InMux I__1955 (
            .O(N__13400),
            .I(\uart_frame_decoder.un1_WDT_cry_0 ));
    InMux I__1954 (
            .O(N__13397),
            .I(N__13394));
    LocalMux I__1953 (
            .O(N__13394),
            .I(\uart_frame_decoder.WDTZ0Z_2 ));
    InMux I__1952 (
            .O(N__13391),
            .I(N__13388));
    LocalMux I__1951 (
            .O(N__13388),
            .I(uart_input_drone_c));
    InMux I__1950 (
            .O(N__13385),
            .I(N__13382));
    LocalMux I__1949 (
            .O(N__13382),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__1948 (
            .O(N__13379),
            .I(N__13376));
    LocalMux I__1947 (
            .O(N__13376),
            .I(N__13373));
    Odrv4 I__1946 (
            .O(N__13373),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__1945 (
            .O(N__13370),
            .I(N__13367));
    LocalMux I__1944 (
            .O(N__13367),
            .I(N__13364));
    Span4Mux_v I__1943 (
            .O(N__13364),
            .I(N__13360));
    InMux I__1942 (
            .O(N__13363),
            .I(N__13357));
    Odrv4 I__1941 (
            .O(N__13360),
            .I(\uart_pc.data_AuxZ0Z_1 ));
    LocalMux I__1940 (
            .O(N__13357),
            .I(\uart_pc.data_AuxZ0Z_1 ));
    InMux I__1939 (
            .O(N__13352),
            .I(N__13349));
    LocalMux I__1938 (
            .O(N__13349),
            .I(N__13345));
    CascadeMux I__1937 (
            .O(N__13348),
            .I(N__13342));
    Span4Mux_v I__1936 (
            .O(N__13345),
            .I(N__13339));
    InMux I__1935 (
            .O(N__13342),
            .I(N__13336));
    Odrv4 I__1934 (
            .O(N__13339),
            .I(\uart_pc.data_AuxZ0Z_0 ));
    LocalMux I__1933 (
            .O(N__13336),
            .I(\uart_pc.data_AuxZ0Z_0 ));
    CascadeMux I__1932 (
            .O(N__13331),
            .I(N__13328));
    InMux I__1931 (
            .O(N__13328),
            .I(N__13324));
    InMux I__1930 (
            .O(N__13327),
            .I(N__13321));
    LocalMux I__1929 (
            .O(N__13324),
            .I(N__13318));
    LocalMux I__1928 (
            .O(N__13321),
            .I(N__13315));
    Odrv4 I__1927 (
            .O(N__13318),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    Odrv4 I__1926 (
            .O(N__13315),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__1925 (
            .O(N__13310),
            .I(N__13306));
    CascadeMux I__1924 (
            .O(N__13309),
            .I(N__13303));
    LocalMux I__1923 (
            .O(N__13306),
            .I(N__13300));
    InMux I__1922 (
            .O(N__13303),
            .I(N__13297));
    Odrv4 I__1921 (
            .O(N__13300),
            .I(\uart_pc.data_AuxZ0Z_2 ));
    LocalMux I__1920 (
            .O(N__13297),
            .I(\uart_pc.data_AuxZ0Z_2 ));
    InMux I__1919 (
            .O(N__13292),
            .I(N__13289));
    LocalMux I__1918 (
            .O(N__13289),
            .I(N__13285));
    InMux I__1917 (
            .O(N__13288),
            .I(N__13282));
    Odrv4 I__1916 (
            .O(N__13285),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__1915 (
            .O(N__13282),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__1914 (
            .O(N__13277),
            .I(N__13274));
    LocalMux I__1913 (
            .O(N__13274),
            .I(N__13270));
    InMux I__1912 (
            .O(N__13273),
            .I(N__13267));
    Odrv4 I__1911 (
            .O(N__13270),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__1910 (
            .O(N__13267),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    InMux I__1909 (
            .O(N__13262),
            .I(N__13258));
    InMux I__1908 (
            .O(N__13261),
            .I(N__13255));
    LocalMux I__1907 (
            .O(N__13258),
            .I(N__13250));
    LocalMux I__1906 (
            .O(N__13255),
            .I(N__13250));
    Odrv4 I__1905 (
            .O(N__13250),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    CascadeMux I__1904 (
            .O(N__13247),
            .I(\uart_pc.N_143_cascade_ ));
    InMux I__1903 (
            .O(N__13244),
            .I(N__13241));
    LocalMux I__1902 (
            .O(N__13241),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1 ));
    InMux I__1901 (
            .O(N__13238),
            .I(N__13234));
    InMux I__1900 (
            .O(N__13237),
            .I(N__13231));
    LocalMux I__1899 (
            .O(N__13234),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__1898 (
            .O(N__13231),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    CascadeMux I__1897 (
            .O(N__13226),
            .I(N__13220));
    InMux I__1896 (
            .O(N__13225),
            .I(N__13215));
    InMux I__1895 (
            .O(N__13224),
            .I(N__13215));
    InMux I__1894 (
            .O(N__13223),
            .I(N__13210));
    InMux I__1893 (
            .O(N__13220),
            .I(N__13210));
    LocalMux I__1892 (
            .O(N__13215),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__1891 (
            .O(N__13210),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    CascadeMux I__1890 (
            .O(N__13205),
            .I(N__13202));
    InMux I__1889 (
            .O(N__13202),
            .I(N__13199));
    LocalMux I__1888 (
            .O(N__13199),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__1887 (
            .O(N__13196),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__1886 (
            .O(N__13193),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__1885 (
            .O(N__13190),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    CascadeMux I__1884 (
            .O(N__13187),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ));
    InMux I__1883 (
            .O(N__13184),
            .I(N__13178));
    InMux I__1882 (
            .O(N__13183),
            .I(N__13175));
    CascadeMux I__1881 (
            .O(N__13182),
            .I(N__13170));
    CascadeMux I__1880 (
            .O(N__13181),
            .I(N__13166));
    LocalMux I__1879 (
            .O(N__13178),
            .I(N__13160));
    LocalMux I__1878 (
            .O(N__13175),
            .I(N__13160));
    InMux I__1877 (
            .O(N__13174),
            .I(N__13156));
    InMux I__1876 (
            .O(N__13173),
            .I(N__13147));
    InMux I__1875 (
            .O(N__13170),
            .I(N__13147));
    InMux I__1874 (
            .O(N__13169),
            .I(N__13147));
    InMux I__1873 (
            .O(N__13166),
            .I(N__13147));
    InMux I__1872 (
            .O(N__13165),
            .I(N__13144));
    Span4Mux_v I__1871 (
            .O(N__13160),
            .I(N__13141));
    InMux I__1870 (
            .O(N__13159),
            .I(N__13138));
    LocalMux I__1869 (
            .O(N__13156),
            .I(N__13133));
    LocalMux I__1868 (
            .O(N__13147),
            .I(N__13133));
    LocalMux I__1867 (
            .O(N__13144),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__1866 (
            .O(N__13141),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__1865 (
            .O(N__13138),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv12 I__1864 (
            .O(N__13133),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__1863 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__1862 (
            .O(N__13121),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    InMux I__1861 (
            .O(N__13118),
            .I(N__13113));
    InMux I__1860 (
            .O(N__13117),
            .I(N__13110));
    InMux I__1859 (
            .O(N__13116),
            .I(N__13107));
    LocalMux I__1858 (
            .O(N__13113),
            .I(N__13104));
    LocalMux I__1857 (
            .O(N__13110),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__1856 (
            .O(N__13107),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    Odrv4 I__1855 (
            .O(N__13104),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__1854 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__1853 (
            .O(N__13094),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    InMux I__1852 (
            .O(N__13091),
            .I(N__13084));
    InMux I__1851 (
            .O(N__13090),
            .I(N__13081));
    InMux I__1850 (
            .O(N__13089),
            .I(N__13076));
    InMux I__1849 (
            .O(N__13088),
            .I(N__13076));
    InMux I__1848 (
            .O(N__13087),
            .I(N__13073));
    LocalMux I__1847 (
            .O(N__13084),
            .I(\uart_pc.N_143 ));
    LocalMux I__1846 (
            .O(N__13081),
            .I(\uart_pc.N_143 ));
    LocalMux I__1845 (
            .O(N__13076),
            .I(\uart_pc.N_143 ));
    LocalMux I__1844 (
            .O(N__13073),
            .I(\uart_pc.N_143 ));
    InMux I__1843 (
            .O(N__13064),
            .I(N__13055));
    InMux I__1842 (
            .O(N__13063),
            .I(N__13055));
    InMux I__1841 (
            .O(N__13062),
            .I(N__13055));
    LocalMux I__1840 (
            .O(N__13055),
            .I(N__13050));
    InMux I__1839 (
            .O(N__13054),
            .I(N__13045));
    InMux I__1838 (
            .O(N__13053),
            .I(N__13045));
    Odrv12 I__1837 (
            .O(N__13050),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__1836 (
            .O(N__13045),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__1835 (
            .O(N__13040),
            .I(N__13036));
    InMux I__1834 (
            .O(N__13039),
            .I(N__13027));
    LocalMux I__1833 (
            .O(N__13036),
            .I(N__13024));
    InMux I__1832 (
            .O(N__13035),
            .I(N__13015));
    InMux I__1831 (
            .O(N__13034),
            .I(N__13015));
    InMux I__1830 (
            .O(N__13033),
            .I(N__13015));
    InMux I__1829 (
            .O(N__13032),
            .I(N__13015));
    InMux I__1828 (
            .O(N__13031),
            .I(N__13012));
    InMux I__1827 (
            .O(N__13030),
            .I(N__13009));
    LocalMux I__1826 (
            .O(N__13027),
            .I(N__13006));
    Span4Mux_v I__1825 (
            .O(N__13024),
            .I(N__13001));
    LocalMux I__1824 (
            .O(N__13015),
            .I(N__13001));
    LocalMux I__1823 (
            .O(N__13012),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__1822 (
            .O(N__13009),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv12 I__1821 (
            .O(N__13006),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__1820 (
            .O(N__13001),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    CascadeMux I__1819 (
            .O(N__12992),
            .I(\uart_pc.N_145_cascade_ ));
    CascadeMux I__1818 (
            .O(N__12989),
            .I(N__12984));
    CascadeMux I__1817 (
            .O(N__12988),
            .I(N__12981));
    InMux I__1816 (
            .O(N__12987),
            .I(N__12977));
    InMux I__1815 (
            .O(N__12984),
            .I(N__12972));
    InMux I__1814 (
            .O(N__12981),
            .I(N__12972));
    InMux I__1813 (
            .O(N__12980),
            .I(N__12969));
    LocalMux I__1812 (
            .O(N__12977),
            .I(N__12964));
    LocalMux I__1811 (
            .O(N__12972),
            .I(N__12964));
    LocalMux I__1810 (
            .O(N__12969),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__1809 (
            .O(N__12964),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__1808 (
            .O(N__12959),
            .I(N__12954));
    InMux I__1807 (
            .O(N__12958),
            .I(N__12951));
    InMux I__1806 (
            .O(N__12957),
            .I(N__12947));
    LocalMux I__1805 (
            .O(N__12954),
            .I(N__12944));
    LocalMux I__1804 (
            .O(N__12951),
            .I(N__12941));
    InMux I__1803 (
            .O(N__12950),
            .I(N__12938));
    LocalMux I__1802 (
            .O(N__12947),
            .I(\uart_pc.N_152 ));
    Odrv4 I__1801 (
            .O(N__12944),
            .I(\uart_pc.N_152 ));
    Odrv4 I__1800 (
            .O(N__12941),
            .I(\uart_pc.N_152 ));
    LocalMux I__1799 (
            .O(N__12938),
            .I(\uart_pc.N_152 ));
    InMux I__1798 (
            .O(N__12929),
            .I(N__12923));
    InMux I__1797 (
            .O(N__12928),
            .I(N__12923));
    LocalMux I__1796 (
            .O(N__12923),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__1795 (
            .O(N__12920),
            .I(N__12913));
    InMux I__1794 (
            .O(N__12919),
            .I(N__12910));
    CascadeMux I__1793 (
            .O(N__12918),
            .I(N__12906));
    InMux I__1792 (
            .O(N__12917),
            .I(N__12901));
    InMux I__1791 (
            .O(N__12916),
            .I(N__12896));
    InMux I__1790 (
            .O(N__12913),
            .I(N__12896));
    LocalMux I__1789 (
            .O(N__12910),
            .I(N__12893));
    InMux I__1788 (
            .O(N__12909),
            .I(N__12890));
    InMux I__1787 (
            .O(N__12906),
            .I(N__12883));
    InMux I__1786 (
            .O(N__12905),
            .I(N__12883));
    InMux I__1785 (
            .O(N__12904),
            .I(N__12883));
    LocalMux I__1784 (
            .O(N__12901),
            .I(N__12878));
    LocalMux I__1783 (
            .O(N__12896),
            .I(N__12878));
    Odrv12 I__1782 (
            .O(N__12893),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__1781 (
            .O(N__12890),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__1780 (
            .O(N__12883),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__1779 (
            .O(N__12878),
            .I(\uart_pc.stateZ0Z_3 ));
    InMux I__1778 (
            .O(N__12869),
            .I(N__12859));
    InMux I__1777 (
            .O(N__12868),
            .I(N__12844));
    InMux I__1776 (
            .O(N__12867),
            .I(N__12844));
    InMux I__1775 (
            .O(N__12866),
            .I(N__12844));
    InMux I__1774 (
            .O(N__12865),
            .I(N__12844));
    InMux I__1773 (
            .O(N__12864),
            .I(N__12844));
    InMux I__1772 (
            .O(N__12863),
            .I(N__12844));
    InMux I__1771 (
            .O(N__12862),
            .I(N__12844));
    LocalMux I__1770 (
            .O(N__12859),
            .I(N__12839));
    LocalMux I__1769 (
            .O(N__12844),
            .I(N__12839));
    Odrv12 I__1768 (
            .O(N__12839),
            .I(\uart_pc.un1_state_2_0 ));
    CascadeMux I__1767 (
            .O(N__12836),
            .I(N__12833));
    InMux I__1766 (
            .O(N__12833),
            .I(N__12830));
    LocalMux I__1765 (
            .O(N__12830),
            .I(N__12826));
    InMux I__1764 (
            .O(N__12829),
            .I(N__12823));
    Odrv4 I__1763 (
            .O(N__12826),
            .I(\uart_pc.N_126_li ));
    LocalMux I__1762 (
            .O(N__12823),
            .I(\uart_pc.N_126_li ));
    InMux I__1761 (
            .O(N__12818),
            .I(N__12813));
    InMux I__1760 (
            .O(N__12817),
            .I(N__12808));
    InMux I__1759 (
            .O(N__12816),
            .I(N__12804));
    LocalMux I__1758 (
            .O(N__12813),
            .I(N__12801));
    InMux I__1757 (
            .O(N__12812),
            .I(N__12796));
    InMux I__1756 (
            .O(N__12811),
            .I(N__12796));
    LocalMux I__1755 (
            .O(N__12808),
            .I(N__12793));
    InMux I__1754 (
            .O(N__12807),
            .I(N__12790));
    LocalMux I__1753 (
            .O(N__12804),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv12 I__1752 (
            .O(N__12801),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__1751 (
            .O(N__12796),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv4 I__1750 (
            .O(N__12793),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__1749 (
            .O(N__12790),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__1748 (
            .O(N__12779),
            .I(\uart_pc.N_126_li_cascade_ ));
    InMux I__1747 (
            .O(N__12776),
            .I(N__12773));
    LocalMux I__1746 (
            .O(N__12773),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__1745 (
            .O(N__12770),
            .I(N__12765));
    InMux I__1744 (
            .O(N__12769),
            .I(N__12760));
    InMux I__1743 (
            .O(N__12768),
            .I(N__12760));
    InMux I__1742 (
            .O(N__12765),
            .I(N__12751));
    LocalMux I__1741 (
            .O(N__12760),
            .I(N__12748));
    InMux I__1740 (
            .O(N__12759),
            .I(N__12737));
    InMux I__1739 (
            .O(N__12758),
            .I(N__12737));
    InMux I__1738 (
            .O(N__12757),
            .I(N__12737));
    InMux I__1737 (
            .O(N__12756),
            .I(N__12737));
    InMux I__1736 (
            .O(N__12755),
            .I(N__12737));
    InMux I__1735 (
            .O(N__12754),
            .I(N__12734));
    LocalMux I__1734 (
            .O(N__12751),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    Odrv4 I__1733 (
            .O(N__12748),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__1732 (
            .O(N__12737),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__1731 (
            .O(N__12734),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    CascadeMux I__1730 (
            .O(N__12725),
            .I(\uart_pc.un1_state_4_0_cascade_ ));
    InMux I__1729 (
            .O(N__12722),
            .I(N__12719));
    LocalMux I__1728 (
            .O(N__12719),
            .I(\uart_pc.CO0 ));
    InMux I__1727 (
            .O(N__12716),
            .I(N__12712));
    InMux I__1726 (
            .O(N__12715),
            .I(N__12709));
    LocalMux I__1725 (
            .O(N__12712),
            .I(\uart_pc.un1_state_7_0 ));
    LocalMux I__1724 (
            .O(N__12709),
            .I(\uart_pc.un1_state_7_0 ));
    CascadeMux I__1723 (
            .O(N__12704),
            .I(N__12696));
    CascadeMux I__1722 (
            .O(N__12703),
            .I(N__12693));
    InMux I__1721 (
            .O(N__12702),
            .I(N__12685));
    InMux I__1720 (
            .O(N__12701),
            .I(N__12685));
    InMux I__1719 (
            .O(N__12700),
            .I(N__12682));
    InMux I__1718 (
            .O(N__12699),
            .I(N__12671));
    InMux I__1717 (
            .O(N__12696),
            .I(N__12671));
    InMux I__1716 (
            .O(N__12693),
            .I(N__12671));
    InMux I__1715 (
            .O(N__12692),
            .I(N__12671));
    InMux I__1714 (
            .O(N__12691),
            .I(N__12671));
    InMux I__1713 (
            .O(N__12690),
            .I(N__12667));
    LocalMux I__1712 (
            .O(N__12685),
            .I(N__12664));
    LocalMux I__1711 (
            .O(N__12682),
            .I(N__12659));
    LocalMux I__1710 (
            .O(N__12671),
            .I(N__12659));
    InMux I__1709 (
            .O(N__12670),
            .I(N__12656));
    LocalMux I__1708 (
            .O(N__12667),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv12 I__1707 (
            .O(N__12664),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    Odrv4 I__1706 (
            .O(N__12659),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__1705 (
            .O(N__12656),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    CascadeMux I__1704 (
            .O(N__12647),
            .I(N__12643));
    CascadeMux I__1703 (
            .O(N__12646),
            .I(N__12640));
    InMux I__1702 (
            .O(N__12643),
            .I(N__12635));
    InMux I__1701 (
            .O(N__12640),
            .I(N__12635));
    LocalMux I__1700 (
            .O(N__12635),
            .I(N__12631));
    InMux I__1699 (
            .O(N__12634),
            .I(N__12628));
    Odrv4 I__1698 (
            .O(N__12631),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__1697 (
            .O(N__12628),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__1696 (
            .O(N__12623),
            .I(N__12610));
    InMux I__1695 (
            .O(N__12622),
            .I(N__12610));
    InMux I__1694 (
            .O(N__12621),
            .I(N__12599));
    InMux I__1693 (
            .O(N__12620),
            .I(N__12599));
    InMux I__1692 (
            .O(N__12619),
            .I(N__12599));
    InMux I__1691 (
            .O(N__12618),
            .I(N__12599));
    InMux I__1690 (
            .O(N__12617),
            .I(N__12599));
    InMux I__1689 (
            .O(N__12616),
            .I(N__12592));
    InMux I__1688 (
            .O(N__12615),
            .I(N__12592));
    LocalMux I__1687 (
            .O(N__12610),
            .I(N__12587));
    LocalMux I__1686 (
            .O(N__12599),
            .I(N__12587));
    InMux I__1685 (
            .O(N__12598),
            .I(N__12582));
    InMux I__1684 (
            .O(N__12597),
            .I(N__12582));
    LocalMux I__1683 (
            .O(N__12592),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv12 I__1682 (
            .O(N__12587),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__1681 (
            .O(N__12582),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    SRMux I__1680 (
            .O(N__12575),
            .I(N__12571));
    SRMux I__1679 (
            .O(N__12574),
            .I(N__12568));
    LocalMux I__1678 (
            .O(N__12571),
            .I(N__12565));
    LocalMux I__1677 (
            .O(N__12568),
            .I(N__12562));
    Odrv4 I__1676 (
            .O(N__12565),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv4 I__1675 (
            .O(N__12562),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__1674 (
            .O(N__12557),
            .I(N__12554));
    LocalMux I__1673 (
            .O(N__12554),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    InMux I__1672 (
            .O(N__12551),
            .I(N__12548));
    LocalMux I__1671 (
            .O(N__12548),
            .I(\uart_pc.data_Auxce_0_3 ));
    InMux I__1670 (
            .O(N__12545),
            .I(N__12542));
    LocalMux I__1669 (
            .O(N__12542),
            .I(\uart_pc.data_Auxce_0_5 ));
    InMux I__1668 (
            .O(N__12539),
            .I(N__12536));
    LocalMux I__1667 (
            .O(N__12536),
            .I(N__12533));
    Odrv4 I__1666 (
            .O(N__12533),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__1665 (
            .O(N__12530),
            .I(N__12524));
    InMux I__1664 (
            .O(N__12529),
            .I(N__12519));
    InMux I__1663 (
            .O(N__12528),
            .I(N__12514));
    InMux I__1662 (
            .O(N__12527),
            .I(N__12514));
    LocalMux I__1661 (
            .O(N__12524),
            .I(N__12511));
    InMux I__1660 (
            .O(N__12523),
            .I(N__12508));
    InMux I__1659 (
            .O(N__12522),
            .I(N__12505));
    LocalMux I__1658 (
            .O(N__12519),
            .I(N__12500));
    LocalMux I__1657 (
            .O(N__12514),
            .I(N__12500));
    Odrv4 I__1656 (
            .O(N__12511),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__1655 (
            .O(N__12508),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__1654 (
            .O(N__12505),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__1653 (
            .O(N__12500),
            .I(\uart_drone.stateZ0Z_4 ));
    CascadeMux I__1652 (
            .O(N__12491),
            .I(N__12488));
    InMux I__1651 (
            .O(N__12488),
            .I(N__12485));
    LocalMux I__1650 (
            .O(N__12485),
            .I(N__12481));
    InMux I__1649 (
            .O(N__12484),
            .I(N__12478));
    Odrv4 I__1648 (
            .O(N__12481),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__1647 (
            .O(N__12478),
            .I(\uart_drone.stateZ0Z_0 ));
    CascadeMux I__1646 (
            .O(N__12473),
            .I(N__12470));
    InMux I__1645 (
            .O(N__12470),
            .I(N__12464));
    InMux I__1644 (
            .O(N__12469),
            .I(N__12461));
    InMux I__1643 (
            .O(N__12468),
            .I(N__12456));
    InMux I__1642 (
            .O(N__12467),
            .I(N__12456));
    LocalMux I__1641 (
            .O(N__12464),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__1640 (
            .O(N__12461),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__1639 (
            .O(N__12456),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__1638 (
            .O(N__12449),
            .I(N__12436));
    InMux I__1637 (
            .O(N__12448),
            .I(N__12436));
    InMux I__1636 (
            .O(N__12447),
            .I(N__12431));
    InMux I__1635 (
            .O(N__12446),
            .I(N__12431));
    InMux I__1634 (
            .O(N__12445),
            .I(N__12424));
    InMux I__1633 (
            .O(N__12444),
            .I(N__12424));
    InMux I__1632 (
            .O(N__12443),
            .I(N__12424));
    InMux I__1631 (
            .O(N__12442),
            .I(N__12417));
    InMux I__1630 (
            .O(N__12441),
            .I(N__12417));
    LocalMux I__1629 (
            .O(N__12436),
            .I(N__12414));
    LocalMux I__1628 (
            .O(N__12431),
            .I(N__12411));
    LocalMux I__1627 (
            .O(N__12424),
            .I(N__12408));
    InMux I__1626 (
            .O(N__12423),
            .I(N__12403));
    InMux I__1625 (
            .O(N__12422),
            .I(N__12403));
    LocalMux I__1624 (
            .O(N__12417),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__1623 (
            .O(N__12414),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv12 I__1622 (
            .O(N__12411),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__1621 (
            .O(N__12408),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__1620 (
            .O(N__12403),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__1619 (
            .O(N__12392),
            .I(N__12389));
    LocalMux I__1618 (
            .O(N__12389),
            .I(\uart_drone.CO0 ));
    InMux I__1617 (
            .O(N__12386),
            .I(N__12382));
    InMux I__1616 (
            .O(N__12385),
            .I(N__12379));
    LocalMux I__1615 (
            .O(N__12382),
            .I(\uart_drone.un1_state_7_0 ));
    LocalMux I__1614 (
            .O(N__12379),
            .I(\uart_drone.un1_state_7_0 ));
    CascadeMux I__1613 (
            .O(N__12374),
            .I(N__12367));
    InMux I__1612 (
            .O(N__12373),
            .I(N__12358));
    InMux I__1611 (
            .O(N__12372),
            .I(N__12358));
    InMux I__1610 (
            .O(N__12371),
            .I(N__12353));
    InMux I__1609 (
            .O(N__12370),
            .I(N__12353));
    InMux I__1608 (
            .O(N__12367),
            .I(N__12346));
    InMux I__1607 (
            .O(N__12366),
            .I(N__12346));
    InMux I__1606 (
            .O(N__12365),
            .I(N__12346));
    InMux I__1605 (
            .O(N__12364),
            .I(N__12342));
    InMux I__1604 (
            .O(N__12363),
            .I(N__12339));
    LocalMux I__1603 (
            .O(N__12358),
            .I(N__12336));
    LocalMux I__1602 (
            .O(N__12353),
            .I(N__12333));
    LocalMux I__1601 (
            .O(N__12346),
            .I(N__12330));
    InMux I__1600 (
            .O(N__12345),
            .I(N__12327));
    LocalMux I__1599 (
            .O(N__12342),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__1598 (
            .O(N__12339),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__1597 (
            .O(N__12336),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__1596 (
            .O(N__12333),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__1595 (
            .O(N__12330),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__1594 (
            .O(N__12327),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__1593 (
            .O(N__12314),
            .I(N__12304));
    InMux I__1592 (
            .O(N__12313),
            .I(N__12304));
    InMux I__1591 (
            .O(N__12312),
            .I(N__12297));
    InMux I__1590 (
            .O(N__12311),
            .I(N__12297));
    InMux I__1589 (
            .O(N__12310),
            .I(N__12297));
    CascadeMux I__1588 (
            .O(N__12309),
            .I(N__12292));
    LocalMux I__1587 (
            .O(N__12304),
            .I(N__12287));
    LocalMux I__1586 (
            .O(N__12297),
            .I(N__12287));
    InMux I__1585 (
            .O(N__12296),
            .I(N__12282));
    InMux I__1584 (
            .O(N__12295),
            .I(N__12282));
    InMux I__1583 (
            .O(N__12292),
            .I(N__12278));
    Sp12to4 I__1582 (
            .O(N__12287),
            .I(N__12273));
    LocalMux I__1581 (
            .O(N__12282),
            .I(N__12273));
    InMux I__1580 (
            .O(N__12281),
            .I(N__12270));
    LocalMux I__1579 (
            .O(N__12278),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv12 I__1578 (
            .O(N__12273),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__1577 (
            .O(N__12270),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__1576 (
            .O(N__12263),
            .I(N__12260));
    LocalMux I__1575 (
            .O(N__12260),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__1574 (
            .O(N__12257),
            .I(N__12254));
    LocalMux I__1573 (
            .O(N__12254),
            .I(\uart_pc.data_Auxce_0_6 ));
    InMux I__1572 (
            .O(N__12251),
            .I(N__12248));
    LocalMux I__1571 (
            .O(N__12248),
            .I(\uart_pc.data_Auxce_0_1 ));
    CascadeMux I__1570 (
            .O(N__12245),
            .I(N__12242));
    InMux I__1569 (
            .O(N__12242),
            .I(N__12233));
    InMux I__1568 (
            .O(N__12241),
            .I(N__12233));
    InMux I__1567 (
            .O(N__12240),
            .I(N__12230));
    InMux I__1566 (
            .O(N__12239),
            .I(N__12225));
    InMux I__1565 (
            .O(N__12238),
            .I(N__12225));
    LocalMux I__1564 (
            .O(N__12233),
            .I(\uart_drone.N_143 ));
    LocalMux I__1563 (
            .O(N__12230),
            .I(\uart_drone.N_143 ));
    LocalMux I__1562 (
            .O(N__12225),
            .I(\uart_drone.N_143 ));
    InMux I__1561 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__1560 (
            .O(N__12215),
            .I(\uart_drone.N_144_1 ));
    CascadeMux I__1559 (
            .O(N__12212),
            .I(\uart_drone.N_144_1_cascade_ ));
    CascadeMux I__1558 (
            .O(N__12209),
            .I(N__12204));
    CascadeMux I__1557 (
            .O(N__12208),
            .I(N__12201));
    CascadeMux I__1556 (
            .O(N__12207),
            .I(N__12197));
    InMux I__1555 (
            .O(N__12204),
            .I(N__12192));
    InMux I__1554 (
            .O(N__12201),
            .I(N__12192));
    InMux I__1553 (
            .O(N__12200),
            .I(N__12187));
    InMux I__1552 (
            .O(N__12197),
            .I(N__12187));
    LocalMux I__1551 (
            .O(N__12192),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__1550 (
            .O(N__12187),
            .I(\uart_drone.stateZ0Z_2 ));
    InMux I__1549 (
            .O(N__12182),
            .I(N__12179));
    LocalMux I__1548 (
            .O(N__12179),
            .I(\uart_drone.N_145 ));
    InMux I__1547 (
            .O(N__12176),
            .I(N__12166));
    InMux I__1546 (
            .O(N__12175),
            .I(N__12163));
    InMux I__1545 (
            .O(N__12174),
            .I(N__12160));
    InMux I__1544 (
            .O(N__12173),
            .I(N__12153));
    InMux I__1543 (
            .O(N__12172),
            .I(N__12153));
    InMux I__1542 (
            .O(N__12171),
            .I(N__12153));
    InMux I__1541 (
            .O(N__12170),
            .I(N__12148));
    InMux I__1540 (
            .O(N__12169),
            .I(N__12148));
    LocalMux I__1539 (
            .O(N__12166),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__1538 (
            .O(N__12163),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__1537 (
            .O(N__12160),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__1536 (
            .O(N__12153),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__1535 (
            .O(N__12148),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    CascadeMux I__1534 (
            .O(N__12137),
            .I(N__12130));
    InMux I__1533 (
            .O(N__12136),
            .I(N__12126));
    InMux I__1532 (
            .O(N__12135),
            .I(N__12123));
    CascadeMux I__1531 (
            .O(N__12134),
            .I(N__12119));
    CascadeMux I__1530 (
            .O(N__12133),
            .I(N__12115));
    InMux I__1529 (
            .O(N__12130),
            .I(N__12112));
    InMux I__1528 (
            .O(N__12129),
            .I(N__12109));
    LocalMux I__1527 (
            .O(N__12126),
            .I(N__12104));
    LocalMux I__1526 (
            .O(N__12123),
            .I(N__12104));
    InMux I__1525 (
            .O(N__12122),
            .I(N__12101));
    InMux I__1524 (
            .O(N__12119),
            .I(N__12094));
    InMux I__1523 (
            .O(N__12118),
            .I(N__12094));
    InMux I__1522 (
            .O(N__12115),
            .I(N__12094));
    LocalMux I__1521 (
            .O(N__12112),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__1520 (
            .O(N__12109),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__1519 (
            .O(N__12104),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__1518 (
            .O(N__12101),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__1517 (
            .O(N__12094),
            .I(\uart_drone.stateZ0Z_3 ));
    InMux I__1516 (
            .O(N__12083),
            .I(N__12079));
    InMux I__1515 (
            .O(N__12082),
            .I(N__12074));
    LocalMux I__1514 (
            .O(N__12079),
            .I(N__12071));
    InMux I__1513 (
            .O(N__12078),
            .I(N__12068));
    InMux I__1512 (
            .O(N__12077),
            .I(N__12065));
    LocalMux I__1511 (
            .O(N__12074),
            .I(\uart_drone.N_152 ));
    Odrv12 I__1510 (
            .O(N__12071),
            .I(\uart_drone.N_152 ));
    LocalMux I__1509 (
            .O(N__12068),
            .I(\uart_drone.N_152 ));
    LocalMux I__1508 (
            .O(N__12065),
            .I(\uart_drone.N_152 ));
    InMux I__1507 (
            .O(N__12056),
            .I(N__12052));
    IoInMux I__1506 (
            .O(N__12055),
            .I(N__12047));
    LocalMux I__1505 (
            .O(N__12052),
            .I(N__12044));
    InMux I__1504 (
            .O(N__12051),
            .I(N__12036));
    InMux I__1503 (
            .O(N__12050),
            .I(N__12033));
    LocalMux I__1502 (
            .O(N__12047),
            .I(N__12030));
    Span4Mux_v I__1501 (
            .O(N__12044),
            .I(N__12027));
    InMux I__1500 (
            .O(N__12043),
            .I(N__12018));
    InMux I__1499 (
            .O(N__12042),
            .I(N__12018));
    InMux I__1498 (
            .O(N__12041),
            .I(N__12018));
    InMux I__1497 (
            .O(N__12040),
            .I(N__12018));
    InMux I__1496 (
            .O(N__12039),
            .I(N__12010));
    LocalMux I__1495 (
            .O(N__12036),
            .I(N__12007));
    LocalMux I__1494 (
            .O(N__12033),
            .I(N__12004));
    IoSpan4Mux I__1493 (
            .O(N__12030),
            .I(N__12001));
    Sp12to4 I__1492 (
            .O(N__12027),
            .I(N__11998));
    LocalMux I__1491 (
            .O(N__12018),
            .I(N__11995));
    InMux I__1490 (
            .O(N__12017),
            .I(N__11990));
    InMux I__1489 (
            .O(N__12016),
            .I(N__11990));
    InMux I__1488 (
            .O(N__12015),
            .I(N__11987));
    InMux I__1487 (
            .O(N__12014),
            .I(N__11984));
    InMux I__1486 (
            .O(N__12013),
            .I(N__11981));
    LocalMux I__1485 (
            .O(N__12010),
            .I(N__11974));
    Span4Mux_v I__1484 (
            .O(N__12007),
            .I(N__11974));
    Span4Mux_h I__1483 (
            .O(N__12004),
            .I(N__11974));
    Span4Mux_s1_v I__1482 (
            .O(N__12001),
            .I(N__11971));
    Span12Mux_h I__1481 (
            .O(N__11998),
            .I(N__11958));
    Sp12to4 I__1480 (
            .O(N__11995),
            .I(N__11958));
    LocalMux I__1479 (
            .O(N__11990),
            .I(N__11958));
    LocalMux I__1478 (
            .O(N__11987),
            .I(N__11958));
    LocalMux I__1477 (
            .O(N__11984),
            .I(N__11958));
    LocalMux I__1476 (
            .O(N__11981),
            .I(N__11958));
    Span4Mux_v I__1475 (
            .O(N__11974),
            .I(N__11955));
    Span4Mux_h I__1474 (
            .O(N__11971),
            .I(N__11952));
    Span12Mux_v I__1473 (
            .O(N__11958),
            .I(N__11947));
    Sp12to4 I__1472 (
            .O(N__11955),
            .I(N__11947));
    Odrv4 I__1471 (
            .O(N__11952),
            .I(uart_input_debug_c));
    Odrv12 I__1470 (
            .O(N__11947),
            .I(uart_input_debug_c));
    InMux I__1469 (
            .O(N__11942),
            .I(N__11934));
    InMux I__1468 (
            .O(N__11941),
            .I(N__11929));
    InMux I__1467 (
            .O(N__11940),
            .I(N__11929));
    CascadeMux I__1466 (
            .O(N__11939),
            .I(N__11923));
    InMux I__1465 (
            .O(N__11938),
            .I(N__11920));
    InMux I__1464 (
            .O(N__11937),
            .I(N__11917));
    LocalMux I__1463 (
            .O(N__11934),
            .I(N__11912));
    LocalMux I__1462 (
            .O(N__11929),
            .I(N__11912));
    InMux I__1461 (
            .O(N__11928),
            .I(N__11905));
    InMux I__1460 (
            .O(N__11927),
            .I(N__11905));
    InMux I__1459 (
            .O(N__11926),
            .I(N__11905));
    InMux I__1458 (
            .O(N__11923),
            .I(N__11902));
    LocalMux I__1457 (
            .O(N__11920),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__1456 (
            .O(N__11917),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__1455 (
            .O(N__11912),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__1454 (
            .O(N__11905),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__1453 (
            .O(N__11902),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__1452 (
            .O(N__11891),
            .I(N__11888));
    LocalMux I__1451 (
            .O(N__11888),
            .I(N__11884));
    InMux I__1450 (
            .O(N__11887),
            .I(N__11881));
    Odrv4 I__1449 (
            .O(N__11884),
            .I(\uart_drone.N_126_li ));
    LocalMux I__1448 (
            .O(N__11881),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__1447 (
            .O(N__11876),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__1446 (
            .O(N__11873),
            .I(N__11870));
    LocalMux I__1445 (
            .O(N__11870),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__1444 (
            .O(N__11867),
            .I(N__11861));
    InMux I__1443 (
            .O(N__11866),
            .I(N__11861));
    LocalMux I__1442 (
            .O(N__11861),
            .I(N__11852));
    InMux I__1441 (
            .O(N__11860),
            .I(N__11847));
    InMux I__1440 (
            .O(N__11859),
            .I(N__11847));
    InMux I__1439 (
            .O(N__11858),
            .I(N__11838));
    InMux I__1438 (
            .O(N__11857),
            .I(N__11838));
    InMux I__1437 (
            .O(N__11856),
            .I(N__11838));
    InMux I__1436 (
            .O(N__11855),
            .I(N__11838));
    Odrv4 I__1435 (
            .O(N__11852),
            .I(\uart_drone.un1_state_2_0 ));
    LocalMux I__1434 (
            .O(N__11847),
            .I(\uart_drone.un1_state_2_0 ));
    LocalMux I__1433 (
            .O(N__11838),
            .I(\uart_drone.un1_state_2_0 ));
    CascadeMux I__1432 (
            .O(N__11831),
            .I(N__11827));
    InMux I__1431 (
            .O(N__11830),
            .I(N__11824));
    InMux I__1430 (
            .O(N__11827),
            .I(N__11821));
    LocalMux I__1429 (
            .O(N__11824),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__1428 (
            .O(N__11821),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    InMux I__1427 (
            .O(N__11816),
            .I(N__11813));
    LocalMux I__1426 (
            .O(N__11813),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__1425 (
            .O(N__11810),
            .I(N__11807));
    LocalMux I__1424 (
            .O(N__11807),
            .I(N__11804));
    Odrv4 I__1423 (
            .O(N__11804),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    SRMux I__1422 (
            .O(N__11801),
            .I(N__11797));
    SRMux I__1421 (
            .O(N__11800),
            .I(N__11794));
    LocalMux I__1420 (
            .O(N__11797),
            .I(N__11790));
    LocalMux I__1419 (
            .O(N__11794),
            .I(N__11787));
    SRMux I__1418 (
            .O(N__11793),
            .I(N__11784));
    Span4Mux_h I__1417 (
            .O(N__11790),
            .I(N__11777));
    Span4Mux_v I__1416 (
            .O(N__11787),
            .I(N__11777));
    LocalMux I__1415 (
            .O(N__11784),
            .I(N__11777));
    Span4Mux_h I__1414 (
            .O(N__11777),
            .I(N__11774));
    Odrv4 I__1413 (
            .O(N__11774),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__1412 (
            .O(N__11771),
            .I(N__11768));
    LocalMux I__1411 (
            .O(N__11768),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    CascadeMux I__1410 (
            .O(N__11765),
            .I(\uart_drone.N_143_cascade_ ));
    CascadeMux I__1409 (
            .O(N__11762),
            .I(N__11756));
    InMux I__1408 (
            .O(N__11761),
            .I(N__11751));
    InMux I__1407 (
            .O(N__11760),
            .I(N__11751));
    InMux I__1406 (
            .O(N__11759),
            .I(N__11746));
    InMux I__1405 (
            .O(N__11756),
            .I(N__11746));
    LocalMux I__1404 (
            .O(N__11751),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__1403 (
            .O(N__11746),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__1402 (
            .O(N__11741),
            .I(N__11736));
    InMux I__1401 (
            .O(N__11740),
            .I(N__11731));
    InMux I__1400 (
            .O(N__11739),
            .I(N__11726));
    InMux I__1399 (
            .O(N__11736),
            .I(N__11726));
    InMux I__1398 (
            .O(N__11735),
            .I(N__11721));
    InMux I__1397 (
            .O(N__11734),
            .I(N__11721));
    LocalMux I__1396 (
            .O(N__11731),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__1395 (
            .O(N__11726),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__1394 (
            .O(N__11721),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__1393 (
            .O(N__11714),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    InMux I__1392 (
            .O(N__11711),
            .I(N__11707));
    InMux I__1391 (
            .O(N__11710),
            .I(N__11704));
    LocalMux I__1390 (
            .O(N__11707),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__1389 (
            .O(N__11704),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    InMux I__1388 (
            .O(N__11699),
            .I(N__11696));
    LocalMux I__1387 (
            .O(N__11696),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    CascadeMux I__1386 (
            .O(N__11693),
            .I(N__11689));
    CascadeMux I__1385 (
            .O(N__11692),
            .I(N__11685));
    InMux I__1384 (
            .O(N__11689),
            .I(N__11682));
    InMux I__1383 (
            .O(N__11688),
            .I(N__11679));
    InMux I__1382 (
            .O(N__11685),
            .I(N__11676));
    LocalMux I__1381 (
            .O(N__11682),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__1380 (
            .O(N__11679),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__1379 (
            .O(N__11676),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__1378 (
            .O(N__11669),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    InMux I__1377 (
            .O(N__11666),
            .I(N__11663));
    LocalMux I__1376 (
            .O(N__11663),
            .I(\uart_pc.state_srsts_0_0_0 ));
    InMux I__1375 (
            .O(N__11660),
            .I(N__11657));
    LocalMux I__1374 (
            .O(N__11657),
            .I(N__11653));
    InMux I__1373 (
            .O(N__11656),
            .I(N__11650));
    Odrv4 I__1372 (
            .O(N__11653),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__1371 (
            .O(N__11650),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__1370 (
            .O(N__11645),
            .I(N__11641));
    InMux I__1369 (
            .O(N__11644),
            .I(N__11638));
    InMux I__1368 (
            .O(N__11641),
            .I(N__11635));
    LocalMux I__1367 (
            .O(N__11638),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__1366 (
            .O(N__11635),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    InMux I__1365 (
            .O(N__11630),
            .I(N__11627));
    LocalMux I__1364 (
            .O(N__11627),
            .I(N__11623));
    CascadeMux I__1363 (
            .O(N__11626),
            .I(N__11620));
    Span12Mux_v I__1362 (
            .O(N__11623),
            .I(N__11617));
    InMux I__1361 (
            .O(N__11620),
            .I(N__11614));
    Odrv12 I__1360 (
            .O(N__11617),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__1359 (
            .O(N__11614),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    CascadeMux I__1358 (
            .O(N__11609),
            .I(N__11605));
    InMux I__1357 (
            .O(N__11608),
            .I(N__11602));
    InMux I__1356 (
            .O(N__11605),
            .I(N__11599));
    LocalMux I__1355 (
            .O(N__11602),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__1354 (
            .O(N__11599),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    InMux I__1353 (
            .O(N__11594),
            .I(N__11591));
    LocalMux I__1352 (
            .O(N__11591),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__1351 (
            .O(N__11588),
            .I(N__11585));
    LocalMux I__1350 (
            .O(N__11585),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__1349 (
            .O(N__11582),
            .I(N__11577));
    InMux I__1348 (
            .O(N__11581),
            .I(N__11572));
    InMux I__1347 (
            .O(N__11580),
            .I(N__11572));
    LocalMux I__1346 (
            .O(N__11577),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__1345 (
            .O(N__11572),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    CascadeMux I__1344 (
            .O(N__11567),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__1343 (
            .O(N__11564),
            .I(N__11559));
    InMux I__1342 (
            .O(N__11563),
            .I(N__11556));
    InMux I__1341 (
            .O(N__11562),
            .I(N__11553));
    LocalMux I__1340 (
            .O(N__11559),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__1339 (
            .O(N__11556),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__1338 (
            .O(N__11553),
            .I(\uart_drone.stateZ0Z_1 ));
    InMux I__1337 (
            .O(N__11546),
            .I(N__11540));
    InMux I__1336 (
            .O(N__11545),
            .I(N__11537));
    InMux I__1335 (
            .O(N__11544),
            .I(N__11532));
    InMux I__1334 (
            .O(N__11543),
            .I(N__11532));
    LocalMux I__1333 (
            .O(N__11540),
            .I(N__11529));
    LocalMux I__1332 (
            .O(N__11537),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__1331 (
            .O(N__11532),
            .I(\reset_module_System.countZ0Z_0 ));
    Odrv4 I__1330 (
            .O(N__11529),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__1329 (
            .O(N__11522),
            .I(N__11517));
    InMux I__1328 (
            .O(N__11521),
            .I(N__11512));
    InMux I__1327 (
            .O(N__11520),
            .I(N__11512));
    LocalMux I__1326 (
            .O(N__11517),
            .I(\reset_module_System.reset6_15 ));
    LocalMux I__1325 (
            .O(N__11512),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__1324 (
            .O(N__11507),
            .I(N__11503));
    InMux I__1323 (
            .O(N__11506),
            .I(N__11496));
    InMux I__1322 (
            .O(N__11503),
            .I(N__11496));
    InMux I__1321 (
            .O(N__11502),
            .I(N__11491));
    InMux I__1320 (
            .O(N__11501),
            .I(N__11491));
    LocalMux I__1319 (
            .O(N__11496),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__1318 (
            .O(N__11491),
            .I(\reset_module_System.reset6_14 ));
    CascadeMux I__1317 (
            .O(N__11486),
            .I(\reset_module_System.count_1_1_cascade_ ));
    InMux I__1316 (
            .O(N__11483),
            .I(N__11475));
    InMux I__1315 (
            .O(N__11482),
            .I(N__11475));
    InMux I__1314 (
            .O(N__11481),
            .I(N__11470));
    InMux I__1313 (
            .O(N__11480),
            .I(N__11470));
    LocalMux I__1312 (
            .O(N__11475),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__1311 (
            .O(N__11470),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__1310 (
            .O(N__11465),
            .I(N__11462));
    InMux I__1309 (
            .O(N__11462),
            .I(N__11458));
    InMux I__1308 (
            .O(N__11461),
            .I(N__11454));
    LocalMux I__1307 (
            .O(N__11458),
            .I(N__11451));
    InMux I__1306 (
            .O(N__11457),
            .I(N__11448));
    LocalMux I__1305 (
            .O(N__11454),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__1304 (
            .O(N__11451),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__1303 (
            .O(N__11448),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__1302 (
            .O(N__11441),
            .I(N__11436));
    InMux I__1301 (
            .O(N__11440),
            .I(N__11431));
    InMux I__1300 (
            .O(N__11439),
            .I(N__11431));
    LocalMux I__1299 (
            .O(N__11436),
            .I(N__11428));
    LocalMux I__1298 (
            .O(N__11431),
            .I(N__11425));
    Odrv12 I__1297 (
            .O(N__11428),
            .I(\uart_drone.state_1_sqmuxa ));
    Odrv4 I__1296 (
            .O(N__11425),
            .I(\uart_drone.state_1_sqmuxa ));
    InMux I__1295 (
            .O(N__11420),
            .I(N__11417));
    LocalMux I__1294 (
            .O(N__11417),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__1293 (
            .O(N__11414),
            .I(N__11411));
    LocalMux I__1292 (
            .O(N__11411),
            .I(\uart_drone.data_Auxce_0_3 ));
    CascadeMux I__1291 (
            .O(N__11408),
            .I(\uart_drone.N_126_li_cascade_ ));
    InMux I__1290 (
            .O(N__11405),
            .I(N__11402));
    LocalMux I__1289 (
            .O(N__11402),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    InMux I__1288 (
            .O(N__11399),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__1287 (
            .O(N__11396),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__1286 (
            .O(N__11393),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__1285 (
            .O(N__11390),
            .I(N__11383));
    InMux I__1284 (
            .O(N__11389),
            .I(N__11383));
    InMux I__1283 (
            .O(N__11388),
            .I(N__11380));
    LocalMux I__1282 (
            .O(N__11383),
            .I(N__11376));
    LocalMux I__1281 (
            .O(N__11380),
            .I(N__11373));
    InMux I__1280 (
            .O(N__11379),
            .I(N__11370));
    Span4Mux_s3_h I__1279 (
            .O(N__11376),
            .I(N__11367));
    Span4Mux_s3_h I__1278 (
            .O(N__11373),
            .I(N__11364));
    LocalMux I__1277 (
            .O(N__11370),
            .I(uart_drone_data_6));
    Odrv4 I__1276 (
            .O(N__11367),
            .I(uart_drone_data_6));
    Odrv4 I__1275 (
            .O(N__11364),
            .I(uart_drone_data_6));
    InMux I__1274 (
            .O(N__11357),
            .I(N__11354));
    LocalMux I__1273 (
            .O(N__11354),
            .I(uart_drone_data_7));
    CEMux I__1272 (
            .O(N__11351),
            .I(N__11348));
    LocalMux I__1271 (
            .O(N__11348),
            .I(N__11344));
    CEMux I__1270 (
            .O(N__11347),
            .I(N__11341));
    Span4Mux_v I__1269 (
            .O(N__11344),
            .I(N__11338));
    LocalMux I__1268 (
            .O(N__11341),
            .I(N__11335));
    Odrv4 I__1267 (
            .O(N__11338),
            .I(\uart_drone.state_1_sqmuxa_0 ));
    Odrv4 I__1266 (
            .O(N__11335),
            .I(\uart_drone.state_1_sqmuxa_0 ));
    SRMux I__1265 (
            .O(N__11330),
            .I(N__11327));
    LocalMux I__1264 (
            .O(N__11327),
            .I(N__11323));
    SRMux I__1263 (
            .O(N__11326),
            .I(N__11320));
    Span4Mux_v I__1262 (
            .O(N__11323),
            .I(N__11315));
    LocalMux I__1261 (
            .O(N__11320),
            .I(N__11315));
    Odrv4 I__1260 (
            .O(N__11315),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    CascadeMux I__1259 (
            .O(N__11312),
            .I(N__11308));
    InMux I__1258 (
            .O(N__11311),
            .I(N__11305));
    InMux I__1257 (
            .O(N__11308),
            .I(N__11302));
    LocalMux I__1256 (
            .O(N__11305),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__1255 (
            .O(N__11302),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    CascadeMux I__1254 (
            .O(N__11297),
            .I(N__11293));
    InMux I__1253 (
            .O(N__11296),
            .I(N__11290));
    InMux I__1252 (
            .O(N__11293),
            .I(N__11287));
    LocalMux I__1251 (
            .O(N__11290),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__1250 (
            .O(N__11287),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__1249 (
            .O(N__11282),
            .I(N__11278));
    InMux I__1248 (
            .O(N__11281),
            .I(N__11275));
    InMux I__1247 (
            .O(N__11278),
            .I(N__11272));
    LocalMux I__1246 (
            .O(N__11275),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__1245 (
            .O(N__11272),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    CascadeMux I__1244 (
            .O(N__11267),
            .I(\uart_drone.data_Auxce_0_0_4_cascade_ ));
    InMux I__1243 (
            .O(N__11264),
            .I(N__11261));
    LocalMux I__1242 (
            .O(N__11261),
            .I(N__11258));
    Span4Mux_v I__1241 (
            .O(N__11258),
            .I(N__11254));
    InMux I__1240 (
            .O(N__11257),
            .I(N__11251));
    Odrv4 I__1239 (
            .O(N__11254),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__1238 (
            .O(N__11251),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    InMux I__1237 (
            .O(N__11246),
            .I(N__11243));
    LocalMux I__1236 (
            .O(N__11243),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__1235 (
            .O(N__11240),
            .I(N__11237));
    LocalMux I__1234 (
            .O(N__11237),
            .I(N__11234));
    Span4Mux_v I__1233 (
            .O(N__11234),
            .I(N__11229));
    InMux I__1232 (
            .O(N__11233),
            .I(N__11226));
    InMux I__1231 (
            .O(N__11232),
            .I(N__11223));
    Odrv4 I__1230 (
            .O(N__11229),
            .I(\frame_dron_decoder_1.stateZ0Z_6 ));
    LocalMux I__1229 (
            .O(N__11226),
            .I(\frame_dron_decoder_1.stateZ0Z_6 ));
    LocalMux I__1228 (
            .O(N__11223),
            .I(\frame_dron_decoder_1.stateZ0Z_6 ));
    IoInMux I__1227 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1226 (
            .O(N__11213),
            .I(N__11210));
    Span12Mux_s1_v I__1225 (
            .O(N__11210),
            .I(N__11207));
    Span12Mux_v I__1224 (
            .O(N__11207),
            .I(N__11203));
    InMux I__1223 (
            .O(N__11206),
            .I(N__11200));
    Odrv12 I__1222 (
            .O(N__11203),
            .I(drone_frame_decoder_data_rdy_debug_c));
    LocalMux I__1221 (
            .O(N__11200),
            .I(drone_frame_decoder_data_rdy_debug_c));
    InMux I__1220 (
            .O(N__11195),
            .I(N__11192));
    LocalMux I__1219 (
            .O(N__11192),
            .I(N__11189));
    Odrv4 I__1218 (
            .O(N__11189),
            .I(uart_drone_data_2));
    CascadeMux I__1217 (
            .O(N__11186),
            .I(\frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ));
    InMux I__1216 (
            .O(N__11183),
            .I(N__11179));
    InMux I__1215 (
            .O(N__11182),
            .I(N__11175));
    LocalMux I__1214 (
            .O(N__11179),
            .I(N__11172));
    InMux I__1213 (
            .O(N__11178),
            .I(N__11169));
    LocalMux I__1212 (
            .O(N__11175),
            .I(N__11164));
    Span4Mux_s3_h I__1211 (
            .O(N__11172),
            .I(N__11164));
    LocalMux I__1210 (
            .O(N__11169),
            .I(N__11161));
    Odrv4 I__1209 (
            .O(N__11164),
            .I(\frame_dron_decoder_1.N_255 ));
    Odrv4 I__1208 (
            .O(N__11161),
            .I(\frame_dron_decoder_1.N_255 ));
    IoInMux I__1207 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__1206 (
            .O(N__11153),
            .I(N__11150));
    Span4Mux_s1_v I__1205 (
            .O(N__11150),
            .I(N__11145));
    CascadeMux I__1204 (
            .O(N__11149),
            .I(N__11142));
    CascadeMux I__1203 (
            .O(N__11148),
            .I(N__11138));
    Sp12to4 I__1202 (
            .O(N__11145),
            .I(N__11131));
    InMux I__1201 (
            .O(N__11142),
            .I(N__11122));
    InMux I__1200 (
            .O(N__11141),
            .I(N__11122));
    InMux I__1199 (
            .O(N__11138),
            .I(N__11122));
    InMux I__1198 (
            .O(N__11137),
            .I(N__11122));
    InMux I__1197 (
            .O(N__11136),
            .I(N__11118));
    InMux I__1196 (
            .O(N__11135),
            .I(N__11115));
    InMux I__1195 (
            .O(N__11134),
            .I(N__11112));
    Span12Mux_h I__1194 (
            .O(N__11131),
            .I(N__11109));
    LocalMux I__1193 (
            .O(N__11122),
            .I(N__11106));
    InMux I__1192 (
            .O(N__11121),
            .I(N__11103));
    LocalMux I__1191 (
            .O(N__11118),
            .I(N__11100));
    LocalMux I__1190 (
            .O(N__11115),
            .I(N__11095));
    LocalMux I__1189 (
            .O(N__11112),
            .I(N__11095));
    Span12Mux_v I__1188 (
            .O(N__11109),
            .I(N__11090));
    Span4Mux_v I__1187 (
            .O(N__11106),
            .I(N__11081));
    LocalMux I__1186 (
            .O(N__11103),
            .I(N__11081));
    Span4Mux_s2_h I__1185 (
            .O(N__11100),
            .I(N__11081));
    Span4Mux_v I__1184 (
            .O(N__11095),
            .I(N__11081));
    InMux I__1183 (
            .O(N__11094),
            .I(N__11076));
    InMux I__1182 (
            .O(N__11093),
            .I(N__11076));
    Odrv12 I__1181 (
            .O(N__11090),
            .I(uart_data_rdy_debug_c));
    Odrv4 I__1180 (
            .O(N__11081),
            .I(uart_data_rdy_debug_c));
    LocalMux I__1179 (
            .O(N__11076),
            .I(uart_data_rdy_debug_c));
    SRMux I__1178 (
            .O(N__11069),
            .I(N__11065));
    SRMux I__1177 (
            .O(N__11068),
            .I(N__11062));
    LocalMux I__1176 (
            .O(N__11065),
            .I(\frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    LocalMux I__1175 (
            .O(N__11062),
            .I(\frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__1174 (
            .O(N__11057),
            .I(N__11054));
    LocalMux I__1173 (
            .O(N__11054),
            .I(N__11051));
    Span4Mux_s3_h I__1172 (
            .O(N__11051),
            .I(N__11046));
    InMux I__1171 (
            .O(N__11050),
            .I(N__11041));
    InMux I__1170 (
            .O(N__11049),
            .I(N__11041));
    Odrv4 I__1169 (
            .O(N__11046),
            .I(uart_drone_data_1));
    LocalMux I__1168 (
            .O(N__11041),
            .I(uart_drone_data_1));
    InMux I__1167 (
            .O(N__11036),
            .I(N__11033));
    LocalMux I__1166 (
            .O(N__11033),
            .I(N__11030));
    Span4Mux_s3_h I__1165 (
            .O(N__11030),
            .I(N__11025));
    InMux I__1164 (
            .O(N__11029),
            .I(N__11020));
    InMux I__1163 (
            .O(N__11028),
            .I(N__11020));
    Odrv4 I__1162 (
            .O(N__11025),
            .I(uart_drone_data_3));
    LocalMux I__1161 (
            .O(N__11020),
            .I(uart_drone_data_3));
    InMux I__1160 (
            .O(N__11015),
            .I(N__11012));
    LocalMux I__1159 (
            .O(N__11012),
            .I(uart_drone_data_0));
    InMux I__1158 (
            .O(N__11009),
            .I(N__11006));
    LocalMux I__1157 (
            .O(N__11006),
            .I(uart_drone_data_5));
    InMux I__1156 (
            .O(N__11003),
            .I(N__10999));
    InMux I__1155 (
            .O(N__11002),
            .I(N__10996));
    LocalMux I__1154 (
            .O(N__10999),
            .I(N__10993));
    LocalMux I__1153 (
            .O(N__10996),
            .I(\reset_module_System.countZ0Z_5 ));
    Odrv4 I__1152 (
            .O(N__10993),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__1151 (
            .O(N__10988),
            .I(N__10984));
    InMux I__1150 (
            .O(N__10987),
            .I(N__10981));
    LocalMux I__1149 (
            .O(N__10984),
            .I(N__10978));
    LocalMux I__1148 (
            .O(N__10981),
            .I(\reset_module_System.countZ0Z_4 ));
    Odrv4 I__1147 (
            .O(N__10978),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__1146 (
            .O(N__10973),
            .I(N__10969));
    InMux I__1145 (
            .O(N__10972),
            .I(N__10966));
    LocalMux I__1144 (
            .O(N__10969),
            .I(\reset_module_System.countZ0Z_18 ));
    LocalMux I__1143 (
            .O(N__10966),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__1142 (
            .O(N__10961),
            .I(N__10957));
    InMux I__1141 (
            .O(N__10960),
            .I(N__10954));
    LocalMux I__1140 (
            .O(N__10957),
            .I(N__10951));
    LocalMux I__1139 (
            .O(N__10954),
            .I(\reset_module_System.countZ0Z_16 ));
    Odrv4 I__1138 (
            .O(N__10951),
            .I(\reset_module_System.countZ0Z_16 ));
    CascadeMux I__1137 (
            .O(N__10946),
            .I(\reset_module_System.reset6_3_cascade_ ));
    InMux I__1136 (
            .O(N__10943),
            .I(N__10940));
    LocalMux I__1135 (
            .O(N__10940),
            .I(\reset_module_System.reset6_13 ));
    InMux I__1134 (
            .O(N__10937),
            .I(N__10934));
    LocalMux I__1133 (
            .O(N__10934),
            .I(N__10930));
    InMux I__1132 (
            .O(N__10933),
            .I(N__10927));
    Odrv12 I__1131 (
            .O(N__10930),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__1130 (
            .O(N__10927),
            .I(\reset_module_System.countZ0Z_12 ));
    CascadeMux I__1129 (
            .O(N__10922),
            .I(\reset_module_System.reset6_17_cascade_ ));
    InMux I__1128 (
            .O(N__10919),
            .I(N__10916));
    LocalMux I__1127 (
            .O(N__10916),
            .I(\reset_module_System.reset6_11 ));
    InMux I__1126 (
            .O(N__10913),
            .I(N__10910));
    LocalMux I__1125 (
            .O(N__10910),
            .I(N__10906));
    InMux I__1124 (
            .O(N__10909),
            .I(N__10903));
    Odrv4 I__1123 (
            .O(N__10906),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__1122 (
            .O(N__10903),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__1121 (
            .O(N__10898),
            .I(N__10895));
    LocalMux I__1120 (
            .O(N__10895),
            .I(N__10891));
    InMux I__1119 (
            .O(N__10894),
            .I(N__10888));
    Odrv4 I__1118 (
            .O(N__10891),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__1117 (
            .O(N__10888),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__1116 (
            .O(N__10883),
            .I(N__10879));
    InMux I__1115 (
            .O(N__10882),
            .I(N__10876));
    LocalMux I__1114 (
            .O(N__10879),
            .I(\reset_module_System.countZ0Z_20 ));
    LocalMux I__1113 (
            .O(N__10876),
            .I(\reset_module_System.countZ0Z_20 ));
    CascadeMux I__1112 (
            .O(N__10871),
            .I(\reset_module_System.reset6_15_cascade_ ));
    InMux I__1111 (
            .O(N__10868),
            .I(N__10865));
    LocalMux I__1110 (
            .O(N__10865),
            .I(N__10862));
    Odrv12 I__1109 (
            .O(N__10862),
            .I(\reset_module_System.count_1_2 ));
    CascadeMux I__1108 (
            .O(N__10859),
            .I(N__10855));
    InMux I__1107 (
            .O(N__10858),
            .I(N__10852));
    InMux I__1106 (
            .O(N__10855),
            .I(N__10849));
    LocalMux I__1105 (
            .O(N__10852),
            .I(N__10846));
    LocalMux I__1104 (
            .O(N__10849),
            .I(\reset_module_System.countZ0Z_2 ));
    Odrv12 I__1103 (
            .O(N__10846),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__1102 (
            .O(N__10841),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__1101 (
            .O(N__10838),
            .I(bfn_2_19_0_));
    InMux I__1100 (
            .O(N__10835),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__1099 (
            .O(N__10832),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__1098 (
            .O(N__10829),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__1097 (
            .O(N__10826),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__1096 (
            .O(N__10823),
            .I(N__10819));
    InMux I__1095 (
            .O(N__10822),
            .I(N__10816));
    LocalMux I__1094 (
            .O(N__10819),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__1093 (
            .O(N__10816),
            .I(\reset_module_System.countZ0Z_13 ));
    CascadeMux I__1092 (
            .O(N__10811),
            .I(N__10808));
    InMux I__1091 (
            .O(N__10808),
            .I(N__10802));
    InMux I__1090 (
            .O(N__10807),
            .I(N__10802));
    LocalMux I__1089 (
            .O(N__10802),
            .I(\reset_module_System.countZ0Z_19 ));
    CascadeMux I__1088 (
            .O(N__10799),
            .I(N__10795));
    InMux I__1087 (
            .O(N__10798),
            .I(N__10790));
    InMux I__1086 (
            .O(N__10795),
            .I(N__10790));
    LocalMux I__1085 (
            .O(N__10790),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__1084 (
            .O(N__10787),
            .I(N__10783));
    InMux I__1083 (
            .O(N__10786),
            .I(N__10780));
    LocalMux I__1082 (
            .O(N__10783),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__1081 (
            .O(N__10780),
            .I(\reset_module_System.countZ0Z_15 ));
    InMux I__1080 (
            .O(N__10775),
            .I(N__10771));
    InMux I__1079 (
            .O(N__10774),
            .I(N__10768));
    LocalMux I__1078 (
            .O(N__10771),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__1077 (
            .O(N__10768),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__1076 (
            .O(N__10763),
            .I(N__10759));
    InMux I__1075 (
            .O(N__10762),
            .I(N__10756));
    LocalMux I__1074 (
            .O(N__10759),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__1073 (
            .O(N__10756),
            .I(\reset_module_System.countZ0Z_10 ));
    CascadeMux I__1072 (
            .O(N__10751),
            .I(N__10748));
    InMux I__1071 (
            .O(N__10748),
            .I(N__10744));
    InMux I__1070 (
            .O(N__10747),
            .I(N__10741));
    LocalMux I__1069 (
            .O(N__10744),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__1068 (
            .O(N__10741),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__1067 (
            .O(N__10736),
            .I(N__10730));
    InMux I__1066 (
            .O(N__10735),
            .I(N__10730));
    LocalMux I__1065 (
            .O(N__10730),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__1064 (
            .O(N__10727),
            .I(N__10723));
    InMux I__1063 (
            .O(N__10726),
            .I(N__10720));
    LocalMux I__1062 (
            .O(N__10723),
            .I(N__10717));
    LocalMux I__1061 (
            .O(N__10720),
            .I(\reset_module_System.countZ0Z_8 ));
    Odrv4 I__1060 (
            .O(N__10717),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__1059 (
            .O(N__10712),
            .I(N__10708));
    InMux I__1058 (
            .O(N__10711),
            .I(N__10705));
    LocalMux I__1057 (
            .O(N__10708),
            .I(N__10702));
    LocalMux I__1056 (
            .O(N__10705),
            .I(\reset_module_System.countZ0Z_7 ));
    Odrv4 I__1055 (
            .O(N__10702),
            .I(\reset_module_System.countZ0Z_7 ));
    CascadeMux I__1054 (
            .O(N__10697),
            .I(N__10693));
    InMux I__1053 (
            .O(N__10696),
            .I(N__10690));
    InMux I__1052 (
            .O(N__10693),
            .I(N__10687));
    LocalMux I__1051 (
            .O(N__10690),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__1050 (
            .O(N__10687),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__1049 (
            .O(N__10682),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__1048 (
            .O(N__10679),
            .I(\reset_module_System.count_1_cry_7 ));
    InMux I__1047 (
            .O(N__10676),
            .I(bfn_2_18_0_));
    InMux I__1046 (
            .O(N__10673),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__1045 (
            .O(N__10670),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__1044 (
            .O(N__10667),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__1043 (
            .O(N__10664),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__1042 (
            .O(N__10661),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__1041 (
            .O(N__10658),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__1040 (
            .O(N__10655),
            .I(N__10651));
    InMux I__1039 (
            .O(N__10654),
            .I(N__10646));
    LocalMux I__1038 (
            .O(N__10651),
            .I(N__10643));
    InMux I__1037 (
            .O(N__10650),
            .I(N__10640));
    InMux I__1036 (
            .O(N__10649),
            .I(N__10637));
    LocalMux I__1035 (
            .O(N__10646),
            .I(\frame_dron_decoder_1.stateZ0Z_0 ));
    Odrv4 I__1034 (
            .O(N__10643),
            .I(\frame_dron_decoder_1.stateZ0Z_0 ));
    LocalMux I__1033 (
            .O(N__10640),
            .I(\frame_dron_decoder_1.stateZ0Z_0 ));
    LocalMux I__1032 (
            .O(N__10637),
            .I(\frame_dron_decoder_1.stateZ0Z_0 ));
    InMux I__1031 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__1030 (
            .O(N__10625),
            .I(\frame_dron_decoder_1.state_ns_i_a2_1_2_0 ));
    CascadeMux I__1029 (
            .O(N__10622),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    InMux I__1028 (
            .O(N__10619),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__1027 (
            .O(N__10616),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__1026 (
            .O(N__10613),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__1025 (
            .O(N__10610),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__1024 (
            .O(N__10607),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__1023 (
            .O(N__10604),
            .I(\frame_dron_decoder_1.un1_WDT_cry_8 ));
    InMux I__1022 (
            .O(N__10601),
            .I(N__10597));
    InMux I__1021 (
            .O(N__10600),
            .I(N__10594));
    LocalMux I__1020 (
            .O(N__10597),
            .I(\frame_dron_decoder_1.WDTZ0Z_10 ));
    LocalMux I__1019 (
            .O(N__10594),
            .I(\frame_dron_decoder_1.WDTZ0Z_10 ));
    InMux I__1018 (
            .O(N__10589),
            .I(\frame_dron_decoder_1.un1_WDT_cry_9 ));
    CascadeMux I__1017 (
            .O(N__10586),
            .I(N__10582));
    InMux I__1016 (
            .O(N__10585),
            .I(N__10578));
    InMux I__1015 (
            .O(N__10582),
            .I(N__10573));
    InMux I__1014 (
            .O(N__10581),
            .I(N__10573));
    LocalMux I__1013 (
            .O(N__10578),
            .I(\frame_dron_decoder_1.WDTZ0Z_11 ));
    LocalMux I__1012 (
            .O(N__10573),
            .I(\frame_dron_decoder_1.WDTZ0Z_11 ));
    InMux I__1011 (
            .O(N__10568),
            .I(\frame_dron_decoder_1.un1_WDT_cry_10 ));
    InMux I__1010 (
            .O(N__10565),
            .I(N__10560));
    InMux I__1009 (
            .O(N__10564),
            .I(N__10555));
    InMux I__1008 (
            .O(N__10563),
            .I(N__10555));
    LocalMux I__1007 (
            .O(N__10560),
            .I(\frame_dron_decoder_1.WDTZ0Z_12 ));
    LocalMux I__1006 (
            .O(N__10555),
            .I(\frame_dron_decoder_1.WDTZ0Z_12 ));
    InMux I__1005 (
            .O(N__10550),
            .I(\frame_dron_decoder_1.un1_WDT_cry_11 ));
    InMux I__1004 (
            .O(N__10547),
            .I(N__10543));
    InMux I__1003 (
            .O(N__10546),
            .I(N__10540));
    LocalMux I__1002 (
            .O(N__10543),
            .I(\frame_dron_decoder_1.WDTZ0Z_13 ));
    LocalMux I__1001 (
            .O(N__10540),
            .I(\frame_dron_decoder_1.WDTZ0Z_13 ));
    InMux I__1000 (
            .O(N__10535),
            .I(\frame_dron_decoder_1.un1_WDT_cry_12 ));
    InMux I__999 (
            .O(N__10532),
            .I(N__10525));
    InMux I__998 (
            .O(N__10531),
            .I(N__10525));
    InMux I__997 (
            .O(N__10530),
            .I(N__10522));
    LocalMux I__996 (
            .O(N__10525),
            .I(N__10519));
    LocalMux I__995 (
            .O(N__10522),
            .I(\frame_dron_decoder_1.WDTZ0Z_14 ));
    Odrv4 I__994 (
            .O(N__10519),
            .I(\frame_dron_decoder_1.WDTZ0Z_14 ));
    InMux I__993 (
            .O(N__10514),
            .I(\frame_dron_decoder_1.un1_WDT_cry_13 ));
    InMux I__992 (
            .O(N__10511),
            .I(\frame_dron_decoder_1.un1_WDT_cry_14 ));
    CascadeMux I__991 (
            .O(N__10508),
            .I(N__10505));
    InMux I__990 (
            .O(N__10505),
            .I(N__10498));
    InMux I__989 (
            .O(N__10504),
            .I(N__10498));
    InMux I__988 (
            .O(N__10503),
            .I(N__10495));
    LocalMux I__987 (
            .O(N__10498),
            .I(N__10492));
    LocalMux I__986 (
            .O(N__10495),
            .I(\frame_dron_decoder_1.WDTZ0Z_15 ));
    Odrv4 I__985 (
            .O(N__10492),
            .I(\frame_dron_decoder_1.WDTZ0Z_15 ));
    InMux I__984 (
            .O(N__10487),
            .I(N__10484));
    LocalMux I__983 (
            .O(N__10484),
            .I(\frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3 ));
    CascadeMux I__982 (
            .O(N__10481),
            .I(N__10478));
    InMux I__981 (
            .O(N__10478),
            .I(N__10473));
    InMux I__980 (
            .O(N__10477),
            .I(N__10470));
    InMux I__979 (
            .O(N__10476),
            .I(N__10467));
    LocalMux I__978 (
            .O(N__10473),
            .I(\frame_dron_decoder_1.stateZ0Z_1 ));
    LocalMux I__977 (
            .O(N__10470),
            .I(\frame_dron_decoder_1.stateZ0Z_1 ));
    LocalMux I__976 (
            .O(N__10467),
            .I(\frame_dron_decoder_1.stateZ0Z_1 ));
    InMux I__975 (
            .O(N__10460),
            .I(N__10456));
    InMux I__974 (
            .O(N__10459),
            .I(N__10453));
    LocalMux I__973 (
            .O(N__10456),
            .I(N__10449));
    LocalMux I__972 (
            .O(N__10453),
            .I(N__10446));
    InMux I__971 (
            .O(N__10452),
            .I(N__10443));
    Span4Mux_v I__970 (
            .O(N__10449),
            .I(N__10436));
    Span4Mux_h I__969 (
            .O(N__10446),
            .I(N__10436));
    LocalMux I__968 (
            .O(N__10443),
            .I(N__10436));
    Span4Mux_v I__967 (
            .O(N__10436),
            .I(N__10433));
    Odrv4 I__966 (
            .O(N__10433),
            .I(uart_drone_data_4));
    CascadeMux I__965 (
            .O(N__10430),
            .I(\frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_ ));
    InMux I__964 (
            .O(N__10427),
            .I(N__10424));
    LocalMux I__963 (
            .O(N__10424),
            .I(N__10421));
    Odrv4 I__962 (
            .O(N__10421),
            .I(\frame_dron_decoder_1.state_ns_0_a3_0_3_3 ));
    InMux I__961 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__960 (
            .O(N__10415),
            .I(\frame_dron_decoder_1.WDTZ0Z_1 ));
    InMux I__959 (
            .O(N__10412),
            .I(\frame_dron_decoder_1.un1_WDT_cry_0 ));
    InMux I__958 (
            .O(N__10409),
            .I(N__10406));
    LocalMux I__957 (
            .O(N__10406),
            .I(\frame_dron_decoder_1.WDTZ0Z_2 ));
    InMux I__956 (
            .O(N__10403),
            .I(\frame_dron_decoder_1.un1_WDT_cry_1 ));
    InMux I__955 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__954 (
            .O(N__10397),
            .I(\frame_dron_decoder_1.WDTZ0Z_3 ));
    InMux I__953 (
            .O(N__10394),
            .I(\frame_dron_decoder_1.un1_WDT_cry_2 ));
    InMux I__952 (
            .O(N__10391),
            .I(N__10387));
    InMux I__951 (
            .O(N__10390),
            .I(N__10384));
    LocalMux I__950 (
            .O(N__10387),
            .I(\frame_dron_decoder_1.WDTZ0Z_4 ));
    LocalMux I__949 (
            .O(N__10384),
            .I(\frame_dron_decoder_1.WDTZ0Z_4 ));
    InMux I__948 (
            .O(N__10379),
            .I(\frame_dron_decoder_1.un1_WDT_cry_3 ));
    InMux I__947 (
            .O(N__10376),
            .I(N__10372));
    InMux I__946 (
            .O(N__10375),
            .I(N__10369));
    LocalMux I__945 (
            .O(N__10372),
            .I(\frame_dron_decoder_1.WDTZ0Z_5 ));
    LocalMux I__944 (
            .O(N__10369),
            .I(\frame_dron_decoder_1.WDTZ0Z_5 ));
    InMux I__943 (
            .O(N__10364),
            .I(\frame_dron_decoder_1.un1_WDT_cry_4 ));
    InMux I__942 (
            .O(N__10361),
            .I(N__10357));
    InMux I__941 (
            .O(N__10360),
            .I(N__10354));
    LocalMux I__940 (
            .O(N__10357),
            .I(\frame_dron_decoder_1.WDTZ0Z_6 ));
    LocalMux I__939 (
            .O(N__10354),
            .I(\frame_dron_decoder_1.WDTZ0Z_6 ));
    InMux I__938 (
            .O(N__10349),
            .I(\frame_dron_decoder_1.un1_WDT_cry_5 ));
    InMux I__937 (
            .O(N__10346),
            .I(N__10342));
    InMux I__936 (
            .O(N__10345),
            .I(N__10339));
    LocalMux I__935 (
            .O(N__10342),
            .I(\frame_dron_decoder_1.WDTZ0Z_7 ));
    LocalMux I__934 (
            .O(N__10339),
            .I(\frame_dron_decoder_1.WDTZ0Z_7 ));
    InMux I__933 (
            .O(N__10334),
            .I(\frame_dron_decoder_1.un1_WDT_cry_6 ));
    InMux I__932 (
            .O(N__10331),
            .I(N__10327));
    InMux I__931 (
            .O(N__10330),
            .I(N__10324));
    LocalMux I__930 (
            .O(N__10327),
            .I(\frame_dron_decoder_1.WDTZ0Z_8 ));
    LocalMux I__929 (
            .O(N__10324),
            .I(\frame_dron_decoder_1.WDTZ0Z_8 ));
    InMux I__928 (
            .O(N__10319),
            .I(bfn_2_15_0_));
    CascadeMux I__927 (
            .O(N__10316),
            .I(N__10312));
    InMux I__926 (
            .O(N__10315),
            .I(N__10309));
    InMux I__925 (
            .O(N__10312),
            .I(N__10306));
    LocalMux I__924 (
            .O(N__10309),
            .I(\frame_dron_decoder_1.WDTZ0Z_9 ));
    LocalMux I__923 (
            .O(N__10306),
            .I(\frame_dron_decoder_1.WDTZ0Z_9 ));
    CascadeMux I__922 (
            .O(N__10301),
            .I(\frame_dron_decoder_1.N_229_cascade_ ));
    InMux I__921 (
            .O(N__10298),
            .I(N__10295));
    LocalMux I__920 (
            .O(N__10295),
            .I(\frame_dron_decoder_1.state_ns_i_a2_0_2_0 ));
    InMux I__919 (
            .O(N__10292),
            .I(N__10289));
    LocalMux I__918 (
            .O(N__10289),
            .I(\frame_dron_decoder_1.N_231 ));
    CascadeMux I__917 (
            .O(N__10286),
            .I(\frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_ ));
    InMux I__916 (
            .O(N__10283),
            .I(N__10280));
    LocalMux I__915 (
            .O(N__10280),
            .I(\frame_dron_decoder_1.state_ns_0_a3_0_3_1 ));
    InMux I__914 (
            .O(N__10277),
            .I(N__10273));
    InMux I__913 (
            .O(N__10276),
            .I(N__10264));
    LocalMux I__912 (
            .O(N__10273),
            .I(N__10261));
    InMux I__911 (
            .O(N__10272),
            .I(N__10256));
    InMux I__910 (
            .O(N__10271),
            .I(N__10256));
    InMux I__909 (
            .O(N__10270),
            .I(N__10247));
    InMux I__908 (
            .O(N__10269),
            .I(N__10247));
    InMux I__907 (
            .O(N__10268),
            .I(N__10247));
    InMux I__906 (
            .O(N__10267),
            .I(N__10247));
    LocalMux I__905 (
            .O(N__10264),
            .I(\frame_dron_decoder_1.N_249 ));
    Odrv4 I__904 (
            .O(N__10261),
            .I(\frame_dron_decoder_1.N_249 ));
    LocalMux I__903 (
            .O(N__10256),
            .I(\frame_dron_decoder_1.N_249 ));
    LocalMux I__902 (
            .O(N__10247),
            .I(\frame_dron_decoder_1.N_249 ));
    CascadeMux I__901 (
            .O(N__10238),
            .I(N__10234));
    CascadeMux I__900 (
            .O(N__10237),
            .I(N__10231));
    InMux I__899 (
            .O(N__10234),
            .I(N__10228));
    InMux I__898 (
            .O(N__10231),
            .I(N__10225));
    LocalMux I__897 (
            .O(N__10228),
            .I(\frame_dron_decoder_1.stateZ0Z_3 ));
    LocalMux I__896 (
            .O(N__10225),
            .I(\frame_dron_decoder_1.stateZ0Z_3 ));
    CascadeMux I__895 (
            .O(N__10220),
            .I(N__10216));
    InMux I__894 (
            .O(N__10219),
            .I(N__10213));
    InMux I__893 (
            .O(N__10216),
            .I(N__10210));
    LocalMux I__892 (
            .O(N__10213),
            .I(\frame_dron_decoder_1.WDT10_0_i ));
    LocalMux I__891 (
            .O(N__10210),
            .I(\frame_dron_decoder_1.WDT10_0_i ));
    InMux I__890 (
            .O(N__10205),
            .I(N__10202));
    LocalMux I__889 (
            .O(N__10202),
            .I(\frame_dron_decoder_1.WDTZ0Z_0 ));
    InMux I__888 (
            .O(N__10199),
            .I(N__10196));
    LocalMux I__887 (
            .O(N__10196),
            .I(\frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4 ));
    CascadeMux I__886 (
            .O(N__10193),
            .I(\frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_ ));
    CascadeMux I__885 (
            .O(N__10190),
            .I(\frame_dron_decoder_1.WDT10lt14_0_cascade_ ));
    InMux I__884 (
            .O(N__10187),
            .I(N__10184));
    LocalMux I__883 (
            .O(N__10184),
            .I(\frame_dron_decoder_1.WDT10lt14_0 ));
    InMux I__882 (
            .O(N__10181),
            .I(N__10178));
    LocalMux I__881 (
            .O(N__10178),
            .I(\frame_dron_decoder_1.WDT10lto13_1 ));
    CascadeMux I__880 (
            .O(N__10175),
            .I(N__10172));
    InMux I__879 (
            .O(N__10172),
            .I(N__10169));
    LocalMux I__878 (
            .O(N__10169),
            .I(N__10165));
    InMux I__877 (
            .O(N__10168),
            .I(N__10162));
    Odrv4 I__876 (
            .O(N__10165),
            .I(\frame_dron_decoder_1.stateZ0Z_7 ));
    LocalMux I__875 (
            .O(N__10162),
            .I(\frame_dron_decoder_1.stateZ0Z_7 ));
    CascadeMux I__874 (
            .O(N__10157),
            .I(\frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_ ));
    CascadeMux I__873 (
            .O(N__10154),
            .I(\frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_ ));
    InMux I__872 (
            .O(N__10151),
            .I(N__10145));
    InMux I__871 (
            .O(N__10150),
            .I(N__10145));
    LocalMux I__870 (
            .O(N__10145),
            .I(\frame_dron_decoder_1.stateZ0Z_2 ));
    CascadeMux I__869 (
            .O(N__10142),
            .I(N__10139));
    InMux I__868 (
            .O(N__10139),
            .I(N__10133));
    InMux I__867 (
            .O(N__10138),
            .I(N__10133));
    LocalMux I__866 (
            .O(N__10133),
            .I(\frame_dron_decoder_1.stateZ0Z_5 ));
    InMux I__865 (
            .O(N__10130),
            .I(N__10124));
    InMux I__864 (
            .O(N__10129),
            .I(N__10124));
    LocalMux I__863 (
            .O(N__10124),
            .I(\frame_dron_decoder_1.stateZ0Z_4 ));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\scaler_3.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\scaler_3.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\scaler_2.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\scaler_2.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\scaler_1.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\scaler_1.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_13 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_13 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_13 ),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_10_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_27_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\uart_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_11_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_28_0_));
    defparam IN_MUX_bfv_11_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_29_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_11_29_0_));
    defparam IN_MUX_bfv_11_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_30_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_11_30_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\frame_dron_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_2_15_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__24213),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB pc_frame_decoder_dv_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__20138),
            .GLOBALBUFFEROUTPUT(pc_frame_decoder_dv_0_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23969),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_228_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \frame_dron_decoder_1.state_2_LC_1_13_0 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_2_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_2_LC_1_13_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \frame_dron_decoder_1.state_2_LC_1_13_0  (
            .in0(N__10150),
            .in1(N__11137),
            .in2(N__10238),
            .in3(N__10267),
            .lcout(\frame_dron_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25295),
            .ce(),
            .sr(N__24755));
    defparam \frame_dron_decoder_1.state_5_LC_1_13_2 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_5_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_5_LC_1_13_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \frame_dron_decoder_1.state_5_LC_1_13_2  (
            .in0(N__10151),
            .in1(N__11141),
            .in2(N__10142),
            .in3(N__10269),
            .lcout(\frame_dron_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25295),
            .ce(),
            .sr(N__24755));
    defparam \frame_dron_decoder_1.state_4_LC_1_13_3 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_4_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_4_LC_1_13_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \frame_dron_decoder_1.state_4_LC_1_13_3  (
            .in0(N__10268),
            .in1(N__10138),
            .in2(N__11148),
            .in3(N__10129),
            .lcout(\frame_dron_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25295),
            .ce(),
            .sr(N__24755));
    defparam \frame_dron_decoder_1.state_7_LC_1_13_7 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_7_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_7_LC_1_13_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \frame_dron_decoder_1.state_7_LC_1_13_7  (
            .in0(N__10270),
            .in1(N__10168),
            .in2(N__11149),
            .in3(N__10130),
            .lcout(\frame_dron_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25295),
            .ce(),
            .sr(N__24755));
    defparam \frame_dron_decoder_1.WDT_RNIMRG3_4_LC_1_14_0 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNIMRG3_4_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNIMRG3_4_LC_1_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \frame_dron_decoder_1.WDT_RNIMRG3_4_LC_1_14_0  (
            .in0(N__10330),
            .in1(N__10375),
            .in2(N__10316),
            .in3(N__10390),
            .lcout(\frame_dron_decoder_1.WDT_RNIMRG3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.WDT_RNI6TFJ1_10_LC_1_14_1 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNI6TFJ1_10_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNI6TFJ1_10_LC_1_14_1 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \frame_dron_decoder_1.WDT_RNI6TFJ1_10_LC_1_14_1  (
            .in0(N__10600),
            .in1(N__10546),
            .in2(N__10586),
            .in3(N__10564),
            .lcout(),
            .ltout(\frame_dron_decoder_1.WDT_RNI6TFJ1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.WDT_RNIA5HI2_7_LC_1_14_2 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNIA5HI2_7_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNIA5HI2_7_LC_1_14_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \frame_dron_decoder_1.WDT_RNIA5HI2_7_LC_1_14_2  (
            .in0(N__10345),
            .in1(N__10199),
            .in2(N__10193),
            .in3(N__10181),
            .lcout(\frame_dron_decoder_1.WDT10lt14_0 ),
            .ltout(\frame_dron_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.WDT_RNI3A9C3_15_LC_1_14_3 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNI3A9C3_15_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNI3A9C3_15_LC_1_14_3 .LUT_INIT=16'b0011001100111111;
    LogicCell40 \frame_dron_decoder_1.WDT_RNI3A9C3_15_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__10504),
            .in2(N__10190),
            .in3(N__10531),
            .lcout(\frame_dron_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.WDT_RNICPRL3_15_LC_1_14_6 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNICPRL3_15_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNICPRL3_15_LC_1_14_6 .LUT_INIT=16'b0000001100010011;
    LogicCell40 \frame_dron_decoder_1.WDT_RNICPRL3_15_LC_1_14_6  (
            .in0(N__10532),
            .in1(N__11136),
            .in2(N__10508),
            .in3(N__10187),
            .lcout(\frame_dron_decoder_1.N_249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.WDT_RNI05KQ_6_LC_1_14_7 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_RNI05KQ_6_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.WDT_RNI05KQ_6_LC_1_14_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \frame_dron_decoder_1.WDT_RNI05KQ_6_LC_1_14_7  (
            .in0(N__10581),
            .in1(N__10563),
            .in2(_gnd_net_),
            .in3(N__10360),
            .lcout(\frame_dron_decoder_1.WDT10lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_6_LC_1_15_0 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_6_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_6_LC_1_15_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \frame_dron_decoder_1.state_6_LC_1_15_0  (
            .in0(N__11233),
            .in1(N__11135),
            .in2(N__10175),
            .in3(N__10271),
            .lcout(\frame_dron_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25290),
            .ce(),
            .sr(N__24764));
    defparam \frame_dron_decoder_1.state_RNIOTUU_6_LC_1_15_4 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNIOTUU_6_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNIOTUU_6_LC_1_15_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \frame_dron_decoder_1.state_RNIOTUU_6_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__11232),
            .in2(_gnd_net_),
            .in3(N__10649),
            .lcout(\frame_dron_decoder_1.state_ns_i_a2_0_2_0 ),
            .ltout(\frame_dron_decoder_1.state_ns_i_a2_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_3_0_LC_1_15_5 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_3_0_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_3_0_LC_1_15_5 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \frame_dron_decoder_1.state_RNO_3_0_LC_1_15_5  (
            .in0(N__10452),
            .in1(N__11389),
            .in2(N__10157),
            .in3(N__10487),
            .lcout(),
            .ltout(\frame_dron_decoder_1.state_ns_i_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_0_0_LC_1_15_6 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_0_0_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_0_0_LC_1_15_6 .LUT_INIT=16'b0101100000000000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_0_0_LC_1_15_6  (
            .in0(N__11390),
            .in1(N__10628),
            .in2(N__10154),
            .in3(N__11178),
            .lcout(),
            .ltout(\frame_dron_decoder_1.N_229_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_0_LC_1_15_7 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_0_LC_1_15_7 .SEQ_MODE=4'b1001;
    defparam \frame_dron_decoder_1.state_0_LC_1_15_7 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \frame_dron_decoder_1.state_0_LC_1_15_7  (
            .in0(N__10272),
            .in1(N__10292),
            .in2(N__10301),
            .in3(N__10654),
            .lcout(\frame_dron_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25290),
            .ce(),
            .sr(N__24764));
    defparam \frame_dron_decoder_1.state_1_LC_1_16_2 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_1_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_1_LC_1_16_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \frame_dron_decoder_1.state_1_LC_1_16_2  (
            .in0(N__10283),
            .in1(N__11183),
            .in2(N__10481),
            .in3(N__10277),
            .lcout(\frame_dron_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25285),
            .ce(),
            .sr(N__24770));
    defparam \frame_dron_decoder_1.state_RNO_1_0_LC_1_16_5 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_1_0_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_1_0_LC_1_16_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_1_0_LC_1_16_5  (
            .in0(N__10476),
            .in1(N__10298),
            .in2(_gnd_net_),
            .in3(N__11134),
            .lcout(\frame_dron_decoder_1.N_231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_1_1_LC_1_17_6 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_1_1_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_1_1_LC_1_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_1_1_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__11388),
            .in2(_gnd_net_),
            .in3(N__11057),
            .lcout(),
            .ltout(\frame_dron_decoder_1.state_ns_0_a3_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_0_1_LC_1_17_7 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_0_1_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_0_1_LC_1_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_0_1_LC_1_17_7  (
            .in0(N__10460),
            .in1(N__10655),
            .in2(N__10286),
            .in3(N__11036),
            .lcout(\frame_dron_decoder_1.state_ns_0_a3_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_4_LC_2_12_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_2_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11264),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25296),
            .ce(N__11351),
            .sr(N__11330));
    defparam \uart_drone.data_esr_2_LC_2_12_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_2_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11630),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25296),
            .ce(N__11351),
            .sr(N__11330));
    defparam \frame_dron_decoder_1.state_3_LC_2_13_3 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_3_LC_2_13_3 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.state_3_LC_2_13_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \frame_dron_decoder_1.state_3_LC_2_13_3  (
            .in0(N__11182),
            .in1(N__10427),
            .in2(N__10237),
            .in3(N__10276),
            .lcout(\frame_dron_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25294),
            .ce(),
            .sr(N__24750));
    defparam \frame_dron_decoder_1.WDT_0_LC_2_14_0 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_0_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_0_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_0_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__10205),
            .in2(N__10220),
            .in3(N__10219),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_0 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_1_LC_2_14_1 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_1_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_1_LC_2_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_1_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__10412),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_0 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_1 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_2_LC_2_14_2 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_2_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_2_LC_2_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_2_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__10409),
            .in2(_gnd_net_),
            .in3(N__10403),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_1 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_2 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_3_LC_2_14_3 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_3_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_3_LC_2_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_3_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__10400),
            .in2(_gnd_net_),
            .in3(N__10394),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_2 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_3 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_4_LC_2_14_4 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_4_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_4_LC_2_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_4_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__10391),
            .in2(_gnd_net_),
            .in3(N__10379),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_3 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_4 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_5_LC_2_14_5 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_5_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_5_LC_2_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_5_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__10376),
            .in2(_gnd_net_),
            .in3(N__10364),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_4 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_5 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_6_LC_2_14_6 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_6_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_6_LC_2_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_6_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__10361),
            .in2(_gnd_net_),
            .in3(N__10349),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_5 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_6 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_7_LC_2_14_7 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_7_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_7_LC_2_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_7_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__10346),
            .in2(_gnd_net_),
            .in3(N__10334),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_6 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_7 ),
            .clk(N__25291),
            .ce(),
            .sr(N__11069));
    defparam \frame_dron_decoder_1.WDT_8_LC_2_15_0 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_8_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_8_LC_2_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_8_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__10331),
            .in2(_gnd_net_),
            .in3(N__10319),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_8 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_9_LC_2_15_1 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_9_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_9_LC_2_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_9_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__10315),
            .in2(_gnd_net_),
            .in3(N__10604),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_8 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_9 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_10_LC_2_15_2 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_10_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_10_LC_2_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_10_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__10601),
            .in2(_gnd_net_),
            .in3(N__10589),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_9 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_10 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_11_LC_2_15_3 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_11_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_11_LC_2_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_11_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__10585),
            .in2(_gnd_net_),
            .in3(N__10568),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_10 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_11 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_12_LC_2_15_4 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_12_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_12_LC_2_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_12_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__10565),
            .in2(_gnd_net_),
            .in3(N__10550),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_11 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_12 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_13_LC_2_15_5 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_13_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_13_LC_2_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_13_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__10547),
            .in2(_gnd_net_),
            .in3(N__10535),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_12 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_13 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_14_LC_2_15_6 .C_ON=1'b1;
    defparam \frame_dron_decoder_1.WDT_14_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_14_LC_2_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \frame_dron_decoder_1.WDT_14_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__10530),
            .in2(_gnd_net_),
            .in3(N__10514),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\frame_dron_decoder_1.un1_WDT_cry_13 ),
            .carryout(\frame_dron_decoder_1.un1_WDT_cry_14 ),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.WDT_15_LC_2_15_7 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.WDT_15_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.WDT_15_LC_2_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \frame_dron_decoder_1.WDT_15_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__10503),
            .in2(_gnd_net_),
            .in3(N__10511),
            .lcout(\frame_dron_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25286),
            .ce(),
            .sr(N__11068));
    defparam \frame_dron_decoder_1.state_ns_0_a3_0_1_3_LC_2_16_2 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_ns_0_a3_0_1_3_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_ns_0_a3_0_1_3_LC_2_16_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \frame_dron_decoder_1.state_ns_0_a3_0_1_3_LC_2_16_2  (
            .in0(N__11049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11028),
            .lcout(\frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3 ),
            .ltout(\frame_dron_decoder_1.state_ns_0_a3_0_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_0_3_LC_2_16_3 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_0_3_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_0_3_LC_2_16_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_0_3_LC_2_16_3  (
            .in0(N__10477),
            .in1(N__10459),
            .in2(N__10430),
            .in3(N__11379),
            .lcout(\frame_dron_decoder_1.state_ns_0_a3_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_RNO_2_0_LC_2_16_5 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_RNO_2_0_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_RNO_2_0_LC_2_16_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \frame_dron_decoder_1.state_RNO_2_0_LC_2_16_5  (
            .in0(N__11029),
            .in1(N__10650),
            .in2(_gnd_net_),
            .in3(N__11050),
            .lcout(\frame_dron_decoder_1.state_ns_i_a2_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_2_16_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_2_16_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_2_16_6  (
            .in0(N__12050),
            .in1(N__11439),
            .in2(_gnd_net_),
            .in3(N__24191),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_2_16_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_2_16_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_2_16_7  (
            .in0(N__11440),
            .in1(_gnd_net_),
            .in2(N__10622),
            .in3(_gnd_net_),
            .lcout(\uart_drone.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_2_17_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_2_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__11546),
            .in2(N__11465),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_2_17_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_2_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__10858),
            .in2(_gnd_net_),
            .in3(N__10619),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_2_17_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_2_17_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_2_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__10894),
            .in2(_gnd_net_),
            .in3(N__10616),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_2_17_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_2_17_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_2_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__10987),
            .in2(_gnd_net_),
            .in3(N__10613),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_2_17_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_2_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__11002),
            .in2(_gnd_net_),
            .in3(N__10610),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_2_17_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_2_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__10909),
            .in2(_gnd_net_),
            .in3(N__10607),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_2_17_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_2_17_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_2_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__10711),
            .in2(_gnd_net_),
            .in3(N__10682),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_2_17_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_2_17_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_2_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__10726),
            .in2(_gnd_net_),
            .in3(N__10679),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__25277),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_2_18_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_2_18_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__10696),
            .in2(_gnd_net_),
            .in3(N__10676),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_2_18_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_2_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__10762),
            .in2(_gnd_net_),
            .in3(N__10673),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_2_18_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_2_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__10747),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_2_18_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_2_18_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_2_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__10933),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_2_18_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_2_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__10823),
            .in2(_gnd_net_),
            .in3(N__10664),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_2_18_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_2_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__10774),
            .in2(_gnd_net_),
            .in3(N__10661),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_2_18_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_2_18_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_2_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__10787),
            .in2(_gnd_net_),
            .in3(N__10658),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_2_18_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_2_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__10960),
            .in2(_gnd_net_),
            .in3(N__10841),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__25272),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_2_19_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_2_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__10735),
            .in2(_gnd_net_),
            .in3(N__10838),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__25268),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_2_19_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_2_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__10973),
            .in2(_gnd_net_),
            .in3(N__10835),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__25268),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_2_19_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_2_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \reset_module_System.count_19_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10811),
            .in3(N__10832),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__25268),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_2_19_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_2_19_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_2_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__10883),
            .in2(_gnd_net_),
            .in3(N__10829),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__25268),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_2_19_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_2_19_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_2_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__10798),
            .in2(_gnd_net_),
            .in3(N__10826),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25268),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_2_19_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_2_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_2_19_5  (
            .in0(N__10822),
            .in1(N__10807),
            .in2(N__10799),
            .in3(N__10786),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_2_19_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_2_19_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_2_19_6  (
            .in0(N__10775),
            .in1(N__10763),
            .in2(N__10751),
            .in3(N__10736),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_2_19_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_2_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_2_19_7  (
            .in0(N__10727),
            .in1(N__10712),
            .in2(N__10697),
            .in3(N__11003),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_2_20_1 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_2_20_1 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_2_20_1  (
            .in0(N__11544),
            .in1(N__11522),
            .in2(N__11507),
            .in3(N__11482),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25262),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_2_20_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_2_20_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__10988),
            .in2(_gnd_net_),
            .in3(N__11457),
            .lcout(),
            .ltout(\reset_module_System.reset6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_2_20_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_2_20_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_2_20_3  (
            .in0(N__10972),
            .in1(N__10961),
            .in2(N__10946),
            .in3(N__10943),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_2_20_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_2_20_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_2_20_4  (
            .in0(N__10937),
            .in1(N__11543),
            .in2(N__10922),
            .in3(N__10919),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_2_20_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_2_20_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_2_20_5  (
            .in0(N__10913),
            .in1(N__10898),
            .in2(N__10859),
            .in3(N__10882),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(\reset_module_System.reset6_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_2_20_6 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_2_20_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \reset_module_System.count_2_LC_2_20_6  (
            .in0(N__11483),
            .in1(N__11506),
            .in2(N__10871),
            .in3(N__10868),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25262),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_2_21_4 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_2_21_4 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.state_1_LC_2_21_4  (
            .in0(N__12056),
            .in1(N__11564),
            .in2(N__12491),
            .in3(N__24919),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25254),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_rdy_LC_3_14_3 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_3_14_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_3_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__12039),
            .in2(_gnd_net_),
            .in3(N__11441),
            .lcout(uart_data_rdy_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25287),
            .ce(),
            .sr(N__24751));
    defparam \frame_dron_decoder_1.source_data_valid_LC_3_14_6 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.source_data_valid_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \frame_dron_decoder_1.source_data_valid_LC_3_14_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \frame_dron_decoder_1.source_data_valid_LC_3_14_6  (
            .in0(N__11206),
            .in1(N__11240),
            .in2(_gnd_net_),
            .in3(N__11121),
            .lcout(drone_frame_decoder_data_rdy_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25287),
            .ce(),
            .sr(N__24751));
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_1 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \frame_dron_decoder_1.state_ns_i_a2_2_0_0_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__11357),
            .in2(_gnd_net_),
            .in3(N__11093),
            .lcout(),
            .ltout(\frame_dron_decoder_1.state_ns_i_a2_2_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_LC_3_15_2 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.state_ns_i_a2_2_0_LC_3_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \frame_dron_decoder_1.state_ns_i_a2_2_0_LC_3_15_2  (
            .in0(N__11009),
            .in1(N__11195),
            .in2(N__11186),
            .in3(N__11015),
            .lcout(\frame_dron_decoder_1.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \frame_dron_decoder_1.source_data_valid_2_sqmuxa_i_LC_3_15_4 .C_ON=1'b0;
    defparam \frame_dron_decoder_1.source_data_valid_2_sqmuxa_i_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \frame_dron_decoder_1.source_data_valid_2_sqmuxa_i_LC_3_15_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \frame_dron_decoder_1.source_data_valid_2_sqmuxa_i_LC_3_15_4  (
            .in0(N__11094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24897),
            .lcout(\frame_dron_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_3_15_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_3_15_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_3_15_6  (
            .in0(N__11656),
            .in1(N__15267),
            .in2(_gnd_net_),
            .in3(N__24896),
            .lcout(\uart_pc.state_srsts_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_1_LC_3_16_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_3_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11296),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_esr_3_LC_3_16_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_3_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11281),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_esr_0_LC_3_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_3_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_3_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11311),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_esr_5_LC_3_16_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_3_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_3_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone.data_esr_5_LC_3_16_5  (
            .in0(N__11830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_esr_6_LC_3_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_3_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11608),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_esr_7_LC_3_16_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_3_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_3_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11644),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25278),
            .ce(N__11347),
            .sr(N__11326));
    defparam \uart_drone.data_Aux_0_LC_3_17_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_3_17_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_0_LC_3_17_0  (
            .in0(N__12040),
            .in1(N__11246),
            .in2(N__11312),
            .in3(N__11855),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25273),
            .ce(),
            .sr(N__11801));
    defparam \uart_drone.data_Aux_1_LC_3_17_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_3_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_3_17_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_3_17_1  (
            .in0(N__11856),
            .in1(N__11420),
            .in2(N__11297),
            .in3(N__12041),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25273),
            .ce(),
            .sr(N__11801));
    defparam \uart_drone.data_Aux_3_LC_3_17_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_3_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_3_17_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_3_17_3  (
            .in0(N__11857),
            .in1(N__11414),
            .in2(N__11282),
            .in3(N__12042),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25273),
            .ce(),
            .sr(N__11801));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_3_17_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_3_17_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_3_17_5  (
            .in0(N__12314),
            .in1(N__12371),
            .in2(_gnd_net_),
            .in3(N__12447),
            .lcout(),
            .ltout(\uart_drone.data_Auxce_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_4_LC_3_17_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_3_17_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \uart_drone.data_Aux_4_LC_3_17_6  (
            .in0(N__12043),
            .in1(N__11257),
            .in2(N__11267),
            .in3(N__11858),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25273),
            .ce(),
            .sr(N__11801));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_3_17_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_3_17_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_3_17_7  (
            .in0(N__12313),
            .in1(N__12370),
            .in2(_gnd_net_),
            .in3(N__12446),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_3_18_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_3_18_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_3_18_0  (
            .in0(N__12310),
            .in1(N__12365),
            .in2(_gnd_net_),
            .in3(N__12443),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_3_18_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_3_18_1 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_3_18_1  (
            .in0(N__12169),
            .in1(N__12527),
            .in2(N__11939),
            .in3(N__11580),
            .lcout(\uart_drone.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_3_18_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_3_18_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_3_18_2  (
            .in0(N__12311),
            .in1(N__12366),
            .in2(_gnd_net_),
            .in3(N__12444),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_3_18_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_3_18_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_3_18_3  (
            .in0(N__12445),
            .in1(_gnd_net_),
            .in2(N__12374),
            .in3(N__12312),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_3_18_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_3_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_3_18_4  (
            .in0(N__11581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12170),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_3_18_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_3_18_5 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_3_18_5  (
            .in0(N__11405),
            .in1(N__12528),
            .in2(N__11408),
            .in3(N__12135),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_3_19_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_3_19_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_3_19_0  (
            .in0(N__11759),
            .in1(N__11710),
            .in2(N__11762),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_3_19_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_3_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__11582),
            .in2(_gnd_net_),
            .in3(N__11399),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_3_19_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_3_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__12174),
            .in2(_gnd_net_),
            .in3(N__11396),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_3_19_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_3_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__11938),
            .in2(_gnd_net_),
            .in3(N__11393),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_3_19_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_3_19_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_3_19_6  (
            .in0(N__11735),
            .in1(N__24120),
            .in2(N__12245),
            .in3(N__11594),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25263),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_3_19_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_3_19_7 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_2_LC_3_19_7  (
            .in0(N__11588),
            .in1(N__12241),
            .in2(N__24169),
            .in3(N__11734),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25263),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_3_20_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_3_20_0 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_3_20_0  (
            .in0(N__12051),
            .in1(N__11562),
            .in2(N__12209),
            .in3(N__24899),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_3_20_1 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_3_20_1 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \uart_drone.state_2_LC_3_20_1  (
            .in0(N__11941),
            .in1(N__12176),
            .in2(N__11567),
            .in3(N__11563),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25255),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_3_20_2 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_3_20_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_3_20_2  (
            .in0(N__11520),
            .in1(N__11501),
            .in2(_gnd_net_),
            .in3(N__11480),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25255),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_3_20_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__11545),
            .in2(_gnd_net_),
            .in3(N__11461),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_3_20_4 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_3_20_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_3_20_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_3_20_4  (
            .in0(N__11521),
            .in1(N__11502),
            .in2(N__11486),
            .in3(N__11481),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25255),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_3_20_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_3_20_6 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_3_20_6  (
            .in0(N__12129),
            .in1(N__11940),
            .in2(N__12208),
            .in3(N__12175),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_3_21_0 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_3_21_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uart_drone.bit_Count_1_LC_3_21_0  (
            .in0(N__12442),
            .in1(N__12363),
            .in2(N__12473),
            .in3(N__12385),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25250),
            .ce(),
            .sr(N__24781));
    defparam \uart_drone.bit_Count_0_LC_3_21_3 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_3_21_3 .LUT_INIT=16'b0100010001100100;
    LogicCell40 \uart_drone.bit_Count_0_LC_3_21_3  (
            .in0(N__12469),
            .in1(N__12441),
            .in2(N__12137),
            .in3(N__12082),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25250),
            .ce(),
            .sr(N__24781));
    defparam \uart_drone_sync.Q_0__0_LC_4_2_2 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_4_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11699),
            .lcout(uart_input_debug_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25304),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_4_2_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_4_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12263),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25304),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_4_13_5 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_4_13_5 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_4_13_5  (
            .in0(N__11660),
            .in1(N__15247),
            .in2(N__11693),
            .in3(N__24918),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25288),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_2_LC_4_14_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_4_14_5 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_4_14_5  (
            .in0(N__12980),
            .in1(N__15246),
            .in2(N__11692),
            .in3(N__24898),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_4_14_6 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_4_14_6 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_pc.state_2_LC_4_14_6  (
            .in0(N__11688),
            .in1(N__13183),
            .in2(N__11669),
            .in3(N__13040),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25282),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_4_15_7 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_4_15_7 .LUT_INIT=16'b1111110101010101;
    LogicCell40 \uart_pc.state_0_LC_4_15_7  (
            .in0(N__11666),
            .in1(N__13184),
            .in2(N__12836),
            .in3(N__12816),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25279),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_7_LC_4_16_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_4_16_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_4_16_0  (
            .in0(N__12015),
            .in1(N__11867),
            .in2(N__11645),
            .in3(N__12083),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25274),
            .ce(),
            .sr(N__11800));
    defparam \uart_drone.data_Aux_2_LC_4_16_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_4_16_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_4_16_6  (
            .in0(N__11810),
            .in1(N__12014),
            .in2(N__11626),
            .in3(N__11866),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25274),
            .ce(),
            .sr(N__11800));
    defparam \uart_drone.data_Aux_6_LC_4_17_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_4_17_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_4_17_1  (
            .in0(N__11816),
            .in1(N__12017),
            .in2(N__11609),
            .in3(N__11860),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25269),
            .ce(),
            .sr(N__11793));
    defparam \uart_drone.data_Aux_5_LC_4_17_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_4_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_4_17_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_5_LC_4_17_3  (
            .in0(N__11873),
            .in1(N__12016),
            .in2(N__11831),
            .in3(N__11859),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25269),
            .ce(),
            .sr(N__11793));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_4_18_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_4_18_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_4_18_1  (
            .in0(N__12296),
            .in1(N__12373),
            .in2(_gnd_net_),
            .in3(N__12449),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_4_18_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_4_18_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_4_18_3  (
            .in0(N__12295),
            .in1(N__12372),
            .in2(_gnd_net_),
            .in3(N__12448),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_4_18_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_4_18_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_4_18_7  (
            .in0(N__12136),
            .in1(N__12529),
            .in2(_gnd_net_),
            .in3(N__24903),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_4_19_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_4_19_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_4_19_2 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \uart_drone.timer_Count_0_LC_4_19_2  (
            .in0(N__24118),
            .in1(N__11761),
            .in2(N__11741),
            .in3(N__12238),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25256),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_4_19_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_4_19_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_4_19_3  (
            .in0(N__11937),
            .in1(N__12523),
            .in2(N__24199),
            .in3(N__11887),
            .lcout(\uart_drone.N_143 ),
            .ltout(\uart_drone.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_4_19_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_4_19_4 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \uart_drone.timer_Count_4_LC_4_19_4  (
            .in0(N__11771),
            .in1(N__24168),
            .in2(N__11765),
            .in3(N__11740),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25256),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_4_19_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_4_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__11760),
            .in2(_gnd_net_),
            .in3(N__11711),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_4_19_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_4_19_7 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_4_19_7  (
            .in0(N__12239),
            .in1(N__11739),
            .in2(N__11714),
            .in3(N__24119),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25256),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_4_20_0 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_4_20_0 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \uart_drone.state_4_LC_4_20_0  (
            .in0(N__24116),
            .in1(N__12218),
            .in2(N__12134),
            .in3(N__12240),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25251),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_4_20_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_4_20_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_4_20_2  (
            .in0(N__11927),
            .in1(N__12078),
            .in2(_gnd_net_),
            .in3(N__12173),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(\uart_drone.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_4_20_3 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_4_20_3 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \uart_drone.state_3_LC_4_20_3  (
            .in0(N__12200),
            .in1(N__12182),
            .in2(N__12212),
            .in3(N__24117),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25251),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_4_20_5 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_4_20_5 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_4_20_5  (
            .in0(N__12172),
            .in1(N__12118),
            .in2(N__12207),
            .in3(N__11928),
            .lcout(\uart_drone.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_4_20_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_4_20_6 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_4_20_6  (
            .in0(N__11926),
            .in1(N__12171),
            .in2(N__12133),
            .in3(N__12522),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_4_21_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_4_21_0 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_4_21_0  (
            .in0(N__12122),
            .in1(N__12468),
            .in2(_gnd_net_),
            .in3(N__12077),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_4_21_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_4_21_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_4_21_2  (
            .in0(N__12281),
            .in1(N__12345),
            .in2(_gnd_net_),
            .in3(N__12422),
            .lcout(\uart_drone.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_4_21_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_4_21_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_4_21_3  (
            .in0(N__12484),
            .in1(N__12013),
            .in2(_gnd_net_),
            .in3(N__24900),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_4_21_4 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_4_21_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_4_21_4 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_4_21_4  (
            .in0(N__11942),
            .in1(N__11891),
            .in2(N__11876),
            .in3(N__12530),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25244),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_4_21_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_4_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_4_21_6  (
            .in0(_gnd_net_),
            .in1(N__12467),
            .in2(_gnd_net_),
            .in3(N__12423),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_2_LC_4_22_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_4_22_5 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uart_drone.bit_Count_2_LC_4_22_5  (
            .in0(N__12392),
            .in1(N__12386),
            .in2(N__12309),
            .in3(N__12364),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25238),
            .ce(),
            .sr(N__24782));
    defparam \uart_drone_sync.aux_2__0__0_LC_5_2_3 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_5_2_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__13379),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25303),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_6_LC_5_9_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_5_9_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_6_LC_5_9_3  (
            .in0(N__12257),
            .in1(N__15266),
            .in2(N__14623),
            .in3(N__12869),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25297),
            .ce(),
            .sr(N__12575));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_10_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_10_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_5_10_2  (
            .in0(N__12702),
            .in1(N__12769),
            .in2(_gnd_net_),
            .in3(N__12623),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_10_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_5_10_4  (
            .in0(N__12701),
            .in1(N__12768),
            .in2(_gnd_net_),
            .in3(N__12622),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_5_11_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_5_11_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_5_11_0  (
            .in0(N__12776),
            .in1(N__15251),
            .in2(N__13348),
            .in3(N__12862),
            .lcout(\uart_pc.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_1_LC_5_11_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_5_11_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_1_LC_5_11_1  (
            .in0(N__12863),
            .in1(N__13363),
            .in2(N__15269),
            .in3(N__12251),
            .lcout(\uart_pc.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_2_LC_5_11_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_5_11_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_5_11_2  (
            .in0(N__12557),
            .in1(N__15252),
            .in2(N__13309),
            .in3(N__12864),
            .lcout(\uart_pc.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_3_LC_5_11_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_5_11_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_3_LC_5_11_3  (
            .in0(N__12865),
            .in1(N__13288),
            .in2(N__15270),
            .in3(N__12551),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_4_LC_5_11_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_5_11_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_5_11_4  (
            .in0(N__12539),
            .in1(N__15253),
            .in2(N__13331),
            .in3(N__12866),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_5_LC_5_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_5_11_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_5_LC_5_11_5  (
            .in0(N__12867),
            .in1(N__13273),
            .in2(N__15271),
            .in3(N__12545),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.data_Aux_7_LC_5_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_5_11_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_7_LC_5_11_7  (
            .in0(N__12868),
            .in1(N__13261),
            .in2(N__15272),
            .in3(N__12959),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25292),
            .ce(),
            .sr(N__12574));
    defparam \uart_pc.state_RNIEAGS_4_LC_5_12_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_5_12_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_5_12_0  (
            .in0(N__12919),
            .in1(N__12818),
            .in2(_gnd_net_),
            .in3(N__24901),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_12_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_5_12_1  (
            .in0(N__12756),
            .in1(N__12692),
            .in2(_gnd_net_),
            .in3(N__12618),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_12_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_12_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_5_12_2  (
            .in0(N__12619),
            .in1(_gnd_net_),
            .in2(N__12703),
            .in3(N__12757),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_12_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_12_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_5_12_3  (
            .in0(N__12759),
            .in1(N__12699),
            .in2(_gnd_net_),
            .in3(N__12621),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_12_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_12_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_5_12_4  (
            .in0(N__12620),
            .in1(_gnd_net_),
            .in2(N__12704),
            .in3(N__12758),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_12_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_12_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_5_12_7  (
            .in0(N__12755),
            .in1(N__12691),
            .in2(_gnd_net_),
            .in3(N__12617),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_5_13_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_5_13_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_2_LC_5_13_2  (
            .in0(N__12722),
            .in1(N__12700),
            .in2(N__12770),
            .in3(N__12716),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25283),
            .ce(),
            .sr(N__24741));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_5_14_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_5_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_5_14_1  (
            .in0(N__12754),
            .in1(N__12670),
            .in2(_gnd_net_),
            .in3(N__12597),
            .lcout(\uart_pc.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_5_14_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_5_14_2 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_5_14_2  (
            .in0(N__13174),
            .in1(N__13039),
            .in2(N__12920),
            .in3(N__12817),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(\uart_pc.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_5_14_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_5_14_3 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__12916),
            .in2(N__12725),
            .in3(N__12950),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_5_14_7 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_5_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__12634),
            .in2(_gnd_net_),
            .in3(N__12598),
            .lcout(\uart_pc.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_1_LC_5_15_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_5_15_2 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uart_pc.bit_Count_1_LC_5_15_2  (
            .in0(N__12690),
            .in1(N__12715),
            .in2(N__12647),
            .in3(N__12616),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25275),
            .ce(),
            .sr(N__24746));
    defparam \uart_pc.bit_Count_0_LC_5_15_6 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_5_15_6 .LUT_INIT=16'b0000111100100000;
    LogicCell40 \uart_pc.bit_Count_0_LC_5_15_6  (
            .in0(N__12917),
            .in1(N__12957),
            .in2(N__12646),
            .in3(N__12615),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25275),
            .ce(),
            .sr(N__24746));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_16_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_16_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_5_16_0  (
            .in0(N__13032),
            .in1(N__13118),
            .in2(N__13181),
            .in3(N__12807),
            .lcout(\uart_pc.state_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_5_16_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_5_16_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_5_16_1  (
            .in0(N__12905),
            .in1(N__13173),
            .in2(N__12989),
            .in3(N__13035),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_5_16_2 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_5_16_2 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_pc.state_3_LC_5_16_2  (
            .in0(N__12987),
            .in1(N__12928),
            .in2(N__12992),
            .in3(N__24193),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25270),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_16_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_5_16_3 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_5_16_3  (
            .in0(N__12904),
            .in1(N__13169),
            .in2(N__12988),
            .in3(N__13034),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_5_16_5 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_5_16_5 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \uart_pc.state_4_LC_5_16_5  (
            .in0(N__12929),
            .in1(N__24192),
            .in2(N__12918),
            .in3(N__13091),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25270),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_16_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_16_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_5_16_6  (
            .in0(N__13033),
            .in1(_gnd_net_),
            .in2(N__13182),
            .in3(N__12958),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_5_17_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_5_17_0 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \uart_pc.timer_Count_0_LC_5_17_0  (
            .in0(N__13225),
            .in1(N__13087),
            .in2(N__24212),
            .in3(N__13053),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25264),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_17_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_5_17_1 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_5_17_1  (
            .in0(N__12812),
            .in1(N__12829),
            .in2(N__13205),
            .in3(N__12909),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_17_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_5_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__13224),
            .in2(_gnd_net_),
            .in3(N__13238),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_17_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_5_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__13030),
            .in2(_gnd_net_),
            .in3(N__13116),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_17_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_5_17_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_5_17_6  (
            .in0(N__13159),
            .in1(N__12811),
            .in2(N__12779),
            .in3(N__24194),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_5_17_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_5_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_5_17_7 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_5_17_7  (
            .in0(N__13054),
            .in1(N__24195),
            .in2(N__13247),
            .in3(N__13244),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25264),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_18_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_5_18_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_5_18_0  (
            .in0(N__13223),
            .in1(N__13237),
            .in2(N__13226),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_18_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_5_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__13117),
            .in2(_gnd_net_),
            .in3(N__13196),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_18_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_5_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__13031),
            .in2(_gnd_net_),
            .in3(N__13193),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_18_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_5_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__13165),
            .in2(_gnd_net_),
            .in3(N__13190),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_5_18_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_5_18_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_pc.timer_Count_4_LC_5_18_4  (
            .in0(N__13064),
            .in1(N__13090),
            .in2(N__13187),
            .in3(N__24184),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25257),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_5_18_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_5_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_5_18_5 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_pc.timer_Count_2_LC_5_18_5  (
            .in0(N__13124),
            .in1(N__13088),
            .in2(N__24210),
            .in3(N__13062),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25257),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_5_18_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_5_18_7 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_pc.timer_Count_3_LC_5_18_7  (
            .in0(N__13097),
            .in1(N__13089),
            .in2(N__24211),
            .in3(N__13063),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25257),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_7_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_7_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13391),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25302),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_7_2_4 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_7_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13385),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25301),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_esr_1_LC_7_10_0 .C_ON=1'b0;
    defparam \uart_pc.data_esr_1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_1_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_1_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13370),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25289),
            .ce(N__14601),
            .sr(N__14808));
    defparam \uart_pc.data_esr_0_LC_7_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_esr_0_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_0_LC_7_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_0_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13352),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25289),
            .ce(N__14601),
            .sr(N__14808));
    defparam \uart_pc.data_esr_4_LC_7_11_0 .C_ON=1'b0;
    defparam \uart_pc.data_esr_4_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_4_LC_7_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_4_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13327),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25284),
            .ce(N__14606),
            .sr(N__14810));
    defparam \uart_pc.data_esr_2_LC_7_11_2 .C_ON=1'b0;
    defparam \uart_pc.data_esr_2_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_2_LC_7_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_2_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13310),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25284),
            .ce(N__14606),
            .sr(N__14810));
    defparam \uart_pc.data_esr_3_LC_7_11_3 .C_ON=1'b0;
    defparam \uart_pc.data_esr_3_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_3_LC_7_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_3_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13292),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25284),
            .ce(N__14606),
            .sr(N__14810));
    defparam \uart_pc.data_esr_5_LC_7_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_esr_5_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_5_LC_7_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc.data_esr_5_LC_7_11_5  (
            .in0(N__13277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25284),
            .ce(N__14606),
            .sr(N__14810));
    defparam \uart_pc.data_esr_7_LC_7_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_esr_7_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_7_LC_7_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc.data_esr_7_LC_7_11_7  (
            .in0(N__13262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25284),
            .ce(N__14606),
            .sr(N__14810));
    defparam \uart_frame_decoder.state_1_1_LC_7_12_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_1_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_1_LC_7_12_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uart_frame_decoder.state_1_1_LC_7_12_3  (
            .in0(N__13763),
            .in1(N__23932),
            .in2(N__13772),
            .in3(N__23904),
            .lcout(\uart_frame_decoder.state_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25280),
            .ce(),
            .sr(N__24740));
    defparam \uart_frame_decoder.state_1_RNIC4PK_6_LC_7_13_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIC4PK_6_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIC4PK_6_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIC4PK_6_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__13852),
            .in2(_gnd_net_),
            .in3(N__23823),
            .lcout(\uart_frame_decoder.source_offset1data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIE6PK_8_LC_7_13_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIE6PK_8_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIE6PK_8_LC_7_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIE6PK_8_LC_7_13_3  (
            .in0(N__23824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13807),
            .lcout(\uart_frame_decoder.source_offset3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNID5PK_7_LC_7_13_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNID5PK_7_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNID5PK_7_LC_7_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNID5PK_7_LC_7_13_5  (
            .in0(N__23825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13828),
            .lcout(\uart_frame_decoder.source_offset2data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIAIVT_7_LC_7_13_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIAIVT_7_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIAIVT_7_LC_7_13_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_frame_decoder.state_1_RNIAIVT_7_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13415),
            .in3(N__24904),
            .lcout(\uart_frame_decoder.source_offset2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI9HVT_6_LC_7_14_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI9HVT_6_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI9HVT_6_LC_7_14_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNI9HVT_6_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__13840),
            .in2(_gnd_net_),
            .in3(N__24905),
            .lcout(\uart_frame_decoder.source_offset1data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIBJVT_8_LC_7_14_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIBJVT_8_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIBJVT_8_LC_7_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNIBJVT_8_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__13792),
            .in2(_gnd_net_),
            .in3(N__24906),
            .lcout(\uart_frame_decoder.source_offset3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_0_LC_7_15_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_0_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_0_LC_7_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_0_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__13412),
            .in2(N__13961),
            .in3(N__13960),
            .lcout(\uart_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_1_LC_7_15_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_1_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_1_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_1_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__13406),
            .in2(_gnd_net_),
            .in3(N__13400),
            .lcout(\uart_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_2_LC_7_15_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_2_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_2_LC_7_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_2_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__13397),
            .in2(_gnd_net_),
            .in3(N__13448),
            .lcout(\uart_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_3_LC_7_15_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_3_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_3_LC_7_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_3_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__13445),
            .in2(_gnd_net_),
            .in3(N__13439),
            .lcout(\uart_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_4_LC_7_15_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_4_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_4_LC_7_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_4_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__13907),
            .in2(_gnd_net_),
            .in3(N__13436),
            .lcout(\uart_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_5_LC_7_15_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_5_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_5_LC_7_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_5_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__13934),
            .in2(_gnd_net_),
            .in3(N__13433),
            .lcout(\uart_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_6_LC_7_15_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_6_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_6_LC_7_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_6_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__14111),
            .in2(_gnd_net_),
            .in3(N__13430),
            .lcout(\uart_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_7_LC_7_15_7 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_7_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_7_LC_7_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_7_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__14042),
            .in2(_gnd_net_),
            .in3(N__13427),
            .lcout(\uart_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__25265),
            .ce(),
            .sr(N__13889));
    defparam \uart_frame_decoder.WDT_8_LC_7_16_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_8_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_8_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_8_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__13946),
            .in2(_gnd_net_),
            .in3(N__13424),
            .lcout(\uart_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_9_LC_7_16_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_9_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_9_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_9_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__13921),
            .in2(_gnd_net_),
            .in3(N__13421),
            .lcout(\uart_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_10_LC_7_16_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_10_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_10_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_10_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__14084),
            .in2(_gnd_net_),
            .in3(N__13418),
            .lcout(\uart_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_11_LC_7_16_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_11_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_11_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_11_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__14099),
            .in2(_gnd_net_),
            .in3(N__13463),
            .lcout(\uart_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_12_LC_7_16_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_12_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_12_LC_7_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_12_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__14057),
            .in2(_gnd_net_),
            .in3(N__13460),
            .lcout(\uart_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_13_LC_7_16_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_13_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_13_LC_7_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_13_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__14071),
            .in2(_gnd_net_),
            .in3(N__13457),
            .lcout(\uart_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_14_LC_7_16_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_14_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_14_LC_7_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_14_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__14008),
            .in2(_gnd_net_),
            .in3(N__13454),
            .lcout(\uart_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.WDT_15_LC_7_16_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_15_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_15_LC_7_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_frame_decoder.WDT_15_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__13981),
            .in2(_gnd_net_),
            .in3(N__13451),
            .lcout(\uart_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25258),
            .ce(),
            .sr(N__13885));
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_7_17_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_0_LC_7_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21103),
            .lcout(frame_decoder_OFF1data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_7_17_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_1_LC_7_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20974),
            .lcout(frame_decoder_OFF1data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_7_17_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_2_LC_7_17_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_2_LC_7_17_2  (
            .in0(N__20898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF1data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_7_17_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_3_LC_7_17_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_3_LC_7_17_3  (
            .in0(N__20812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF1data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_7_17_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_4_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20727),
            .lcout(frame_decoder_OFF1data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_7_17_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_5_LC_7_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_5_LC_7_17_5  (
            .in0(N__26360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF1data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_7_17_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_6_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20632),
            .lcout(frame_decoder_OFF1data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_7_17_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset1data_esr_7_LC_7_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset1data_esr_7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20527),
            .lcout(frame_decoder_OFF1data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25252),
            .ce(N__13475),
            .sr(N__24756));
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_7_18_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_0_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_0_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(frame_decoder_CH1data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_7_18_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_1_LC_7_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_1_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20975),
            .lcout(frame_decoder_CH1data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_7_18_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_2_LC_7_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_2_LC_7_18_2  (
            .in0(N__20899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH1data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_7_18_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_3_LC_7_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_3_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20813),
            .lcout(frame_decoder_CH1data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_7_18_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_4_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_4_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20716),
            .lcout(frame_decoder_CH1data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_7_18_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_5_LC_7_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_5_LC_7_18_5  (
            .in0(N__26361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH1data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_7_18_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_6_LC_7_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_6_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20633),
            .lcout(frame_decoder_CH1data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25245),
            .ce(N__14312),
            .sr(N__24759));
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_7_19_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH1data_esr_7_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH1data_esr_7_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20536),
            .lcout(frame_decoder_CH1data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25239),
            .ce(N__14308),
            .sr(N__24765));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_7_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_7_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_7_20_7  (
            .in0(N__26102),
            .in1(N__14327),
            .in2(_gnd_net_),
            .in3(N__15421),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_7_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14981),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25228),
            .ce(N__21739),
            .sr(N__24774));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_7_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_7_21_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_7_21_4  (
            .in0(N__23594),
            .in1(_gnd_net_),
            .in2(N__22771),
            .in3(N__22330),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_7_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_7_21_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_7_21_5  (
            .in0(N__19418),
            .in1(N__22705),
            .in2(_gnd_net_),
            .in3(N__23592),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_7_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_7_21_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_7_21_6  (
            .in0(N__23593),
            .in1(_gnd_net_),
            .in2(N__22770),
            .in3(N__19417),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_7_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_7_21_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_7_21_7  (
            .in0(N__23086),
            .in1(N__22704),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_7_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_7_22_1 .LUT_INIT=16'b0100101000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_7_22_1  (
            .in0(N__22188),
            .in1(N__26071),
            .in2(N__23192),
            .in3(N__25800),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_22_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_22_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_7_22_2  (
            .in0(N__24920),
            .in1(N__22189),
            .in2(N__13478),
            .in3(N__23589),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25224),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_22_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_7_22_3  (
            .in0(N__23160),
            .in1(N__26072),
            .in2(N__25807),
            .in3(N__22693),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIE3D21_LC_7_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIE3D21_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIE3D21_LC_7_22_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIE3D21_LC_7_22_6  (
            .in0(N__15626),
            .in1(N__22239),
            .in2(N__22195),
            .in3(N__23156),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_162_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_7_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_7_23_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_7_23_0  (
            .in0(N__23508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14510),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIGD613_LC_7_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIGD613_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIGD613_LC_7_23_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIGD613_LC_7_23_1  (
            .in0(N__14512),
            .in1(N__15997),
            .in2(_gnd_net_),
            .in3(N__23510),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_7_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_7_23_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__15404),
            .in2(N__22695),
            .in3(N__25931),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_7_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_7_23_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13484),
            .in3(N__23506),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_7_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_7_23_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22190),
            .in3(N__14351),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_7_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_7_23_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13481),
            .in3(N__23505),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_7_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_7_23_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_7_23_6  (
            .in0(N__23507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14509),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_7_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_7_23_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_7_23_7  (
            .in0(N__14511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23509),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR7352_3_LC_7_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR7352_3_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR7352_3_LC_7_24_0 .LUT_INIT=16'b1101001000101101;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR7352_3_LC_7_24_0  (
            .in0(N__18637),
            .in1(N__19988),
            .in2(N__22511),
            .in3(N__16124),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI60223_3_LC_7_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI60223_3_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI60223_3_LC_7_24_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI60223_3_LC_7_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13499),
            .in3(N__15763),
            .lcout(\ppm_encoder_1.init_pulses_RNI60223Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_7_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_7_24_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_7_24_2  (
            .in0(N__22649),
            .in1(N__22503),
            .in2(_gnd_net_),
            .in3(N__23511),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_7_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_7_24_3 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_7_24_3  (
            .in0(N__23512),
            .in1(_gnd_net_),
            .in2(N__22510),
            .in3(N__22650),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_1_LC_7_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_7_24_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_7_24_4  (
            .in0(_gnd_net_),
            .in1(N__19989),
            .in2(_gnd_net_),
            .in3(N__25542),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25214),
            .ce(),
            .sr(N__24787));
    defparam \ppm_encoder_1.throttle_2_LC_7_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_7_24_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_7_24_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_7_24_5  (
            .in0(N__25543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13496),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25214),
            .ce(),
            .sr(N__24787));
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_7_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_7_24_6 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ppm_encoder_1.throttle_RNIR7352_2_LC_7_24_6  (
            .in0(N__13494),
            .in1(N__22136),
            .in2(N__18665),
            .in3(N__16123),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_7_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_7_24_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_7_24_7  (
            .in0(N__26063),
            .in1(N__25808),
            .in2(_gnd_net_),
            .in3(N__13495),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_7_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_7_25_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_7_25_0  (
            .in0(N__22345),
            .in1(N__23655),
            .in2(N__14525),
            .in3(N__16139),
            .lcout(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_6_LC_7_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_7_25_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_7_25_1 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_7_25_1  (
            .in0(N__19515),
            .in1(N__19700),
            .in2(N__13625),
            .in3(N__15674),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25208),
            .ce(),
            .sr(N__24793));
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_7_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_7_25_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIERUS_6_LC_7_25_2  (
            .in0(N__22344),
            .in1(N__22779),
            .in2(_gnd_net_),
            .in3(N__23653),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_7_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_7_25_3 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_7_25_3  (
            .in0(N__23656),
            .in1(N__22414),
            .in2(N__16147),
            .in3(N__14524),
            .lcout(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_7_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_7_25_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_7_25_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_7_25_4  (
            .in0(N__19699),
            .in1(N__13565),
            .in2(N__19549),
            .in3(N__15872),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25208),
            .ce(),
            .sr(N__24793));
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_7_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_7_25_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISFRP_13_LC_7_25_5  (
            .in0(N__23654),
            .in1(_gnd_net_),
            .in2(N__22822),
            .in3(N__22413),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_7_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_7_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(N__13553),
            .in2(N__14537),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_7_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_7_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_7_26_1  (
            .in0(_gnd_net_),
            .in1(N__13544),
            .in2(_gnd_net_),
            .in3(N__13535),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_7_26_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_7_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(N__14483),
            .in2(N__13532),
            .in3(N__13520),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_7_26_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_7_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_7_26_3  (
            .in0(_gnd_net_),
            .in1(N__13517),
            .in2(_gnd_net_),
            .in3(N__13508),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_7_26_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_7_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__14633),
            .in2(_gnd_net_),
            .in3(N__13505),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_7_26_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_7_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_7_26_5  (
            .in0(_gnd_net_),
            .in1(N__19721),
            .in2(_gnd_net_),
            .in3(N__13502),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_7_26_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_7_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__13643),
            .in2(N__13634),
            .in3(N__13616),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_7_26_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_7_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_7_26_7  (
            .in0(_gnd_net_),
            .in1(N__13613),
            .in2(_gnd_net_),
            .in3(N__13604),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_7_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_7_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(N__17402),
            .in2(_gnd_net_),
            .in3(N__13601),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_7_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_7_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(N__17354),
            .in2(_gnd_net_),
            .in3(N__13598),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_7_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_7_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__14408),
            .in2(_gnd_net_),
            .in3(N__13595),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_7_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_7_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(N__14447),
            .in2(_gnd_net_),
            .in3(N__13592),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_7_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_7_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__14576),
            .in2(_gnd_net_),
            .in3(N__13589),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_7_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_7_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(N__13586),
            .in2(N__13577),
            .in3(N__13556),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(N__13691),
            .in2(_gnd_net_),
            .in3(N__13679),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_7_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_7_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__14552),
            .in2(_gnd_net_),
            .in3(N__13676),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_7_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_7_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__13658),
            .in2(_gnd_net_),
            .in3(N__13673),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_7_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_7_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__13664),
            .in2(_gnd_net_),
            .in3(N__13670),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_7_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_7_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_7_28_2 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_7_28_2  (
            .in0(N__23707),
            .in1(N__15985),
            .in2(N__22840),
            .in3(N__13667),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_7_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_7_28_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_7_28_4  (
            .in0(N__23706),
            .in1(_gnd_net_),
            .in2(N__22839),
            .in3(N__16072),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_7_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_7_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_7_28_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_7_28_7  (
            .in0(N__15956),
            .in1(N__22827),
            .in2(_gnd_net_),
            .in3(N__23705),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_8_3_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_8_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_8_3_2  (
            .in0(N__13652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25300),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_8_4_3 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_8_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13721),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25299),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_8_4_6 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_8_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13727),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25299),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_8_5_0 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_8_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13715),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25298),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_8_8_0 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_8_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13709),
            .lcout(uart_input_pc_sync),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25293),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_10_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_8_10_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_8_10_0  (
            .in0(N__15221),
            .in1(N__15166),
            .in2(_gnd_net_),
            .in3(N__24173),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIE94V3_2_LC_8_10_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIE94V3_2_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIE94V3_2_LC_8_10_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_pc.timer_Count_RNIE94V3_2_LC_8_10_1  (
            .in0(N__15167),
            .in1(_gnd_net_),
            .in2(N__13700),
            .in3(_gnd_net_),
            .lcout(\uart_pc.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_8_11_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_8_11_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_0_LC_8_11_1  (
            .in0(N__13762),
            .in1(N__15317),
            .in2(_gnd_net_),
            .in3(N__14770),
            .lcout(\uart_frame_decoder.N_39_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_11_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_8_11_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_3_0_LC_8_11_3  (
            .in0(N__13761),
            .in1(N__15316),
            .in2(_gnd_net_),
            .in3(N__13781),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_RNO_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_8_11_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_8_11_4 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_1_0_LC_8_11_4  (
            .in0(N__13739),
            .in1(N__23953),
            .in2(N__13697),
            .in3(N__23931),
            .lcout(\uart_frame_decoder.state_1_ns_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_8_11_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_8_11_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__26310),
            .in2(_gnd_net_),
            .in3(N__21065),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIDPNH_1_LC_8_11_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIDPNH_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIDPNH_1_LC_8_11_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIDPNH_1_LC_8_11_6  (
            .in0(N__20483),
            .in1(N__13760),
            .in2(N__13694),
            .in3(N__20851),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_8_12_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_8_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_8_12_2  (
            .in0(N__26309),
            .in1(N__20850),
            .in2(N__20505),
            .in3(N__21069),
            .lcout(\uart_frame_decoder.N_138_4 ),
            .ltout(\uart_frame_decoder.N_138_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_8_12_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_8_12_3 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_1_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__14769),
            .in2(N__13775),
            .in3(_gnd_net_),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_8_12_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_8_12_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_2_0_LC_8_12_4  (
            .in0(N__15309),
            .in1(N__13759),
            .in2(N__14771),
            .in3(N__23826),
            .lcout(\uart_frame_decoder.state_1_RNO_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_8_12_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_8_12_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_8_12_6  (
            .in0(N__20599),
            .in1(N__20955),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_8_12_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_8_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_8_12_7  (
            .in0(N__23827),
            .in1(N__20673),
            .in2(N__13733),
            .in3(N__20766),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNI5CUL2_15_LC_8_13_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNI5CUL2_15_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNI5CUL2_15_LC_8_13_0 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \uart_frame_decoder.WDT_RNI5CUL2_15_LC_8_13_0  (
            .in0(N__14012),
            .in1(N__13985),
            .in2(N__23831),
            .in3(N__14021),
            .lcout(\uart_frame_decoder.N_85 ),
            .ltout(\uart_frame_decoder.N_85_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_3_LC_8_13_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_3_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_3_LC_8_13_1 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \uart_frame_decoder.state_1_3_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__14893),
            .in2(N__13730),
            .in3(N__21362),
            .lcout(\uart_frame_decoder.state_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_4_LC_8_13_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_4_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_4_LC_8_13_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uart_frame_decoder.state_1_4_LC_8_13_2  (
            .in0(N__14879),
            .in1(N__23845),
            .in2(_gnd_net_),
            .in3(N__23898),
            .lcout(\uart_frame_decoder.state_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_5_LC_8_13_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_5_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_5_LC_8_13_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \uart_frame_decoder.state_1_5_LC_8_13_3  (
            .in0(N__23899),
            .in1(N__17794),
            .in2(_gnd_net_),
            .in3(N__26381),
            .lcout(\uart_frame_decoder.state_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_6_LC_8_13_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_6_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_6_LC_8_13_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uart_frame_decoder.state_1_6_LC_8_13_4  (
            .in0(N__13853),
            .in1(N__17780),
            .in2(_gnd_net_),
            .in3(N__23900),
            .lcout(\uart_frame_decoder.state_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_7_LC_8_13_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_7_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_7_LC_8_13_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uart_frame_decoder.state_1_7_LC_8_13_5  (
            .in0(N__23901),
            .in1(N__13841),
            .in2(_gnd_net_),
            .in3(N__13829),
            .lcout(\uart_frame_decoder.state_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_8_LC_8_13_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_8_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_8_LC_8_13_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uart_frame_decoder.state_1_8_LC_8_13_6  (
            .in0(N__13817),
            .in1(N__13808),
            .in2(_gnd_net_),
            .in3(N__23902),
            .lcout(\uart_frame_decoder.state_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.state_1_9_LC_8_13_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_9_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_9_LC_8_13_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \uart_frame_decoder.state_1_9_LC_8_13_7  (
            .in0(N__23903),
            .in1(_gnd_net_),
            .in2(N__13796),
            .in3(N__14753),
            .lcout(\uart_frame_decoder.state_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25271),
            .ce(),
            .sr(N__24743));
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_8_14_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_0_LC_8_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_0_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21101),
            .lcout(frame_decoder_OFF2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_8_14_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_1_LC_8_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_1_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20988),
            .lcout(frame_decoder_OFF2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_8_14_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_2_LC_8_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_2_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20882),
            .lcout(frame_decoder_OFF2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_8_14_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_7_LC_8_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_7_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20507),
            .lcout(frame_decoder_OFF2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_8_14_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_4_LC_8_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_4_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20725),
            .lcout(frame_decoder_OFF2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_8_14_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_5_LC_8_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_5_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26342),
            .lcout(frame_decoder_OFF2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_8_14_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_6_LC_8_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_6_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20619),
            .lcout(frame_decoder_OFF2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_8_14_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset2data_esr_3_LC_8_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset2data_esr_3_LC_8_14_7  (
            .in0(N__20798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25266),
            .ce(N__13868),
            .sr(N__24747));
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_8_15_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_0_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_0_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21102),
            .lcout(frame_decoder_OFF3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_8_15_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_1_LC_8_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_1_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20989),
            .lcout(frame_decoder_OFF3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_8_15_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_2_LC_8_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_2_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20897),
            .lcout(frame_decoder_OFF3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_8_15_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_3_LC_8_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_3_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20811),
            .lcout(frame_decoder_OFF3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_8_15_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_4_LC_8_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_4_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20726),
            .lcout(frame_decoder_OFF3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_8_15_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_5_LC_8_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_5_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26359),
            .lcout(frame_decoder_OFF3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_8_15_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_6_LC_8_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_6_LC_8_15_6  (
            .in0(N__20620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_8_15_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset3data_esr_7_LC_8_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset3data_esr_7_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20526),
            .lcout(frame_decoder_OFF3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25259),
            .ce(N__14117),
            .sr(N__24752));
    defparam \uart_frame_decoder.WDT_RNIBI7E_6_LC_8_16_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIBI7E_6_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIBI7E_6_LC_8_16_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_frame_decoder.WDT_RNIBI7E_6_LC_8_16_0  (
            .in0(N__14055),
            .in1(N__14097),
            .in2(_gnd_net_),
            .in3(N__14110),
            .lcout(\uart_frame_decoder.WDT8lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_8_16_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIAGPB_10_LC_8_16_1 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \uart_frame_decoder.WDT_RNIAGPB_10_LC_8_16_1  (
            .in0(N__14098),
            .in1(N__14083),
            .in2(N__14072),
            .in3(N__14056),
            .lcout(),
            .ltout(\uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIM8N32_7_LC_8_16_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIM8N32_7_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIM8N32_7_LC_8_16_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \uart_frame_decoder.WDT_RNIM8N32_7_LC_8_16_2  (
            .in0(N__14041),
            .in1(N__13895),
            .in2(N__14030),
            .in3(N__14027),
            .lcout(\uart_frame_decoder.WDT8lt14_0 ),
            .ltout(\uart_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_8_16_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNI17K92_15_LC_8_16_3 .LUT_INIT=16'b0000001111111111;
    LogicCell40 \uart_frame_decoder.WDT_RNI17K92_15_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__14004),
            .in2(N__13988),
            .in3(N__13977),
            .lcout(\uart_frame_decoder.WDT8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_8_16_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_8_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_frame_decoder.WDT_RNIQAB11_4_LC_8_16_4  (
            .in0(N__13945),
            .in1(N__13933),
            .in2(N__13922),
            .in3(N__13906),
            .lcout(\uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_RNIHJ501_0_LC_8_16_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNIHJ501_0_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNIHJ501_0_LC_8_16_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uart_frame_decoder.count_RNIHJ501_0_LC_8_16_5  (
            .in0(N__16618),
            .in1(N__23816),
            .in2(_gnd_net_),
            .in3(N__15327),
            .lcout(\uart_frame_decoder.count_RNIHJ501Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_8_16_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_8_16_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_8_16_6  (
            .in0(N__23817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24902),
            .lcout(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_8_17_0 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__16536),
            .in2(N__16583),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\scaler_1.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_8_17_1 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_8_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__14231),
            .in2(N__14225),
            .in3(N__14216),
            .lcout(\scaler_1.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_0 ),
            .carryout(\scaler_1.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_8_17_2 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__14213),
            .in2(N__14207),
            .in3(N__14198),
            .lcout(\scaler_1.un3_source_data_0_cry_1_c_RNIISC11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_1 ),
            .carryout(\scaler_1.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_8_17_3 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__14195),
            .in2(N__14189),
            .in3(N__14180),
            .lcout(\scaler_1.un3_source_data_0_cry_2_c_RNIL0E11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_2 ),
            .carryout(\scaler_1.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_8_17_4 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__14177),
            .in2(N__14171),
            .in3(N__14162),
            .lcout(\scaler_1.un3_source_data_0_cry_3_c_RNIO4F11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_3 ),
            .carryout(\scaler_1.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_8_17_5 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__14159),
            .in2(N__14153),
            .in3(N__14144),
            .lcout(\scaler_1.un3_source_data_0_cry_4_c_RNIR8G11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_4 ),
            .carryout(\scaler_1.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_8_17_6 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__14141),
            .in2(N__14135),
            .in3(N__14126),
            .lcout(\scaler_1.un3_source_data_0_cry_5_c_RNIUCH11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_5 ),
            .carryout(\scaler_1.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_8_17_7 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_8_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__14288),
            .in2(_gnd_net_),
            .in3(N__14123),
            .lcout(\scaler_1.un3_source_data_0_cry_6_c_RNI1HI11 ),
            .ltout(),
            .carryin(\scaler_1.un3_source_data_0_cry_6 ),
            .carryout(\scaler_1.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_8_18_0 .C_ON=1'b1;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__14261),
            .in2(N__21850),
            .in3(N__14120),
            .lcout(\scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\scaler_1.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_8_18_1 .C_ON=1'b0;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_8_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14291),
            .lcout(\scaler_1.un3_source_data_0_cry_8_c_RNIPB6F ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_1_LC_8_18_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_1_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_1_LC_8_18_4 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \uart_frame_decoder.count_1_LC_8_18_4  (
            .in0(N__14254),
            .in1(N__14697),
            .in2(_gnd_net_),
            .in3(N__16635),
            .lcout(\uart_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25240),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_8_18_5 .C_ON=1'b0;
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_8_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__14269),
            .in2(_gnd_net_),
            .in3(N__14281),
            .lcout(\scaler_1.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.N_508_i_l_ofx_LC_8_18_6 .C_ON=1'b0;
    defparam \scaler_1.N_508_i_l_ofx_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \scaler_1.N_508_i_l_ofx_LC_8_18_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \scaler_1.N_508_i_l_ofx_LC_8_18_6  (
            .in0(N__14282),
            .in1(_gnd_net_),
            .in2(N__14273),
            .in3(_gnd_net_),
            .lcout(\scaler_1.N_508_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_2_LC_8_18_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_2_LC_8_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_2_LC_8_18_7 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \uart_frame_decoder.count_2_LC_8_18_7  (
            .in0(N__16636),
            .in1(N__14255),
            .in2(N__14704),
            .in3(N__14725),
            .lcout(\uart_frame_decoder.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25240),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_0_c_LC_8_19_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_8_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__16694),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\uart_frame_decoder.count8_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_8_19_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_8_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_1_c_inv_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__14243),
            .in2(_gnd_net_),
            .in3(N__14693),
            .lcout(\uart_frame_decoder.count8_axb_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_0 ),
            .carryout(\uart_frame_decoder.count8_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_8_19_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_8_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_inv_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__14237),
            .in2(N__21848),
            .in3(N__14721),
            .lcout(\uart_frame_decoder.count_i_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_1 ),
            .carryout(\uart_frame_decoder.count8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_8_19_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_8_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.count8_THRU_LUT4_0_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14315),
            .lcout(\uart_frame_decoder.count8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_4_LC_8_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_4_LC_8_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_4_LC_8_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_4_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15020),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.elevator_esr_4_LC_8_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_4_LC_8_20_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_4_LC_8_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_4_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14999),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_20_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_8_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16226),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_20_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_4_LC_8_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_4_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15104),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_5_LC_8_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_5_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15116),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_20_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_5_LC_8_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_5_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15128),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25229),
            .ce(N__21707),
            .sr(N__24775));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_8_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_8_21_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_8_21_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_8_21_0  (
            .in0(N__23628),
            .in1(N__23166),
            .in2(N__14396),
            .in3(N__24215),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25225),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_8_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_8_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_8_21_3 .LUT_INIT=16'b1111000111111010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_8_21_3  (
            .in0(N__22240),
            .in1(N__22751),
            .in2(N__24930),
            .in3(N__23630),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25225),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI5DVT_2_LC_8_21_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI5DVT_2_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI5DVT_2_LC_8_21_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.state_1_RNI5DVT_2_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(N__21361),
            .in2(_gnd_net_),
            .in3(N__24912),
            .lcout(\uart_frame_decoder.source_CH1data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_8_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_8_21_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_8_21_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_8_21_6  (
            .in0(N__23629),
            .in1(N__24916),
            .in2(N__26090),
            .in3(N__15476),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25225),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_8_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_8_21_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_8_21_7  (
            .in0(N__22024),
            .in1(N__22750),
            .in2(_gnd_net_),
            .in3(N__23627),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_8_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_8_22_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14369),
            .in3(N__14348),
            .lcout(\ppm_encoder_1.N_230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_22_1 .LUT_INIT=16'b1111000111111010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_22_1  (
            .in0(N__15457),
            .in1(N__22694),
            .in2(N__24931),
            .in3(N__23556),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25220),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_8_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_8_22_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_8_22_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_8_22_2  (
            .in0(N__23554),
            .in1(N__24214),
            .in2(N__14395),
            .in3(N__14350),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25220),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_8_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_8_22_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_8_22_3 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_8_22_3  (
            .in0(N__14368),
            .in1(N__14378),
            .in2(N__24932),
            .in3(N__23555),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25220),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_8_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_8_22_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_8_22_4  (
            .in0(N__14367),
            .in1(N__14349),
            .in2(N__15458),
            .in3(N__15474),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_8_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_8_22_5 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_8_22_5  (
            .in0(N__18517),
            .in1(N__23553),
            .in2(N__14333),
            .in3(N__18440),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_8_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_8_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_8_22_6 .LUT_INIT=16'b1010111100001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIALN65_1_LC_8_22_6  (
            .in0(N__19995),
            .in1(N__15518),
            .in2(N__14330),
            .in3(N__18644),
            .lcout(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_8_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_8_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_8_22_7  (
            .in0(N__15437),
            .in1(N__15392),
            .in2(_gnd_net_),
            .in3(N__15624),
            .lcout(\ppm_encoder_1.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_8_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_8_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_8_23_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_8_23_0  (
            .in0(N__22242),
            .in1(N__25932),
            .in2(N__15625),
            .in3(N__23995),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_8_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_8_23_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_8_23_2 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_8_23_2  (
            .in0(N__19473),
            .in1(N__19701),
            .in2(N__14426),
            .in3(N__15491),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25215),
            .ce(),
            .sr(N__24788));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_8_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_8_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_8_23_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_8_23_3  (
            .in0(N__22687),
            .in1(N__23079),
            .in2(_gnd_net_),
            .in3(N__23572),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_8_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_8_23_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_8_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21468),
            .in3(N__23994),
            .lcout(\ppm_encoder_1.PPM_STATE_62_d ),
            .ltout(\ppm_encoder_1.PPM_STATE_62_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_8_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_8_23_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_8_23_5  (
            .in0(N__22241),
            .in1(N__25930),
            .in2(N__14414),
            .in3(N__15617),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_8_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_8_23_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_8_23_6 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_8_23_6  (
            .in0(N__24257),
            .in1(N__21467),
            .in2(N__24027),
            .in3(N__24280),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25215),
            .ce(),
            .sr(N__24788));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_8_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_8_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_8_23_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_8_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24284),
            .in3(N__24019),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25215),
            .ce(),
            .sr(N__24788));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_24_0 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_8_24_0  (
            .in0(N__20026),
            .in1(N__16127),
            .in2(N__23676),
            .in3(N__14513),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_8_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_8_24_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_8_24_1 .LUT_INIT=16'b0001000000110010;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_8_24_1  (
            .in0(N__19497),
            .in1(N__19694),
            .in2(N__14411),
            .in3(N__15530),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25209),
            .ce(),
            .sr(N__24794));
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_8_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_8_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_8_24_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_8_24_2  (
            .in0(N__20025),
            .in1(N__14514),
            .in2(N__23677),
            .in3(N__16125),
            .lcout(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_8_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_8_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_8_24_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_8_24_3  (
            .in0(N__23683),
            .in1(_gnd_net_),
            .in2(N__22752),
            .in3(N__20024),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_8_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_8_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_8_24_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_8_24_4  (
            .in0(N__22138),
            .in1(N__14515),
            .in2(N__23678),
            .in3(N__16126),
            .lcout(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_8_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_8_24_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_8_24_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_8_24_5  (
            .in0(N__19496),
            .in1(N__14474),
            .in2(N__15782),
            .in3(N__19695),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25209),
            .ce(),
            .sr(N__24794));
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_8_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_8_24_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIANUS_2_LC_8_24_6  (
            .in0(N__22137),
            .in1(N__22683),
            .in2(_gnd_net_),
            .in3(N__23682),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_8_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_8_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_8_24_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5V123_2_LC_8_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14465),
            .in3(N__14462),
            .lcout(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_11_LC_8_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_8_25_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_8_25_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_8_25_0  (
            .in0(N__19692),
            .in1(N__14456),
            .in2(N__19551),
            .in3(N__15890),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25204),
            .ce(),
            .sr(N__24798));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_8_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_8_25_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_8_25_1  (
            .in0(N__22548),
            .in1(N__23686),
            .in2(_gnd_net_),
            .in3(N__22787),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_8_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_8_25_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_8_25_2  (
            .in0(N__23684),
            .in1(_gnd_net_),
            .in2(N__22823),
            .in3(N__22549),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_12_LC_8_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_8_25_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_8_25_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_8_25_3  (
            .in0(N__19550),
            .in1(N__14435),
            .in2(N__19706),
            .in3(N__15881),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25204),
            .ce(),
            .sr(N__24798));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_8_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_8_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_8_25_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_12_LC_8_25_4  (
            .in0(N__23687),
            .in1(_gnd_net_),
            .in2(N__22824),
            .in3(N__22458),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_8_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_8_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_8_25_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_8_25_5  (
            .in0(N__22459),
            .in1(N__23685),
            .in2(_gnd_net_),
            .in3(N__22786),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_8_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_8_25_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_8_25_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_8_25_6  (
            .in0(N__19693),
            .in1(N__14567),
            .in2(N__19552),
            .in3(N__15857),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25204),
            .ce(),
            .sr(N__24798));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_8_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_8_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_8_25_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_14_LC_8_25_7  (
            .in0(N__22317),
            .in1(N__23688),
            .in2(_gnd_net_),
            .in3(N__22791),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_8_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_8_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_8_26_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_8_26_0  (
            .in0(N__23692),
            .in1(N__16050),
            .in2(N__22826),
            .in3(N__16146),
            .lcout(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_8_26_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_8_26_1  (
            .in0(N__19576),
            .in1(N__14558),
            .in2(N__19702),
            .in3(N__15833),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25200),
            .ce(),
            .sr(N__24801));
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_8_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_8_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_8_26_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_8_26_2  (
            .in0(N__23690),
            .in1(_gnd_net_),
            .in2(N__22825),
            .in3(N__16051),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_8_26_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_8_26_4  (
            .in0(N__19670),
            .in1(N__14546),
            .in2(N__19583),
            .in3(N__16154),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25200),
            .ce(),
            .sr(N__24801));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_8_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_8_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_8_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_8_26_5  (
            .in0(_gnd_net_),
            .in1(N__22796),
            .in2(_gnd_net_),
            .in3(N__23691),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_8_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_26_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_8_26_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_8_26_6  (
            .in0(N__19669),
            .in1(N__19575),
            .in2(N__14663),
            .in3(N__15932),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25200),
            .ce(),
            .sr(N__24801));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_8_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_8_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_8_26_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_8_26_7  (
            .in0(N__22017),
            .in1(N__22792),
            .in2(_gnd_net_),
            .in3(N__23689),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_8_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_8_27_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_8_27_0 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_8_27_0  (
            .in0(N__19561),
            .in1(N__19667),
            .in2(N__14654),
            .in3(N__15824),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25196),
            .ce(),
            .sr(N__24804));
    defparam \ppm_encoder_1.init_pulses_17_LC_8_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_27_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_8_27_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_8_27_2  (
            .in0(N__19562),
            .in1(N__19668),
            .in2(N__15809),
            .in3(N__14645),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25196),
            .ce(),
            .sr(N__24804));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_8_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_8_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_8_27_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_8_27_3  (
            .in0(N__23681),
            .in1(_gnd_net_),
            .in2(N__22821),
            .in3(N__16071),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_8_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_8_27_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_8_27_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_8_27_5  (
            .in0(N__19666),
            .in1(N__14639),
            .in2(N__19580),
            .in3(N__15701),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25196),
            .ce(),
            .sr(N__24804));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_8_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_8_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_8_27_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_4_LC_8_27_6  (
            .in0(N__19071),
            .in1(N__22772),
            .in2(_gnd_net_),
            .in3(N__23679),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_8_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_8_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_8_27_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_8_27_7  (
            .in0(N__23680),
            .in1(_gnd_net_),
            .in2(N__22820),
            .in3(N__19072),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_esr_6_LC_9_10_1 .C_ON=1'b0;
    defparam \uart_pc.data_esr_6_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_esr_6_LC_9_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc.data_esr_6_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14627),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25281),
            .ce(N__14602),
            .sr(N__14809));
    defparam \uart_frame_decoder.state_1_0_LC_9_11_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_0_LC_9_11_0 .SEQ_MODE=4'b1001;
    defparam \uart_frame_decoder.state_1_0_LC_9_11_0 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \uart_frame_decoder.state_1_0_LC_9_11_0  (
            .in0(N__14671),
            .in1(N__14786),
            .in2(N__14780),
            .in3(N__23913),
            .lcout(\uart_frame_decoder.state_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25276),
            .ce(),
            .sr(N__24742));
    defparam \uart_frame_decoder.state_1_10_LC_9_11_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_10_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_10_LC_9_11_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \uart_frame_decoder.state_1_10_LC_9_11_3  (
            .in0(N__23914),
            .in1(N__14672),
            .in2(N__14741),
            .in3(N__15318),
            .lcout(\uart_frame_decoder.state_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25276),
            .ce(),
            .sr(N__24742));
    defparam \uart_frame_decoder.state_1_RNIF7PK_9_LC_9_12_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIF7PK_9_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIF7PK_9_LC_9_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIF7PK_9_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__14752),
            .in2(_gnd_net_),
            .in3(N__23821),
            .lcout(\uart_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNICKVT_9_LC_9_12_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNICKVT_9_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNICKVT_9_LC_9_12_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_frame_decoder.state_1_RNICKVT_9_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14732),
            .in3(N__24907),
            .lcout(\uart_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_9_12_3 .C_ON=1'b0;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_9_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_9_12_3  (
            .in0(N__16202),
            .in1(N__15039),
            .in2(_gnd_net_),
            .in3(N__15080),
            .lcout(\scaler_2.un2_source_data_0_cry_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNINMHJ_10_LC_9_12_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNINMHJ_10_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNINMHJ_10_LC_9_12_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uart_frame_decoder.state_1_RNINMHJ_10_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__23820),
            .in2(_gnd_net_),
            .in3(N__15315),
            .lcout(\uart_frame_decoder.state_1_RNINMHJZ0Z_10 ),
            .ltout(\uart_frame_decoder.state_1_RNINMHJZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_RNI8GDP1_2_LC_9_12_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNI8GDP1_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNI8GDP1_2_LC_9_12_5 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \uart_frame_decoder.count_RNI8GDP1_2_LC_9_12_5  (
            .in0(N__14729),
            .in1(N__14705),
            .in2(N__14675),
            .in3(N__16622),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_o2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_9_13_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_0_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21094),
            .lcout(frame_decoder_CH2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_9_13_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_1_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20976),
            .lcout(frame_decoder_CH2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_9_13_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_2_LC_9_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20892),
            .lcout(frame_decoder_CH2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_9_13_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_3_LC_9_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_3_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20809),
            .lcout(frame_decoder_CH2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_9_13_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_4_LC_9_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20720),
            .lcout(frame_decoder_CH2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_9_13_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_5_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26355),
            .lcout(frame_decoder_CH2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_9_13_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_6_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20606),
            .lcout(frame_decoder_CH2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25267),
            .ce(N__17815),
            .sr(N__24748));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_9_14_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__15038),
            .in2(N__15085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_9_14_1 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__14864),
            .in2(N__14858),
            .in3(N__14849),
            .lcout(\scaler_2.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_0 ),
            .carryout(\scaler_2.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_9_14_2 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__14846),
            .in2(N__14840),
            .in3(N__14831),
            .lcout(\scaler_2.un3_source_data_0_cry_1_c_RNILSPH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_1 ),
            .carryout(\scaler_2.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_9_14_3 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__14828),
            .in2(N__14822),
            .in3(N__14813),
            .lcout(\scaler_2.un3_source_data_0_cry_2_c_RNIO0RH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_2 ),
            .carryout(\scaler_2.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_9_14_4 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_9_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__14960),
            .in2(N__14954),
            .in3(N__14945),
            .lcout(\scaler_2.un3_source_data_0_cry_3_c_RNIR4SH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_3 ),
            .carryout(\scaler_2.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_9_14_5 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_9_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__14942),
            .in2(N__14936),
            .in3(N__14927),
            .lcout(\scaler_2.un3_source_data_0_cry_4_c_RNIU8TH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_4 ),
            .carryout(\scaler_2.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_9_14_6 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_9_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__14924),
            .in2(N__14918),
            .in3(N__14909),
            .lcout(\scaler_2.un3_source_data_0_cry_5_c_RNI1DUH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_5 ),
            .carryout(\scaler_2.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_9_14_7 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__17846),
            .in2(_gnd_net_),
            .in3(N__14906),
            .lcout(\scaler_2.un3_source_data_0_cry_6_c_RNI4HVH ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_6 ),
            .carryout(\scaler_2.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_9_15_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__15134),
            .in2(N__21916),
            .in3(N__14903),
            .lcout(\scaler_2.un3_source_data_0_cry_7_c_RNI5J0I ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_9_15_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_9_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14900),
            .lcout(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI91PK_3_LC_9_15_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI91PK_3_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI91PK_3_LC_9_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNI91PK_3_LC_9_15_2  (
            .in0(N__23792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14897),
            .lcout(\uart_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(\uart_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI6EVT_3_LC_9_15_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI6EVT_3_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI6EVT_3_LC_9_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_frame_decoder.state_1_RNI6EVT_3_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14867),
            .in3(N__24908),
            .lcout(\uart_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_9_15_6 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_9_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__16669),
            .in2(_gnd_net_),
            .in3(N__21379),
            .lcout(\scaler_3.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.N_520_i_l_ofx_LC_9_15_7 .C_ON=1'b0;
    defparam \scaler_2.N_520_i_l_ofx_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.N_520_i_l_ofx_LC_9_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_2.N_520_i_l_ofx_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__17860),
            .in2(_gnd_net_),
            .in3(N__17837),
            .lcout(\scaler_2.N_520_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.source_data_1_esr_5_LC_9_16_0 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_5_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_5_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_1.source_data_1_esr_5_LC_9_16_0  (
            .in0(N__16502),
            .in1(N__16592),
            .in2(_gnd_net_),
            .in3(N__16555),
            .lcout(scaler_1_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25246),
            .ce(N__21142),
            .sr(N__24760));
    defparam \scaler_2.source_data_1_esr_5_LC_9_16_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_5_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_5_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.source_data_1_esr_5_LC_9_16_1  (
            .in0(N__16201),
            .in1(N__15081),
            .in2(_gnd_net_),
            .in3(N__15047),
            .lcout(scaler_2_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25246),
            .ce(N__21142),
            .sr(N__24760));
    defparam \scaler_3.source_data_1_esr_5_LC_9_16_2 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_5_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_5_LC_9_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.source_data_1_esr_5_LC_9_16_2  (
            .in0(N__21026),
            .in1(N__18069),
            .in2(_gnd_net_),
            .in3(N__16451),
            .lcout(scaler_3_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25246),
            .ce(N__21142),
            .sr(N__24760));
    defparam \scaler_1.source_data_1_4_LC_9_17_1 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_4_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_4_LC_9_17_1 .LUT_INIT=16'b0101110010101100;
    LogicCell40 \scaler_1.source_data_1_4_LC_9_17_1  (
            .in0(N__16587),
            .in1(N__15097),
            .in2(N__20176),
            .in3(N__16556),
            .lcout(scaler_1_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25241),
            .ce(),
            .sr(N__24766));
    defparam \scaler_2.source_data_1_4_LC_9_17_3 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_4_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_4_LC_9_17_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_2.source_data_1_4_LC_9_17_3  (
            .in0(N__20167),
            .in1(N__15086),
            .in2(N__15016),
            .in3(N__15046),
            .lcout(scaler_2_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25241),
            .ce(),
            .sr(N__24766));
    defparam \scaler_3.source_data_1_4_LC_9_17_5 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_4_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_4_LC_9_17_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \scaler_3.source_data_1_4_LC_9_17_5  (
            .in0(N__20168),
            .in1(N__21025),
            .in2(N__16460),
            .in3(N__14998),
            .lcout(scaler_3_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25241),
            .ce(),
            .sr(N__24766));
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_9_17_6 .C_ON=1'b0;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_9_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_9_17_6  (
            .in0(N__18074),
            .in1(N__16455),
            .in2(_gnd_net_),
            .in3(N__21018),
            .lcout(\scaler_3.un2_source_data_0_cry_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_4_LC_9_17_7 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_9_17_7 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_9_17_7  (
            .in0(N__20169),
            .in1(N__17900),
            .in2(N__14977),
            .in3(N__17936),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25241),
            .ce(),
            .sr(N__24766));
    defparam \ppm_encoder_1.rudder_10_LC_9_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_9_18_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_9_18_1  (
            .in0(N__20279),
            .in1(N__18110),
            .in2(N__25494),
            .in3(N__22042),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25233),
            .ce(),
            .sr(N__24771));
    defparam \scaler_1.source_data_valid_LC_9_18_3 .C_ON=1'b0;
    defparam \scaler_1.source_data_valid_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_valid_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_1.source_data_valid_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20165),
            .lcout(scaler_1_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25233),
            .ce(),
            .sr(N__24771));
    defparam \uart_frame_decoder.source_data_valid_LC_9_18_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_data_valid_LC_9_18_5 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \uart_frame_decoder.source_data_valid_LC_9_18_5  (
            .in0(N__15281),
            .in1(N__15329),
            .in2(N__23787),
            .in3(N__20166),
            .lcout(pc_frame_decoder_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25233),
            .ce(),
            .sr(N__24771));
    defparam \uart_frame_decoder.count8_cry_2_c_RNIU1C61_LC_9_18_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_2_c_RNIU1C61_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_RNIU1C61_LC_9_18_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_RNIU1C61_LC_9_18_6  (
            .in0(N__15328),
            .in1(N__24177),
            .in2(N__23818),
            .in3(N__15280),
            .lcout(\uart_frame_decoder.count8_cry_2_c_RNIU1CZ0Z61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_rdy_LC_9_18_7 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_9_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__15268),
            .in2(_gnd_net_),
            .in3(N__15165),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25233),
            .ce(),
            .sr(N__24771));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_9_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_9_19_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_9_19_0  (
            .in0(N__16960),
            .in1(N__25777),
            .in2(_gnd_net_),
            .in3(N__16982),
            .lcout(\ppm_encoder_1.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_19_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_19_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_9_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_9_19_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(_gnd_net_),
            .in3(N__24911),
            .lcout(\ppm_encoder_1.scaler_1_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_9_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_9_20_1 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNIG4JI2_11_LC_9_20_1  (
            .in0(N__16917),
            .in1(N__22531),
            .in2(N__18689),
            .in3(N__18769),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_9_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_9_20_2 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIALRT5_11_LC_9_20_2  (
            .in0(N__15923),
            .in1(_gnd_net_),
            .in2(N__15137),
            .in3(N__15362),
            .lcout(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_9_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_9_20_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI03DH2_11_LC_9_20_3  (
            .in0(N__16936),
            .in1(N__15351),
            .in2(N__18543),
            .in3(N__18452),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_9_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_9_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_9_20_4  (
            .in0(N__25787),
            .in1(N__16918),
            .in2(_gnd_net_),
            .in3(N__16937),
            .lcout(),
            .ltout(\ppm_encoder_1.N_306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_9_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_9_20_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__26101),
            .in2(N__15356),
            .in3(N__15352),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_9_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_9_20_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_9_20_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_9_20_6  (
            .in0(N__15353),
            .in1(N__25473),
            .in2(N__19217),
            .in3(N__19190),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25226),
            .ce(),
            .sr(N__24778));
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_9_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_9_21_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.throttle_RNIS5KK2_8_LC_9_21_0  (
            .in0(N__21640),
            .in1(N__18746),
            .in2(N__19037),
            .in3(N__18674),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_9_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_9_21_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIONI96_8_LC_9_21_1  (
            .in0(N__17423),
            .in1(_gnd_net_),
            .in2(N__15341),
            .in3(N__15338),
            .lcout(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_9_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_9_21_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNICKVN2_8_LC_9_21_2  (
            .in0(N__16849),
            .in1(N__16876),
            .in2(N__18451),
            .in3(N__18513),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_9_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_9_21_3 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \ppm_encoder_1.throttle_RNIU7KK2_9_LC_9_21_3  (
            .in0(N__18673),
            .in1(N__19133),
            .in2(N__18768),
            .in3(N__25633),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_9_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_9_21_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNITSI96_9_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__17372),
            .in2(N__15332),
            .in3(N__15482),
            .lcout(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_9_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_9_21_5 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \ppm_encoder_1.elevator_RNIEMVN2_9_LC_9_21_5  (
            .in0(N__18512),
            .in1(N__16903),
            .in2(N__25656),
            .in3(N__18435),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_9_LC_9_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_9_21_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_9_21_7  (
            .in0(N__18251),
            .in1(N__18275),
            .in2(N__25528),
            .in3(N__25658),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25221),
            .ce(),
            .sr(N__24783));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_9_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_9_22_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_9_22_0  (
            .in0(N__15475),
            .in1(N__15456),
            .in2(N__23590),
            .in3(N__25929),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_9_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_9_22_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_9_22_1  (
            .in0(N__15436),
            .in1(N__15422),
            .in2(N__15407),
            .in3(N__18429),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_9_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_9_22_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_9_22_2 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_9_22_2  (
            .in0(N__15616),
            .in1(N__24927),
            .in2(N__26100),
            .in3(N__23588),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25216),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_9_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_9_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__23503),
            .in2(_gnd_net_),
            .in3(N__15403),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI62ME2_4_LC_9_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI62ME2_4_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI62ME2_4_LC_9_22_4 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI62ME2_4_LC_9_22_4  (
            .in0(N__15391),
            .in1(N__19054),
            .in2(N__15374),
            .in3(N__18643),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI8CGI5_4_LC_9_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI8CGI5_4_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI8CGI5_4_LC_9_22_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI8CGI5_4_LC_9_22_5  (
            .in0(N__15737),
            .in1(_gnd_net_),
            .in2(N__15371),
            .in3(N__15368),
            .lcout(\ppm_encoder_1.aileron_esr_RNI8CGI5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_9_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_9_22_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_9_22_6  (
            .in0(N__23504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.N_614_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_9_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_9_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_9_22_7  (
            .in0(N__22233),
            .in1(N__15615),
            .in2(N__25936),
            .in3(N__23499),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI84ME2_5_LC_9_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI84ME2_5_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI84ME2_5_LC_9_23_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI84ME2_5_LC_9_23_0  (
            .in0(N__15568),
            .in1(N__22081),
            .in2(N__18766),
            .in3(N__18656),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIDHGI5_5_LC_9_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIDHGI5_5_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIDHGI5_5_LC_9_23_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIDHGI5_5_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__18916),
            .in2(N__15590),
            .in3(N__15587),
            .lcout(\ppm_encoder_1.aileron_esr_RNIDHGI5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_9_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_9_23_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_9_23_2  (
            .in0(N__15580),
            .in1(N__18505),
            .in2(N__15545),
            .in3(N__18431),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_9_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_9_23_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_9_23_3  (
            .in0(N__25805),
            .in1(N__15581),
            .in2(_gnd_net_),
            .in3(N__15569),
            .lcout(),
            .ltout(\ppm_encoder_1.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_9_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_9_23_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_9_23_4  (
            .in0(N__26062),
            .in1(_gnd_net_),
            .in2(N__15557),
            .in3(N__15544),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_5_LC_9_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_5_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_5_LC_9_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_5_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15554),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25210),
            .ce(N__21731),
            .sr(N__24795));
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_0_LC_9_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_0_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_0_LC_9_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8LUS_0_0_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__15529),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__15514),
            .in2(N__15503),
            .in3(N__15485),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__15797),
            .in2(N__15791),
            .in3(N__15770),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__15767),
            .in2(N__15752),
            .in3(N__15740),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__15736),
            .in2(N__15713),
            .in3(N__15689),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__18917),
            .in2(N__15686),
            .in3(N__15677),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__17083),
            .in2(N__17057),
            .in3(N__15662),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__17162),
            .in2(N__17188),
            .in3(N__15659),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_25_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__17419),
            .in2(N__15656),
            .in3(N__15644),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_25_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__17365),
            .in2(N__15641),
            .in3(N__15629),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_25_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__17221),
            .in2(N__17204),
            .in3(N__15926),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_25_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__15919),
            .in2(N__15902),
            .in3(N__15884),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_25_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__17038),
            .in2(N__17024),
            .in3(N__15875),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_25_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__17314),
            .in2(N__17297),
            .in3(N__15860),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_25_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__18577),
            .in2(N__18563),
            .in3(N__15851),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_25_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__15848),
            .in2(N__15842),
            .in3(N__15827),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_26_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__15941),
            .in2(_gnd_net_),
            .in3(N__15818),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_26_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__15815),
            .in2(_gnd_net_),
            .in3(N__15800),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__16094),
            .in2(_gnd_net_),
            .in3(N__16157),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_9_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_9_26_5 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_9_26_5  (
            .in0(N__22813),
            .in1(N__16148),
            .in2(N__15978),
            .in3(N__23675),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_9_26_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_9_26_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_9_26_7  (
            .in0(N__22910),
            .in1(N__26192),
            .in2(N__16037),
            .in3(N__22886),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_9_27_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_9_27_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__16088),
            .in2(_gnd_net_),
            .in3(N__24239),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_16_LC_9_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_9_28_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_9_28_1  (
            .in0(N__15955),
            .in1(N__17564),
            .in2(N__16019),
            .in3(N__23712),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25190),
            .ce(),
            .sr(N__24808));
    defparam \ppm_encoder_1.pulses2count_17_LC_9_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_9_28_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_9_28_2  (
            .in0(N__23709),
            .in1(N__16016),
            .in2(N__16076),
            .in3(N__17551),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25190),
            .ce(),
            .sr(N__24808));
    defparam \ppm_encoder_1.pulses2count_15_LC_9_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_9_28_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_9_28_3  (
            .in0(N__16055),
            .in1(N__16033),
            .in2(N__16018),
            .in3(N__23711),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25190),
            .ce(),
            .sr(N__24808));
    defparam \ppm_encoder_1.pulses2count_18_LC_9_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_9_28_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_9_28_4  (
            .in0(N__23710),
            .in1(N__16017),
            .in2(N__15986),
            .in3(N__17531),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25190),
            .ce(),
            .sr(N__24808));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_9_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_9_28_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_9_28_7  (
            .in0(N__15954),
            .in1(N__22837),
            .in2(_gnd_net_),
            .in3(N__23708),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_10_12_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_0_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21107),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_1_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_1_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20980),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_10_12_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_7_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_7_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20535),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_3_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_3_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20810),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_5_LC_10_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_5_LC_10_12_5  (
            .in0(N__26363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_10_12_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_6_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_6_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20613),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_10_12_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_2_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_2_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20893),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25260),
            .ce(N__20119),
            .sr(N__24744));
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_10_13_0 .C_ON=1'b1;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__16190),
            .in2(N__16211),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_6_LC_10_13_1 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_6_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_6_LC_10_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_6_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__16165),
            .in2(N__16200),
            .in3(N__16172),
            .lcout(scaler_2_data_6),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_1 ),
            .carryout(\scaler_2.un2_source_data_0_cry_2 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_7_LC_10_13_2 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_7_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_7_LC_10_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_7_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__16327),
            .in2(N__16169),
            .in3(N__16334),
            .lcout(scaler_2_data_7),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_2 ),
            .carryout(\scaler_2.un2_source_data_0_cry_3 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_8_LC_10_13_3 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_8_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_8_LC_10_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_8_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__16312),
            .in2(N__16331),
            .in3(N__16319),
            .lcout(scaler_2_data_8),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_3 ),
            .carryout(\scaler_2.un2_source_data_0_cry_4 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_9_LC_10_13_4 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_9_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_9_LC_10_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_9_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__16297),
            .in2(N__16316),
            .in3(N__16304),
            .lcout(scaler_2_data_9),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_4 ),
            .carryout(\scaler_2.un2_source_data_0_cry_5 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_10_LC_10_13_5 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_10_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_10_LC_10_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_10_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__16282),
            .in2(N__16301),
            .in3(N__16289),
            .lcout(scaler_2_data_10),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_5 ),
            .carryout(\scaler_2.un2_source_data_0_cry_6 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_11_LC_10_13_6 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_11_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_11_LC_10_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_11_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__16267),
            .in2(N__16286),
            .in3(N__16274),
            .lcout(scaler_2_data_11),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_6 ),
            .carryout(\scaler_2.un2_source_data_0_cry_7 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_12_LC_10_13_7 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_12_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_12_LC_10_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_12_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__16256),
            .in2(N__16271),
            .in3(N__16259),
            .lcout(scaler_2_data_12),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_7 ),
            .carryout(\scaler_2.un2_source_data_0_cry_8 ),
            .clk(N__25253),
            .ce(N__21137),
            .sr(N__24749));
    defparam \scaler_2.source_data_1_esr_13_LC_10_14_0 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_13_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_13_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_13_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__16255),
            .in2(N__16241),
            .in3(N__16232),
            .lcout(scaler_2_data_13),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_9 ),
            .clk(N__25248),
            .ce(N__21138),
            .sr(N__24753));
    defparam \scaler_2.source_data_1_esr_14_LC_10_14_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_14_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_14_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_2.source_data_1_esr_14_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16229),
            .lcout(scaler_2_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25248),
            .ce(N__21138),
            .sr(N__24753));
    defparam \scaler_4.source_data_1_esr_5_LC_10_14_4 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_10_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_10_14_4  (
            .in0(N__20441),
            .in1(N__17896),
            .in2(_gnd_net_),
            .in3(N__17935),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25248),
            .ce(N__21138),
            .sr(N__24753));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_10_15_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_10_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__21017),
            .in2(N__16459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_10_15_1 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__20909),
            .in2(N__16427),
            .in3(N__16415),
            .lcout(\scaler_3.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_0 ),
            .carryout(\scaler_3.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_10_15_2 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__20822),
            .in2(N__16412),
            .in3(N__16400),
            .lcout(\scaler_3.un3_source_data_0_cry_1_c_RNIOS6I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_1 ),
            .carryout(\scaler_3.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_10_15_3 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(N__20741),
            .in3(N__16388),
            .lcout(\scaler_3.un3_source_data_0_cry_2_c_RNIR08I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_2 ),
            .carryout(\scaler_3.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_10_15_4 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__16385),
            .in2(N__20645),
            .in3(N__16376),
            .lcout(\scaler_3.un3_source_data_0_cry_3_c_RNIU49I ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_3 ),
            .carryout(\scaler_3.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_10_15_5 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__26279),
            .in2(N__16373),
            .in3(N__16358),
            .lcout(\scaler_3.un3_source_data_0_cry_4_c_RNI19AI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_4 ),
            .carryout(\scaler_3.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_10_15_6 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__16355),
            .in2(N__20549),
            .in3(N__16346),
            .lcout(\scaler_3.un3_source_data_0_cry_5_c_RNI4DBI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_5 ),
            .carryout(\scaler_3.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_10_15_7 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_10_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__16343),
            .in2(_gnd_net_),
            .in3(N__16337),
            .lcout(\scaler_3.un3_source_data_0_cry_6_c_RNI7HCI ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_6 ),
            .carryout(\scaler_3.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_10_16_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__16658),
            .in2(N__21922),
            .in3(N__16700),
            .lcout(\scaler_3.un3_source_data_0_cry_7_c_RNI8JDI ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_10_16_1 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_10_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16697),
            .lcout(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_10_16_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_10_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_inv_LC_10_16_2  (
            .in0(N__21893),
            .in1(N__16690),
            .in2(_gnd_net_),
            .in3(N__16610),
            .lcout(\uart_frame_decoder.count8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.N_532_i_l_ofx_LC_10_16_3 .C_ON=1'b0;
    defparam \scaler_3.N_532_i_l_ofx_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.N_532_i_l_ofx_LC_10_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_3.N_532_i_l_ofx_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__16676),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(\scaler_3.N_532_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_0_LC_10_16_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_0_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_0_LC_10_16_5 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \uart_frame_decoder.count_0_LC_10_16_5  (
            .in0(N__16611),
            .in1(N__16652),
            .in2(_gnd_net_),
            .in3(N__16640),
            .lcout(\uart_frame_decoder.count8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25235),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_10_16_7 .C_ON=1'b0;
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_10_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_10_16_7  (
            .in0(N__16511),
            .in1(N__16591),
            .in2(_gnd_net_),
            .in3(N__16554),
            .lcout(\scaler_1.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_10_17_0 .C_ON=1'b1;
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \scaler_1.un2_source_data_0_cry_1_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_1.un2_source_data_0_cry_1_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__16503),
            .in2(N__16520),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\scaler_1.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_1.source_data_1_esr_6_LC_10_17_1 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_6_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_6_LC_10_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_6_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__16474),
            .in2(N__16510),
            .in3(N__16481),
            .lcout(scaler_1_data_6),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_1 ),
            .carryout(\scaler_1.un2_source_data_0_cry_2 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_7_LC_10_17_2 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_7_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_7_LC_10_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_7_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__16822),
            .in2(N__16478),
            .in3(N__16463),
            .lcout(scaler_1_data_7),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_2 ),
            .carryout(\scaler_1.un2_source_data_0_cry_3 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_8_LC_10_17_3 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_8_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_8_LC_10_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_8_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__16804),
            .in2(N__16826),
            .in3(N__16811),
            .lcout(scaler_1_data_8),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_3 ),
            .carryout(\scaler_1.un2_source_data_0_cry_4 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_9_LC_10_17_4 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_9_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_9_LC_10_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_9_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__16786),
            .in2(N__16808),
            .in3(N__16793),
            .lcout(scaler_1_data_9),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_4 ),
            .carryout(\scaler_1.un2_source_data_0_cry_5 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_10_LC_10_17_5 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_10_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_10_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_10_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__16768),
            .in2(N__16790),
            .in3(N__16775),
            .lcout(scaler_1_data_10),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_5 ),
            .carryout(\scaler_1.un2_source_data_0_cry_6 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_11_LC_10_17_6 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_11_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_11_LC_10_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_11_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__16750),
            .in2(N__16772),
            .in3(N__16757),
            .lcout(scaler_1_data_11),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_6 ),
            .carryout(\scaler_1.un2_source_data_0_cry_7 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_12_LC_10_17_7 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_12_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_12_LC_10_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_12_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__16735),
            .in2(N__16754),
            .in3(N__16739),
            .lcout(scaler_1_data_12),
            .ltout(),
            .carryin(\scaler_1.un2_source_data_0_cry_7 ),
            .carryout(\scaler_1.un2_source_data_0_cry_8 ),
            .clk(N__25231),
            .ce(N__21141),
            .sr(N__24767));
    defparam \scaler_1.source_data_1_esr_13_LC_10_18_0 .C_ON=1'b1;
    defparam \scaler_1.source_data_1_esr_13_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_13_LC_10_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_1.source_data_1_esr_13_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__16736),
            .in2(N__16718),
            .in3(N__16706),
            .lcout(scaler_1_data_13),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\scaler_1.un2_source_data_0_cry_9 ),
            .clk(N__25227),
            .ce(N__21143),
            .sr(N__24772));
    defparam \scaler_1.source_data_1_esr_14_LC_10_18_1 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_14_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \scaler_1.source_data_1_esr_14_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_1.source_data_1_esr_14_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16703),
            .lcout(scaler_1_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25227),
            .ce(N__21143),
            .sr(N__24772));
    defparam \ppm_encoder_1.aileron_8_LC_10_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_10_19_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_10_19_0  (
            .in0(N__19325),
            .in1(N__19304),
            .in2(N__16850),
            .in3(N__25424),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.rudder_8_LC_10_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_10_19_1 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_10_19_1  (
            .in0(N__25430),
            .in1(N__20351),
            .in2(N__19032),
            .in3(N__18125),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.aileron_9_LC_10_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_10_19_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_10_19_2  (
            .in0(N__19285),
            .in1(N__19265),
            .in2(N__16904),
            .in3(N__25425),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.elevator_11_LC_10_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_10_19_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_10_19_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_10_19_3  (
            .in0(N__18197),
            .in1(N__18176),
            .in2(N__25495),
            .in3(N__16935),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.elevator_8_LC_10_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_10_19_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_10_19_4  (
            .in0(N__18284),
            .in1(N__18302),
            .in2(N__16877),
            .in3(N__25429),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.throttle_11_LC_10_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_10_19_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_10_19_5  (
            .in0(N__21275),
            .in1(N__21257),
            .in2(N__25496),
            .in3(N__16919),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.throttle_7_LC_10_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_10_19_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_10_19_6  (
            .in0(N__21299),
            .in1(N__21317),
            .in2(N__17147),
            .in3(N__25434),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25222),
            .ce(),
            .sr(N__24776));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_10_20_1  (
            .in0(N__26099),
            .in1(N__25610),
            .in2(_gnd_net_),
            .in3(N__16899),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_10_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_10_20_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__25897),
            .in2(N__16880),
            .in3(N__19112),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25218),
            .ce(N__26175),
            .sr(N__24779));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_3  (
            .in0(N__25794),
            .in1(N__21641),
            .in2(_gnd_net_),
            .in3(N__16872),
            .lcout(),
            .ltout(\ppm_encoder_1.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_4  (
            .in0(N__26092),
            .in1(_gnd_net_),
            .in2(N__16853),
            .in3(N__16845),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_10_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_10_20_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_10_20_5  (
            .in0(N__25898),
            .in1(_gnd_net_),
            .in2(N__17048),
            .in3(N__18974),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25218),
            .ce(N__26175),
            .sr(N__24779));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_10_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_10_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_10_20_6  (
            .in0(N__26091),
            .in1(N__17126),
            .in2(_gnd_net_),
            .in3(N__17102),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_10_21_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_10_21_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNII6JI2_12_LC_10_21_0  (
            .in0(N__16953),
            .in1(N__22444),
            .in2(N__18773),
            .in3(N__18690),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_10_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_10_21_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIFQRT5_12_LC_10_21_1  (
            .in0(N__17045),
            .in1(_gnd_net_),
            .in2(N__17027),
            .in3(N__17009),
            .lcout(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_10_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_10_21_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI25DH2_12_LC_10_21_2  (
            .in0(N__16974),
            .in1(N__16992),
            .in2(N__18536),
            .in3(N__18444),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_21_4  (
            .in0(N__26073),
            .in1(N__17003),
            .in2(_gnd_net_),
            .in3(N__16993),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_10_21_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_10_21_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_10_21_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_10_21_5  (
            .in0(N__16994),
            .in1(N__25477),
            .in2(N__19877),
            .in3(N__19850),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25212),
            .ce(),
            .sr(N__24784));
    defparam \ppm_encoder_1.elevator_12_LC_10_21_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_10_21_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_10_21_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_10_21_6  (
            .in0(N__16975),
            .in1(N__18896),
            .in2(N__25529),
            .in3(N__18875),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25212),
            .ce(),
            .sr(N__24784));
    defparam \ppm_encoder_1.throttle_12_LC_10_21_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_10_21_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_10_21_7  (
            .in0(N__21242),
            .in1(N__21218),
            .in2(N__16961),
            .in3(N__25481),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25212),
            .ce(),
            .sr(N__24784));
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_10_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_10_22_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_10_22_0  (
            .in0(N__17145),
            .in1(N__19092),
            .in2(N__18765),
            .in3(N__18687),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_10_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_10_22_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIJII96_7_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__17189),
            .in2(N__17165),
            .in3(N__17153),
            .lcout(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_10_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_10_22_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIAIVN2_7_LC_10_22_2  (
            .in0(N__17115),
            .in1(N__17097),
            .in2(N__18530),
            .in3(N__18430),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_10_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_10_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_10_22_3  (
            .in0(N__25747),
            .in1(N__17146),
            .in2(_gnd_net_),
            .in3(N__17116),
            .lcout(\ppm_encoder_1.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_7_LC_10_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_10_22_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_10_22_4 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_10_22_4  (
            .in0(N__25522),
            .in1(N__17117),
            .in2(N__18320),
            .in3(N__18341),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25206),
            .ce(),
            .sr(N__24789));
    defparam \ppm_encoder_1.aileron_7_LC_10_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_10_22_6 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_10_22_6  (
            .in0(N__25521),
            .in1(N__17098),
            .in2(N__19364),
            .in3(N__19337),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25206),
            .ce(),
            .sr(N__24789));
    defparam \ppm_encoder_1.rudder_7_LC_10_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_10_22_7 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_10_22_7  (
            .in0(N__19093),
            .in1(N__18140),
            .in2(N__20399),
            .in3(N__25523),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25206),
            .ce(),
            .sr(N__24789));
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_10_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_10_23_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIO1KK2_6_LC_10_23_0  (
            .in0(N__17235),
            .in1(N__26233),
            .in2(N__18767),
            .in3(N__18672),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_10_23_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_10_23_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEDI96_6_LC_10_23_1  (
            .in0(N__17084),
            .in1(_gnd_net_),
            .in2(N__17060),
            .in3(N__17255),
            .lcout(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_10_23_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_10_23_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNI8GVN2_6_LC_10_23_2  (
            .in0(N__17247),
            .in1(N__22569),
            .in2(N__18531),
            .in3(N__18436),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_10_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_10_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_10_23_3  (
            .in0(N__25785),
            .in1(N__17236),
            .in2(_gnd_net_),
            .in3(N__17248),
            .lcout(\ppm_encoder_1.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_10_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_10_23_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_10_23_5 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_10_23_5  (
            .in0(N__22570),
            .in1(N__25516),
            .in2(_gnd_net_),
            .in3(N__19396),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25202),
            .ce(),
            .sr(N__24796));
    defparam \ppm_encoder_1.elevator_6_LC_10_23_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_10_23_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_10_23_6 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_10_23_6  (
            .in0(N__17249),
            .in1(_gnd_net_),
            .in2(N__25548),
            .in3(N__18362),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25202),
            .ce(),
            .sr(N__24796));
    defparam \ppm_encoder_1.throttle_6_LC_10_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_10_23_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_10_23_7 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_10_23_7  (
            .in0(N__21335),
            .in1(N__25520),
            .in2(_gnd_net_),
            .in3(N__17237),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25202),
            .ce(),
            .sr(N__24796));
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_10_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_10_24_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIE2JI2_10_LC_10_24_0  (
            .in0(N__21550),
            .in1(N__22054),
            .in2(N__18781),
            .in3(N__18691),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_10_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_10_24_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI5GRT5_10_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__17225),
            .in2(N__17207),
            .in3(N__17195),
            .lcout(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_10_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_10_24_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNIU0DH2_10_LC_10_24_2  (
            .in0(N__17325),
            .in1(N__17337),
            .in2(N__18544),
            .in3(N__18454),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_24_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_24_3  (
            .in0(N__25786),
            .in1(N__21551),
            .in2(_gnd_net_),
            .in3(N__17326),
            .lcout(),
            .ltout(\ppm_encoder_1.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_24_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_24_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__26011),
            .in2(N__17342),
            .in3(N__17338),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_10_LC_10_24_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_10_24_5 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_10_24_5  (
            .in0(N__17339),
            .in1(N__25554),
            .in2(N__19250),
            .in3(N__19226),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25198),
            .ce(),
            .sr(N__24799));
    defparam \ppm_encoder_1.elevator_10_LC_10_24_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_10_24_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_10_24_6  (
            .in0(N__17327),
            .in1(N__18212),
            .in2(N__25559),
            .in3(N__18236),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25198),
            .ce(),
            .sr(N__24799));
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_10_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_10_25_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIK8JI2_13_LC_10_25_0  (
            .in0(N__17265),
            .in1(N__22396),
            .in2(N__18785),
            .in3(N__18692),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_10_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_10_25_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIKVRT5_13_LC_10_25_1  (
            .in0(N__17315),
            .in1(_gnd_net_),
            .in2(N__17300),
            .in3(N__17288),
            .lcout(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_10_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_10_25_2 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNI47DH2_13_LC_10_25_2  (
            .in0(N__25321),
            .in1(N__17277),
            .in2(N__18548),
            .in3(N__18455),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_10_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_10_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_10_25_3  (
            .in0(N__17278),
            .in1(N__25806),
            .in2(_gnd_net_),
            .in3(N__17266),
            .lcout(),
            .ltout(\ppm_encoder_1.N_308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_10_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_10_25_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_10_25_4  (
            .in0(N__25322),
            .in1(_gnd_net_),
            .in2(N__17282),
            .in3(N__26048),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_13_LC_10_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_10_25_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_10_25_6 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_10_25_6  (
            .in0(N__18836),
            .in1(N__25524),
            .in2(N__18863),
            .in3(N__17279),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25194),
            .ce(),
            .sr(N__24802));
    defparam \ppm_encoder_1.throttle_13_LC_10_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_10_25_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_10_25_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_10_25_7  (
            .in0(N__21985),
            .in1(N__21788),
            .in2(N__25549),
            .in3(N__17267),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25194),
            .ce(),
            .sr(N__24802));
    defparam \ppm_encoder_1.init_pulses_8_LC_10_26_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_26_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_26_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_10_26_0  (
            .in0(N__19671),
            .in1(N__17441),
            .in2(N__19581),
            .in3(N__17429),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25192),
            .ce(),
            .sr(N__24805));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_10_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_10_26_1 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_10_26_1  (
            .in0(N__23701),
            .in1(N__18988),
            .in2(N__22838),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_10_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_10_26_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_10_26_2  (
            .in0(N__18987),
            .in1(N__22814),
            .in2(_gnd_net_),
            .in3(N__23699),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_10_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_10_26_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_10_26_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_10_26_4  (
            .in0(N__19672),
            .in1(N__17390),
            .in2(N__19582),
            .in3(N__17378),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25192),
            .ce(),
            .sr(N__24805));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_10_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_10_26_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_10_26_5  (
            .in0(N__22819),
            .in1(_gnd_net_),
            .in2(N__23714),
            .in3(N__19147),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_10_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_10_26_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_10_26_6  (
            .in0(N__19146),
            .in1(N__23700),
            .in2(_gnd_net_),
            .in3(N__22815),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_27_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_10_27_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_10_27_0  (
            .in0(_gnd_net_),
            .in1(N__20039),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_27_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_27_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_10_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(N__17576),
            .in2(N__21955),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_27_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_10_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__17570),
            .in2(N__21949),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_27_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_10_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(N__19727),
            .in2(N__21952),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_27_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_10_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__17582),
            .in2(N__21950),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_27_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_10_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(N__17615),
            .in2(N__21953),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_27_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_10_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_10_27_6  (
            .in0(_gnd_net_),
            .in1(N__19733),
            .in2(N__21951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_27_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_10_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(N__17477),
            .in2(N__21954),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_10_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_10_28_0  (
            .in0(_gnd_net_),
            .in1(N__17537),
            .in2(N__21965),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_28_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_10_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_10_28_1  (
            .in0(_gnd_net_),
            .in1(N__21964),
            .in2(N__17519),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_28_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_10_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17471),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_10_28_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_10_28_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_10_28_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_10_28_3  (
            .in0(N__24348),
            .in1(N__17468),
            .in2(N__17453),
            .in3(N__24459),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_10_28_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_10_28_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_10_28_4  (
            .in0(N__17495),
            .in1(N__20096),
            .in2(N__19964),
            .in3(N__19898),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_10_28_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_10_28_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_10_28_5  (
            .in0(N__23034),
            .in1(N__19784),
            .in2(N__19763),
            .in3(N__22992),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_28_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_28_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_10_28_6  (
            .in0(N__17563),
            .in1(N__22976),
            .in2(N__17552),
            .in3(N__22955),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_10_28_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_10_28_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_10_28_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_10_28_7  (
            .in0(N__17530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22933),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_10_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_10_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_10_29_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_10_29_0  (
            .in0(N__19933),
            .in1(N__19899),
            .in2(N__20102),
            .in3(N__21481),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_10_29_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_10_29_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_10_29_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_10_29_1  (
            .in0(N__19900),
            .in1(N__24023),
            .in2(N__19934),
            .in3(N__20100),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_10_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_10_29_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_10_29_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_10_29_3  (
            .in0(N__25893),
            .in1(N__17510),
            .in2(_gnd_net_),
            .in3(N__22118),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25185),
            .ce(N__26177),
            .sr(N__24811));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_10_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_10_29_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_10_29_4  (
            .in0(N__17489),
            .in1(N__25894),
            .in2(_gnd_net_),
            .in3(N__22001),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25185),
            .ce(N__26177),
            .sr(N__24811));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_10_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_10_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_10_29_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_10_29_5  (
            .in0(N__17621),
            .in1(N__24327),
            .in2(N__17591),
            .in3(N__24366),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_10_29_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_10_29_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_10_29_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_10_29_6  (
            .in0(N__17606),
            .in1(N__25895),
            .in2(_gnd_net_),
            .in3(N__22361),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25185),
            .ce(N__26177),
            .sr(N__24811));
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_11_11_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_0_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21108),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_11_11_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_1_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_1_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20981),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_11_11_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_2_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20872),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_11_11_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_3_LC_11_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_3_LC_11_11_3  (
            .in0(N__20788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_11_11_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_4_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_4_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20721),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_11_11_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_5_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_5_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26332),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_11_11_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_6_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_6_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20621),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_11_11_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH4data_esr_7_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH4data_esr_7_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20506),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25261),
            .ce(N__17948),
            .sr(N__24745));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_12_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__17915),
            .in2(N__17895),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_11_12_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_11_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__17723),
            .in2(N__17717),
            .in3(N__17708),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_11_12_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_11_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__17705),
            .in2(N__17699),
            .in3(N__17690),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNIRSJI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_11_12_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_11_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__17687),
            .in2(N__17681),
            .in3(N__17672),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIU0LI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_11_12_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_11_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__17669),
            .in2(N__20132),
            .in3(N__17663),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNI15MI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_11_12_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_11_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__17660),
            .in2(N__17654),
            .in3(N__17645),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNI49NI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_11_12_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_11_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__17642),
            .in2(N__17636),
            .in3(N__17627),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNI7DOI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_11_12_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_11_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__17732),
            .in2(_gnd_net_),
            .in3(N__17624),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIAHPI ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_11_13_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_11_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__17867),
            .in2(N__21948),
            .in3(N__17954),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIBJQI ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_13_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17951),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI8GVT_5_LC_11_13_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI8GVT_5_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI8GVT_5_LC_11_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_RNI8GVT_5_LC_11_13_2  (
            .in0(N__17773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24909),
            .lcout(\uart_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_13_3 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_11_13_3  (
            .in0(N__20439),
            .in1(N__17925),
            .in2(_gnd_net_),
            .in3(N__17888),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_544_i_l_ofx_LC_11_13_6 .C_ON=1'b0;
    defparam \scaler_4.N_544_i_l_ofx_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_544_i_l_ofx_LC_11_13_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_544_i_l_ofx_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__17761),
            .in2(_gnd_net_),
            .in3(N__17747),
            .lcout(\scaler_4.N_544_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_14_0 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__17861),
            .in2(_gnd_net_),
            .in3(N__17830),
            .lcout(\scaler_2.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_11_14_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH2data_esr_7_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH2data_esr_7_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20531),
            .lcout(frame_decoder_CH2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25243),
            .ce(N__17819),
            .sr(N__24757));
    defparam \uart_frame_decoder.state_1_RNIB3PK_5_LC_11_14_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIB3PK_5_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIB3PK_5_LC_11_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIB3PK_5_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__17798),
            .in2(_gnd_net_),
            .in3(N__23822),
            .lcout(\uart_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_14_7 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__17762),
            .in2(_gnd_net_),
            .in3(N__17746),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_15_0 .C_ON=1'b1;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__18065),
            .in2(N__18089),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.source_data_1_esr_6_LC_11_15_1 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_6_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_6_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_6_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__18040),
            .in2(N__18073),
            .in3(N__18047),
            .lcout(scaler_3_data_6),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_1 ),
            .carryout(\scaler_3.un2_source_data_0_cry_2 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_7_LC_11_15_2 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_7_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_7_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_7_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__18025),
            .in2(N__18044),
            .in3(N__18032),
            .lcout(scaler_3_data_7),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_2 ),
            .carryout(\scaler_3.un2_source_data_0_cry_3 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_8_LC_11_15_3 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_8_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_8_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_8_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__18010),
            .in2(N__18029),
            .in3(N__18017),
            .lcout(scaler_3_data_8),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_3 ),
            .carryout(\scaler_3.un2_source_data_0_cry_4 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_9_LC_11_15_4 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_9_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_9_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_9_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__17995),
            .in2(N__18014),
            .in3(N__18002),
            .lcout(scaler_3_data_9),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_4 ),
            .carryout(\scaler_3.un2_source_data_0_cry_5 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_10_LC_11_15_5 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_10_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_10_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_10_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__17980),
            .in2(N__17999),
            .in3(N__17987),
            .lcout(scaler_3_data_10),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_5 ),
            .carryout(\scaler_3.un2_source_data_0_cry_6 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_11_LC_11_15_6 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_11_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_11_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_11_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__17965),
            .in2(N__17984),
            .in3(N__17972),
            .lcout(scaler_3_data_11),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_6 ),
            .carryout(\scaler_3.un2_source_data_0_cry_7 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_12_LC_11_15_7 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_12_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_12_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_12_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__18166),
            .in2(N__17969),
            .in3(N__17957),
            .lcout(scaler_3_data_12),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_7 ),
            .carryout(\scaler_3.un2_source_data_0_cry_8 ),
            .clk(N__25236),
            .ce(N__21139),
            .sr(N__24761));
    defparam \scaler_3.source_data_1_esr_13_LC_11_16_0 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_13_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_13_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_13_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__18167),
            .in2(N__18155),
            .in3(N__18146),
            .lcout(scaler_3_data_13),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_9 ),
            .clk(N__25232),
            .ce(N__21140),
            .sr(N__24768));
    defparam \scaler_3.source_data_1_esr_14_LC_11_16_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_14_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_14_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_3.source_data_1_esr_14_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18143),
            .lcout(scaler_3_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25232),
            .ce(N__21140),
            .sr(N__24768));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_11_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__26257),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_11_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__20389),
            .in2(_gnd_net_),
            .in3(N__18128),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_11_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__20347),
            .in2(_gnd_net_),
            .in3(N__18116),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_11_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__20311),
            .in2(_gnd_net_),
            .in3(N__18113),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_11_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__20278),
            .in2(_gnd_net_),
            .in3(N__18098),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_11_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__21607),
            .in2(_gnd_net_),
            .in3(N__18095),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_11_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__21523),
            .in2(_gnd_net_),
            .in3(N__18092),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_11_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__21178),
            .in2(N__21920),
            .in3(N__18368),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_11_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_11_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__21155),
            .in2(_gnd_net_),
            .in3(N__18365),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25223),
            .ce(N__21738),
            .sr(N__24777));
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_11_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__18358),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_11_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__18337),
            .in2(_gnd_net_),
            .in3(N__18305),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_11_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_11_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__18301),
            .in2(_gnd_net_),
            .in3(N__18278),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_11_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__18268),
            .in2(_gnd_net_),
            .in3(N__18239),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_11_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_11_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__18229),
            .in2(_gnd_net_),
            .in3(N__18200),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_11_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_11_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18196),
            .in3(N__18170),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_11_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_11_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__18892),
            .in2(_gnd_net_),
            .in3(N__18866),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_11_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_11_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__21849),
            .in2(N__18856),
            .in3(N__18824),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_11_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_11_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__18821),
            .in2(_gnd_net_),
            .in3(N__18809),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25213),
            .ce(N__21726),
            .sr(N__24785));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__24256),
            .in2(_gnd_net_),
            .in3(N__24028),
            .lcout(\ppm_encoder_1.N_143_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_13_LC_11_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_11_21_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_11_21_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_11_21_2  (
            .in0(N__21182),
            .in1(N__18806),
            .in2(N__25550),
            .in3(N__22389),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25207),
            .ce(),
            .sr(N__24790));
    defparam \ppm_encoder_1.rudder_9_LC_11_21_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_11_21_4 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_11_21_4  (
            .in0(N__20315),
            .in1(N__25533),
            .in2(N__18797),
            .in3(N__19132),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25207),
            .ce(),
            .sr(N__24790));
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_11_22_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_11_22_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_11_22_0  (
            .in0(N__22294),
            .in1(N__21757),
            .in2(N__18780),
            .in3(N__18688),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_11_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_11_22_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_11_22_1  (
            .in0(N__18584),
            .in1(_gnd_net_),
            .in2(N__18566),
            .in3(N__18374),
            .lcout(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_11_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_11_22_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_11_22_2  (
            .in0(N__22270),
            .in1(N__18535),
            .in2(N__19175),
            .in3(N__18453),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_11_22_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_11_22_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_11_22_3  (
            .in0(N__19174),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__21758),
            .lcout(\ppm_encoder_1.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_22_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_22_4 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_22_4  (
            .in0(N__23222),
            .in1(N__19154),
            .in2(N__23277),
            .in3(N__19131),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_11_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_11_22_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_11_22_5  (
            .in0(N__19411),
            .in1(N__23220),
            .in2(N__19100),
            .in3(N__23258),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_11_22_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_11_22_6 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_11_22_6  (
            .in0(N__23219),
            .in1(N__19079),
            .in2(N__23276),
            .in3(N__19058),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_22_7 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_22_7  (
            .in0(N__19036),
            .in1(N__23259),
            .in2(N__19001),
            .in3(N__23221),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_11_23_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_11_23_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_11_23_0  (
            .in0(N__19703),
            .in1(N__18965),
            .in2(N__19566),
            .in3(N__18953),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25199),
            .ce(),
            .sr(N__24800));
    defparam \ppm_encoder_1.init_pulses_5_LC_11_23_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_11_23_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_11_23_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_11_23_3  (
            .in0(N__19704),
            .in1(N__18941),
            .in2(N__19567),
            .in3(N__18929),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25199),
            .ce(),
            .sr(N__24800));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_11_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_11_23_4 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_11_23_4  (
            .in0(N__22760),
            .in1(N__22098),
            .in2(N__23693),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_11_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_11_23_5 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__23631),
            .in2(N__22103),
            .in3(N__22759),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_11_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_11_23_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_11_23_7  (
            .in0(N__19705),
            .in1(N__19595),
            .in2(N__19568),
            .in3(N__19430),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25199),
            .ce(),
            .sr(N__24800));
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_11_24_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_11_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_c_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__19397),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_24_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__19360),
            .in2(_gnd_net_),
            .in3(N__19328),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_24_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__19324),
            .in2(_gnd_net_),
            .in3(N__19289),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_24_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__19253),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_24_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__19246),
            .in2(_gnd_net_),
            .in3(N__19220),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_24_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__19213),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_24_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__19873),
            .in2(_gnd_net_),
            .in3(N__19838),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_24_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__25591),
            .in2(N__21923),
            .in3(N__19835),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_25_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__19832),
            .in2(_gnd_net_),
            .in3(N__19814),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25193),
            .ce(N__21740),
            .sr(N__24806));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_11_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_11_26_1  (
            .in0(N__25884),
            .in1(N__19811),
            .in2(_gnd_net_),
            .in3(N__19796),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25189),
            .ce(N__26171),
            .sr(N__24807));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_11_26_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_11_26_2  (
            .in0(N__19775),
            .in1(N__25885),
            .in2(_gnd_net_),
            .in3(N__22064),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25189),
            .ce(N__26171),
            .sr(N__24807));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_26_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_11_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_11_26_3  (
            .in0(N__25883),
            .in1(N__19748),
            .in2(_gnd_net_),
            .in3(N__22373),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25189),
            .ce(N__26171),
            .sr(N__24807));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_11_26_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_11_26_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_11_26_4  (
            .in0(N__23318),
            .in1(N__22862),
            .in2(N__19742),
            .in3(N__24440),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_26_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_26_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_11_26_6  (
            .in0(N__23017),
            .in1(N__23348),
            .in2(N__23372),
            .in3(N__23057),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_11_27_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_11_27_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_11_27_1  (
            .in0(N__26066),
            .in1(N__25781),
            .in2(_gnd_net_),
            .in3(N__20003),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_27_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_27_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_11_27_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_11_27_2  (
            .in0(_gnd_net_),
            .in1(N__25891),
            .in2(N__20051),
            .in3(N__23063),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25188),
            .ce(N__26176),
            .sr(N__24809));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_27_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_27_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_11_27_3  (
            .in0(N__19925),
            .in1(N__24309),
            .in2(N__20048),
            .in3(N__20009),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_27_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_11_27_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_11_27_4  (
            .in0(N__23310),
            .in1(N__23225),
            .in2(_gnd_net_),
            .in3(N__20033),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25188),
            .ce(N__26176),
            .sr(N__24809));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_11_27_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_11_27_6 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(N__20002),
            .in2(N__25804),
            .in3(N__26067),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_27_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_11_27_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_11_27_7  (
            .in0(N__22475),
            .in1(_gnd_net_),
            .in2(N__19967),
            .in3(N__25892),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25188),
            .ce(N__26176),
            .sr(N__24809));
    defparam \ppm_encoder_1.counter_0_LC_11_28_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_11_28_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_11_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_11_28_0  (
            .in0(_gnd_net_),
            .in1(N__24311),
            .in2(N__19955),
            .in3(N__19954),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_28_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_1_LC_11_28_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_11_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_11_28_1  (
            .in0(_gnd_net_),
            .in1(N__19932),
            .in2(_gnd_net_),
            .in3(N__19904),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_2_LC_11_28_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_11_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_11_28_2  (
            .in0(_gnd_net_),
            .in1(N__19901),
            .in2(_gnd_net_),
            .in3(N__19880),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_3_LC_11_28_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_11_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_11_28_3  (
            .in0(_gnd_net_),
            .in1(N__20101),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_4_LC_11_28_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_11_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_11_28_4  (
            .in0(_gnd_net_),
            .in1(N__22994),
            .in2(_gnd_net_),
            .in3(N__20075),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_5_LC_11_28_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_11_28_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_11_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_11_28_5  (
            .in0(_gnd_net_),
            .in1(N__23036),
            .in2(_gnd_net_),
            .in3(N__20072),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_6_LC_11_28_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_11_28_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_11_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_11_28_6  (
            .in0(_gnd_net_),
            .in1(N__23056),
            .in2(_gnd_net_),
            .in3(N__20069),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_7_LC_11_28_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_11_28_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_11_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_11_28_7  (
            .in0(_gnd_net_),
            .in1(N__23016),
            .in2(_gnd_net_),
            .in3(N__20066),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__25186),
            .ce(),
            .sr(N__20201));
    defparam \ppm_encoder_1.counter_8_LC_11_29_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_11_29_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_11_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_11_29_0  (
            .in0(_gnd_net_),
            .in1(N__24461),
            .in2(_gnd_net_),
            .in3(N__20063),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_29_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_9_LC_11_29_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_11_29_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_11_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_11_29_1  (
            .in0(_gnd_net_),
            .in1(N__24350),
            .in2(_gnd_net_),
            .in3(N__20060),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_10_LC_11_29_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_11_29_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_11_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_11_29_2  (
            .in0(_gnd_net_),
            .in1(N__24368),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_11_LC_11_29_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_11_29_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_11_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_11_29_3  (
            .in0(_gnd_net_),
            .in1(N__24331),
            .in2(_gnd_net_),
            .in3(N__20054),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_12_LC_11_29_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_11_29_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_11_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_11_29_4  (
            .in0(_gnd_net_),
            .in1(N__24439),
            .in2(_gnd_net_),
            .in3(N__20222),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_13_LC_11_29_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_11_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_11_29_5  (
            .in0(_gnd_net_),
            .in1(N__22861),
            .in2(_gnd_net_),
            .in3(N__20219),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_14_LC_11_29_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_11_29_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_11_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_11_29_6  (
            .in0(_gnd_net_),
            .in1(N__22882),
            .in2(_gnd_net_),
            .in3(N__20216),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_15_LC_11_29_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_11_29_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_11_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_11_29_7  (
            .in0(_gnd_net_),
            .in1(N__22906),
            .in2(_gnd_net_),
            .in3(N__20213),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__25184),
            .ce(),
            .sr(N__20200));
    defparam \ppm_encoder_1.counter_16_LC_11_30_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_11_30_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_11_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_11_30_0  (
            .in0(_gnd_net_),
            .in1(N__22954),
            .in2(_gnd_net_),
            .in3(N__20210),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_30_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__25183),
            .ce(),
            .sr(N__20199));
    defparam \ppm_encoder_1.counter_17_LC_11_30_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_11_30_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_11_30_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_11_30_1  (
            .in0(_gnd_net_),
            .in1(N__22975),
            .in2(_gnd_net_),
            .in3(N__20207),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__25183),
            .ce(),
            .sr(N__20199));
    defparam \ppm_encoder_1.counter_18_LC_11_30_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_11_30_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_11_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_11_30_2  (
            .in0(_gnd_net_),
            .in1(N__22932),
            .in2(_gnd_net_),
            .in3(N__20204),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25183),
            .ce(),
            .sr(N__20199));
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_12_1_2 .C_ON=1'b0;
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \scaler_1.source_data_1_esr_ctle_14_LC_12_1_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_1.source_data_1_esr_ctle_14_LC_12_1_2  (
            .in0(_gnd_net_),
            .in1(N__20186),
            .in2(_gnd_net_),
            .in3(N__24895),
            .lcout(pc_frame_decoder_dv_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_12_12_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_offset4data_esr_4_LC_12_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_offset4data_esr_4_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20729),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25247),
            .ce(N__20123),
            .sr(N__24754));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_13_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__20432),
            .in2(N__20450),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_12_13_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_12_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__20407),
            .in2(N__20440),
            .in3(N__20414),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_7_LC_12_13_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__20359),
            .in2(N__20411),
            .in3(N__20366),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_8_LC_12_13_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_12_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__20323),
            .in2(N__20363),
            .in3(N__20330),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_9_LC_12_13_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_12_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__20287),
            .in2(N__20327),
            .in3(N__20294),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_10_LC_12_13_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_12_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__20248),
            .in2(N__20291),
            .in3(N__20255),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_11_LC_12_13_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_12_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__20233),
            .in2(N__20252),
            .in3(N__20240),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_12_LC_12_13_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_12_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(N__20237),
            .in3(N__20225),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__25242),
            .ce(N__21135),
            .sr(N__24758));
    defparam \scaler_4.source_data_1_esr_13_LC_12_14_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_12_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__21203),
            .in2(N__21191),
            .in3(N__21161),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__25234),
            .ce(N__21136),
            .sr(N__24762));
    defparam \scaler_4.source_data_1_esr_14_LC_12_14_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21158),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25234),
            .ce(N__21136),
            .sr(N__24762));
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_12_15_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_0_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_0_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(frame_decoder_CH3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_12_15_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_1_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_1_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(frame_decoder_CH3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_12_15_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_2_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_2_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20900),
            .lcout(frame_decoder_CH3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_12_15_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_3_LC_12_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_3_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20808),
            .lcout(frame_decoder_CH3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_12_15_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_4_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_4_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20728),
            .lcout(frame_decoder_CH3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_12_15_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_6_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_6_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(frame_decoder_CH3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_12_15_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_7_LC_12_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_7_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20537),
            .lcout(frame_decoder_CH3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25230),
            .ce(N__26270),
            .sr(N__24769));
    defparam \uart_frame_decoder.state_1_RNI80PK_2_LC_12_16_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI80PK_2_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI80PK_2_LC_12_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNI80PK_2_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__23866),
            .in2(_gnd_net_),
            .in3(N__23788),
            .lcout(\uart_frame_decoder.source_CH1data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_12_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_c_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_c_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__21334),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__21316),
            .in2(_gnd_net_),
            .in3(N__21287),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__21655),
            .in2(_gnd_net_),
            .in3(N__21284),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__21400),
            .in2(_gnd_net_),
            .in3(N__21281),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__21568),
            .in2(_gnd_net_),
            .in3(N__21278),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__21274),
            .in2(_gnd_net_),
            .in3(N__21245),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21238),
            .in3(N__21206),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__21986),
            .in2(N__21921),
            .in3(N__21773),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__21770),
            .in2(_gnd_net_),
            .in3(N__21761),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25217),
            .ce(N__21730),
            .sr(N__24780));
    defparam \ppm_encoder_1.throttle_8_LC_12_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_12_19_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_12_19_2  (
            .in0(N__21668),
            .in1(N__21659),
            .in2(N__25547),
            .in3(N__21633),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25211),
            .ce(),
            .sr(N__24786));
    defparam \ppm_encoder_1.rudder_11_LC_12_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_12_20_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_12_20_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_12_20_2  (
            .in0(N__21611),
            .in1(N__21590),
            .in2(N__25544),
            .in3(N__22530),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25205),
            .ce(),
            .sr(N__24791));
    defparam \ppm_encoder_1.throttle_10_LC_12_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_12_20_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_12_20_5  (
            .in0(N__21581),
            .in1(N__21572),
            .in2(N__21549),
            .in3(N__25505),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25205),
            .ce(),
            .sr(N__24791));
    defparam \ppm_encoder_1.rudder_12_LC_12_21_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_12_21_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_12_21_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_12_21_1  (
            .in0(N__21527),
            .in1(N__21503),
            .in2(N__25545),
            .in3(N__22443),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25201),
            .ce(),
            .sr(N__24797));
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_21_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_12_21_2 .LUT_INIT=16'b1110111101000100;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_12_21_2  (
            .in0(N__24380),
            .in1(N__21491),
            .in2(N__21485),
            .in3(N__21424),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25201),
            .ce(),
            .sr(N__24797));
    defparam \ppm_encoder_1.throttle_9_LC_12_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_12_21_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_12_21_3  (
            .in0(N__21413),
            .in1(N__21404),
            .in2(N__25546),
            .in3(N__25632),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25201),
            .ce(),
            .sr(N__24797));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_12_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_12_22_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_12_22_1  (
            .in0(N__25732),
            .in1(N__22249),
            .in2(_gnd_net_),
            .in3(N__22194),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_22_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_22_2 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_22_2  (
            .in0(N__23223),
            .in1(N__22331),
            .in2(N__22301),
            .in3(N__22298),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_22_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_12_22_5  (
            .in0(N__26031),
            .in1(N__22277),
            .in2(_gnd_net_),
            .in3(N__22271),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_12_22_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_12_22_7 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_12_22_7  (
            .in0(N__25733),
            .in1(N__24928),
            .in2(N__26065),
            .in3(N__23698),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25197),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_12_23_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_12_23_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_12_23_4  (
            .in0(N__22253),
            .in1(N__25734),
            .in2(_gnd_net_),
            .in3(N__22199),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_12_23_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_12_23_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_12_23_5  (
            .in0(N__23251),
            .in1(N__23211),
            .in2(N__22148),
            .in3(N__22145),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_23_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_23_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_12_23_7  (
            .in0(N__23212),
            .in1(N__22102),
            .in2(N__23275),
            .in3(N__22085),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_12_24_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_12_24_0 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_12_24_0  (
            .in0(N__22055),
            .in1(N__23206),
            .in2(N__23299),
            .in3(N__22028),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_24_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_24_1 .LUT_INIT=16'b1010111110111010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_24_1  (
            .in0(N__24929),
            .in1(N__22841),
            .in2(N__23713),
            .in3(N__25979),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25191),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_24_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_24_2  (
            .in0(N__25978),
            .in1(N__22592),
            .in2(_gnd_net_),
            .in3(N__22580),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_24_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_24_7  (
            .in0(N__23205),
            .in1(N__22556),
            .in2(_gnd_net_),
            .in3(N__22535),
            .lcout(\ppm_encoder_1.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_12_25_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_12_25_1 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_12_25_1  (
            .in0(N__23308),
            .in1(N__23209),
            .in2(N__23116),
            .in3(N__22502),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_12_25_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_12_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_12_25_2  (
            .in0(N__23207),
            .in1(N__22463),
            .in2(_gnd_net_),
            .in3(N__22445),
            .lcout(),
            .ltout(\ppm_encoder_1.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_25_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_25_3 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_25_3  (
            .in0(N__23109),
            .in1(_gnd_net_),
            .in2(N__22421),
            .in3(N__23301),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_12_25_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_12_25_4 .LUT_INIT=16'b1110111101001111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_12_25_4  (
            .in0(N__23208),
            .in1(N__22418),
            .in2(N__23311),
            .in3(N__22400),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_25_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_25_5  (
            .in0(N__23108),
            .in1(N__23300),
            .in2(_gnd_net_),
            .in3(N__22367),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_25_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_25_6 .LUT_INIT=16'b1110111101001111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_12_25_6  (
            .in0(N__23210),
            .in1(N__22349),
            .in2(N__23312),
            .in3(N__26234),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_25_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_25_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_25_7  (
            .in0(_gnd_net_),
            .in1(N__24917),
            .in2(_gnd_net_),
            .in3(N__23694),
            .lcout(\ppm_encoder_1.N_614_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_12_26_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_12_26_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_12_26_1  (
            .in0(N__23396),
            .in1(N__25863),
            .in2(_gnd_net_),
            .in3(N__23384),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25187),
            .ce(N__26160),
            .sr(N__24810));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_12_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_12_26_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_12_26_2  (
            .in0(N__25862),
            .in1(N__23363),
            .in2(_gnd_net_),
            .in3(N__23354),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25187),
            .ce(N__26160),
            .sr(N__24810));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_12_26_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_12_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_12_26_5  (
            .in0(N__25861),
            .in1(N__23342),
            .in2(_gnd_net_),
            .in3(N__23324),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25187),
            .ce(N__26160),
            .sr(N__24810));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_12_27_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_12_27_0 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_12_27_0  (
            .in0(N__23309),
            .in1(N__23224),
            .in2(N__23120),
            .in3(N__23090),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_28_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_12_28_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_12_28_1  (
            .in0(N__23055),
            .in1(N__23035),
            .in2(N__23018),
            .in3(N__22993),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_12_29_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_12_29_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_12_29_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_12_29_0  (
            .in0(N__22974),
            .in1(N__22953),
            .in2(N__22934),
            .in3(N__22905),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_12_29_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_12_29_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_12_29_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_12_29_2  (
            .in0(_gnd_net_),
            .in1(N__22881),
            .in2(_gnd_net_),
            .in3(N__22860),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_12_29_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_12_29_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_12_29_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_12_29_3  (
            .in0(N__24467),
            .in1(N__24460),
            .in2(N__24443),
            .in3(N__24438),
            .lcout(\ppm_encoder_1.N_148_17 ),
            .ltout(\ppm_encoder_1.N_148_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_12_29_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_12_29_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_12_29_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_12_29_4  (
            .in0(N__24292),
            .in1(N__24406),
            .in2(N__24419),
            .in3(N__24416),
            .lcout(\ppm_encoder_1.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_12_29_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_12_29_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_12_29_5  (
            .in0(N__24407),
            .in1(N__24398),
            .in2(N__24392),
            .in3(N__24293),
            .lcout(\ppm_encoder_1.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_12_29_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_12_29_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_12_29_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_12_29_7  (
            .in0(N__24367),
            .in1(N__24349),
            .in2(N__24332),
            .in3(N__24310),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_12_30_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_12_30_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_12_30_1 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_12_30_1  (
            .in0(N__24268),
            .in1(N__24252),
            .in2(N__24203),
            .in3(N__24029),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_2_LC_13_13_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_2_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_2_LC_13_13_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_2_LC_13_13_0  (
            .in0(N__23963),
            .in1(N__23942),
            .in2(N__23867),
            .in3(N__23915),
            .lcout(\uart_frame_decoder.state_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25249),
            .ce(),
            .sr(N__24763));
    defparam \uart_frame_decoder.state_1_RNIA2PK_4_LC_13_13_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIA2PK_4_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIA2PK_4_LC_13_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNIA2PK_4_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__23846),
            .in2(_gnd_net_),
            .in3(N__23819),
            .lcout(\uart_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI7FVT_4_LC_13_14_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI7FVT_4_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI7FVT_4_LC_13_14_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_frame_decoder.state_1_RNI7FVT_4_LC_13_14_3  (
            .in0(N__26374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24910),
            .lcout(\uart_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_13_15_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_CH3data_esr_5_LC_13_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.source_CH3data_esr_5_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26362),
            .lcout(frame_decoder_CH3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25237),
            .ce(N__26269),
            .sr(N__24773));
    defparam \ppm_encoder_1.rudder_6_LC_13_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_13_19_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_13_19_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_13_19_0  (
            .in0(N__25512),
            .in1(N__26258),
            .in2(_gnd_net_),
            .in3(N__26226),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25219),
            .ce(),
            .sr(N__24792));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_13_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_13_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_13_22_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_13_22_1  (
            .in0(N__26204),
            .in1(N__25896),
            .in2(_gnd_net_),
            .in3(N__26198),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25203),
            .ce(N__26167),
            .sr(N__24803));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_13_26_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_13_26_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_13_26_2  (
            .in0(N__26064),
            .in1(N__25795),
            .in2(_gnd_net_),
            .in3(N__25943),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_21_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_21_2  (
            .in0(N__25796),
            .in1(N__25657),
            .in2(_gnd_net_),
            .in3(N__25634),
            .lcout(\ppm_encoder_1.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_14_25_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_14_25_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_14_25_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_14_25_5  (
            .in0(N__25598),
            .in1(N__25571),
            .in2(N__25558),
            .in3(N__25320),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25195),
            .ce(),
            .sr(N__24812));
endmodule // Pc2drone
