-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 10 2019 19:42:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2Drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2Drone
entity Pc2Drone is
port (
    data : out std_logic_vector(7 downto 0);
    uart_input : in std_logic;
    data_rdy : out std_logic;
    uart_input_debug : out std_logic;
    clk_system : in std_logic);
end Pc2Drone;

-- Architecture of Pc2Drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2Drone is

signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2014\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1917\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1884\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1844\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1837\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1659\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1611\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1529\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1476\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1393\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1376\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1372\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1367\ : std_logic;
signal \N__1366\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1356\ : std_logic;
signal \N__1355\ : std_logic;
signal \N__1350\ : std_logic;
signal \N__1345\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1337\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1325\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1313\ : std_logic;
signal \N__1310\ : std_logic;
signal \N__1307\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1303\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1295\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1280\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1271\ : std_logic;
signal \N__1268\ : std_logic;
signal \N__1265\ : std_logic;
signal \N__1262\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1260\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1253\ : std_logic;
signal \N__1244\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1237\ : std_logic;
signal \N__1236\ : std_logic;
signal \N__1229\ : std_logic;
signal \N__1226\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1214\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1208\ : std_logic;
signal \N__1205\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \uart.CO0_0_cascade_\ : std_logic;
signal \uart.bit_Count_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \uart.CO1_1_cascade_\ : std_logic;
signal \uart.bit_Count_RNO_2Z0Z_2\ : std_logic;
signal \uart.bit_Count_RNO_1Z0Z_1\ : std_logic;
signal \uart.state_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \uart.state_RNO_2Z0Z_2\ : std_logic;
signal \uart.N_170_cascade_\ : std_logic;
signal \uart.stateZ0Z_2\ : std_logic;
signal \uart.stateZ0Z_1\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \uart.N_44_0\ : std_logic;
signal \uart.N_147_0_cascade_\ : std_logic;
signal \uart.timer_Count_RNITC202Z0Z_6\ : std_logic;
signal \uart.timer_Count_RNIGLM11Z0Z_6_cascade_\ : std_logic;
signal \uart.un1_state_7_0_0\ : std_logic;
signal \uart.un1_state_7_0_0_cascade_\ : std_logic;
signal \uart.N_177\ : std_logic;
signal \uart.un1_state_5\ : std_logic;
signal \uart.state_RNO_0Z0Z_3\ : std_logic;
signal \uart.state_RNO_1Z0Z_3\ : std_logic;
signal \uart.N_147_0\ : std_logic;
signal \uart.N_159\ : std_logic;
signal \uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_\ : std_logic;
signal \uart.un1_state_2_0_a3_0_cascade_\ : std_logic;
signal \uart.timer_CountZ0Z_6\ : std_logic;
signal \uart.timer_Count_fastZ0Z_6\ : std_logic;
signal \uart.un1_state_4_0_a2_iso_cascade_\ : std_logic;
signal \uart.N_38_0\ : std_logic;
signal \uart.N_165_1\ : std_logic;
signal \uart.timer_Count_RNIICSG1Z0Z_6\ : std_logic;
signal \uart.N_175_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_1\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \uart.timer_Count_6_repZ0Z1\ : std_logic;
signal \uart.un4_timer_Count_1_c2\ : std_logic;
signal \uart.timer_Count_RNIMLMA1Z0Z_1_cascade_\ : std_logic;
signal \uart.un4_timer_Count_1_c5\ : std_logic;
signal \uart.un4_timer_Count_1_c5_cascade_\ : std_logic;
signal \uart.timer_CountZ0Z_3\ : std_logic;
signal \uart.timer_CountZ0Z_2\ : std_logic;
signal \uart.stateZ0Z_3\ : std_logic;
signal \uart.timer_Count_RNIHJ661Z0Z_3_cascade_\ : std_logic;
signal \uart.timer_CountZ0Z_5\ : std_logic;
signal \uart.state_0_sqmuxa_1_d\ : std_logic;
signal \uart.timer_CountZ0Z_0\ : std_logic;
signal \uart.timer_CountZ0Z_1\ : std_logic;
signal \uart.un1_timer_Count_0_sqmuxa_0\ : std_logic;
signal \uart.timer_CountZ0Z_4\ : std_logic;
signal \uart.timer_CountZ0Z_7\ : std_logic;
signal \uart.N_28_mux_i_i_0\ : std_logic;
signal \uart.N_22_mux\ : std_logic;
signal data_rdy_c : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_0\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_4\ : std_logic;
signal \uart.N_39_0\ : std_logic;
signal \uart.N_40_0\ : std_logic;
signal \uart.timer_Count_6_rep1_RNI1B4SZ0\ : std_logic;
signal \uart.timer_Count_6_rep1_RNI02QZ0Z61\ : std_logic;
signal \uart.N_145_0\ : std_logic;
signal \uart.timer_Count28\ : std_logic;
signal \uart.timer_Count28_cascade_\ : std_logic;
signal \uart.stateZ0Z_4\ : std_logic;
signal \uart.bit_CountZ0Z_1\ : std_logic;
signal \uart.bit_CountZ0Z_0\ : std_logic;
signal \uart.bit_CountZ0Z_2\ : std_logic;
signal \uart.N_175\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \uart.data_Aux_esr_RNO_0Z0Z_6\ : std_logic;
signal \uart.state_1_sqmuxa\ : std_logic;
signal \uart.N_42_0\ : std_logic;
signal \uart.N_41_0\ : std_logic;
signal \uart.N_37_0\ : std_logic;
signal \uart.data_AuxZ0Z_0\ : std_logic;
signal data_c_0 : std_logic;
signal \uart.data_AuxZ0Z_1\ : std_logic;
signal data_c_1 : std_logic;
signal \uart.data_AuxZ0Z_2\ : std_logic;
signal data_c_2 : std_logic;
signal \uart.data_AuxZ0Z_3\ : std_logic;
signal data_c_3 : std_logic;
signal \uart.data_AuxZ0Z_5\ : std_logic;
signal data_c_5 : std_logic;
signal data_c_6 : std_logic;
signal \uart.data_AuxZ0Z_7\ : std_logic;
signal data_c_7 : std_logic;
signal \uart.data_AuxZ0Z_4\ : std_logic;
signal data_c_4 : std_logic;
signal \uart.state_1_sqmuxa_0\ : std_logic;
signal \uart.state_RNIVF8I3Z0Z_4\ : std_logic;
signal uart_input_c : std_logic;
signal \uart.data_AuxZ0Z_6\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal \uart.N_43_0\ : std_logic;
signal \uart.un1_state_4_0_a2_iso\ : std_logic;

signal clk_system_wire : std_logic;
signal data_wire : std_logic_vector(7 downto 0);
signal uart_input_wire : std_logic;
signal data_rdy_wire : std_logic;
signal uart_input_debug_wire : std_logic;

begin
    clk_system_wire <= clk_system;
    data <= data_wire;
    uart_input_wire <= uart_input;
    data_rdy <= data_rdy_wire;
    uart_input_debug <= uart_input_debug_wire;

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3231\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3233\,
            DIN => \N__3232\,
            DOUT => \N__3231\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3233\,
            PADOUT => \N__3232\,
            PADIN => \N__3231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3222\,
            DIN => \N__3221\,
            DOUT => \N__3220\,
            PACKAGEPIN => data_wire(2)
        );

    \data_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3222\,
            PADOUT => \N__3221\,
            PADIN => \N__3220\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3213\,
            DIN => \N__3212\,
            DOUT => \N__3211\,
            PACKAGEPIN => data_wire(6)
        );

    \data_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3213\,
            PADOUT => \N__3212\,
            PADIN => \N__3211\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3032\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3204\,
            DIN => \N__3203\,
            DOUT => \N__3202\,
            PACKAGEPIN => uart_input_wire
        );

    \uart_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3204\,
            PADOUT => \N__3203\,
            PADIN => \N__3202\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3195\,
            DIN => \N__3194\,
            DOUT => \N__3193\,
            PACKAGEPIN => data_wire(1)
        );

    \data_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3195\,
            PADOUT => \N__3194\,
            PADIN => \N__3193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2330\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3186\,
            DIN => \N__3185\,
            DOUT => \N__3184\,
            PACKAGEPIN => data_wire(5)
        );

    \data_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3186\,
            PADOUT => \N__3185\,
            PADIN => \N__3184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3047\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3177\,
            DIN => \N__3176\,
            DOUT => \N__3175\,
            PACKAGEPIN => data_wire(0)
        );

    \data_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3177\,
            PADOUT => \N__3176\,
            PADIN => \N__3175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2357\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3168\,
            DIN => \N__3167\,
            DOUT => \N__3166\,
            PACKAGEPIN => data_wire(4)
        );

    \data_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3168\,
            PADOUT => \N__3167\,
            PADIN => \N__3166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2972\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_rdy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3159\,
            DIN => \N__3158\,
            DOUT => \N__3157\,
            PACKAGEPIN => data_rdy_wire
        );

    \data_rdy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3159\,
            PADOUT => \N__3158\,
            PADIN => \N__3157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2309\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3150\,
            DIN => \N__3149\,
            DOUT => \N__3148\,
            PACKAGEPIN => data_wire(3)
        );

    \data_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3150\,
            PADOUT => \N__3149\,
            PADIN => \N__3148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3141\,
            DIN => \N__3140\,
            DOUT => \N__3139\,
            PACKAGEPIN => uart_input_debug_wire
        );

    \uart_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3141\,
            PADOUT => \N__3140\,
            PADIN => \N__3139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2806\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \data_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3132\,
            DIN => \N__3131\,
            DOUT => \N__3130\,
            PACKAGEPIN => data_wire(7)
        );

    \data_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3132\,
            PADOUT => \N__3131\,
            PADIN => \N__3130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__739\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3110\,
            I => \uart.data_AuxZ0Z_2\
        );

    \I__737\ : IoInMux
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__735\ : Span4Mux_s3_v
    port map (
            O => \N__3101\,
            I => \N__3098\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__733\ : Span12Mux_s8_h
    port map (
            O => \N__3095\,
            I => \N__3092\
        );

    \I__732\ : Span12Mux_v
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__3089\,
            I => data_c_2
        );

    \I__730\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3083\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__728\ : IoInMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__726\ : Span4Mux_s3_v
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__725\ : Span4Mux_h
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__724\ : Span4Mux_h
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__723\ : Sp12to4
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__722\ : Span12Mux_v
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__3059\,
            I => data_c_3
        );

    \I__720\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__718\ : Odrv4
    port map (
            O => \N__3050\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__717\ : IoInMux
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__715\ : Sp12to4
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__714\ : Span12Mux_v
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__713\ : Odrv12
    port map (
            O => \N__3035\,
            I => data_c_5
        );

    \I__712\ : IoInMux
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__710\ : IoSpan4Mux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__709\ : Span4Mux_s0_v
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__708\ : Sp12to4
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__707\ : Span12Mux_v
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__706\ : Odrv12
    port map (
            O => \N__3014\,
            I => data_c_6
        );

    \I__705\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__3002\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__701\ : IoInMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__699\ : IoSpan4Mux
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__698\ : Sp12to4
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__697\ : Span12Mux_v
    port map (
            O => \N__2987\,
            I => \N__2984\
        );

    \I__696\ : Odrv12
    port map (
            O => \N__2984\,
            I => data_c_7
        );

    \I__695\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__2975\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__692\ : IoInMux
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__690\ : Span4Mux_s3_v
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__688\ : Span4Mux_v
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__2957\,
            I => data_c_4
        );

    \I__686\ : CEMux
    port map (
            O => \N__2954\,
            I => \N__2950\
        );

    \I__685\ : CEMux
    port map (
            O => \N__2953\,
            I => \N__2947\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2944\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__2944\,
            I => \uart.state_1_sqmuxa_0\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__2941\,
            I => \uart.state_1_sqmuxa_0\
        );

    \I__680\ : SRMux
    port map (
            O => \N__2936\,
            I => \N__2933\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__678\ : Span4Mux_v
    port map (
            O => \N__2930\,
            I => \N__2926\
        );

    \I__677\ : SRMux
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__2926\,
            I => \N__2917\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__2923\,
            I => \N__2917\
        );

    \I__674\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2914\
        );

    \I__673\ : Odrv12
    port map (
            O => \N__2917\,
            I => \uart.state_RNIVF8I3Z0Z_4\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__2914\,
            I => \uart.state_RNIVF8I3Z0Z_4\
        );

    \I__671\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2903\
        );

    \I__670\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2898\
        );

    \I__669\ : InMux
    port map (
            O => \N__2907\,
            I => \N__2894\
        );

    \I__668\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2891\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__2903\,
            I => \N__2887\
        );

    \I__666\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2884\
        );

    \I__665\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2881\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__2898\,
            I => \N__2878\
        );

    \I__663\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2875\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2870\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__2891\,
            I => \N__2870\
        );

    \I__660\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2867\
        );

    \I__659\ : Span4Mux_h
    port map (
            O => \N__2887\,
            I => \N__2859\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__2884\,
            I => \N__2859\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__2881\,
            I => \N__2859\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__2878\,
            I => \N__2851\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__2875\,
            I => \N__2851\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__2870\,
            I => \N__2846\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__2867\,
            I => \N__2846\
        );

    \I__652\ : InMux
    port map (
            O => \N__2866\,
            I => \N__2843\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__2859\,
            I => \N__2840\
        );

    \I__650\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2837\
        );

    \I__649\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2834\
        );

    \I__648\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2831\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__2851\,
            I => \N__2828\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__2846\,
            I => \N__2825\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__2843\,
            I => \N__2822\
        );

    \I__644\ : Span4Mux_h
    port map (
            O => \N__2840\,
            I => \N__2819\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__2837\,
            I => \N__2812\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__2834\,
            I => \N__2812\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__2831\,
            I => \N__2812\
        );

    \I__640\ : Sp12to4
    port map (
            O => \N__2828\,
            I => \N__2807\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__2825\,
            I => \N__2807\
        );

    \I__638\ : Span12Mux_h
    port map (
            O => \N__2822\,
            I => \N__2803\
        );

    \I__637\ : Sp12to4
    port map (
            O => \N__2819\,
            I => \N__2798\
        );

    \I__636\ : Span12Mux_h
    port map (
            O => \N__2812\,
            I => \N__2798\
        );

    \I__635\ : Span12Mux_h
    port map (
            O => \N__2807\,
            I => \N__2795\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__2806\,
            I => \N__2792\
        );

    \I__633\ : Span12Mux_v
    port map (
            O => \N__2803\,
            I => \N__2789\
        );

    \I__632\ : Span12Mux_v
    port map (
            O => \N__2798\,
            I => \N__2786\
        );

    \I__631\ : Span12Mux_v
    port map (
            O => \N__2795\,
            I => \N__2783\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__2792\,
            I => \N__2780\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__2789\,
            I => uart_input_c
        );

    \I__628\ : Odrv12
    port map (
            O => \N__2786\,
            I => uart_input_c
        );

    \I__627\ : Odrv12
    port map (
            O => \N__2783\,
            I => uart_input_c
        );

    \I__626\ : Odrv4
    port map (
            O => \N__2780\,
            I => uart_input_c
        );

    \I__625\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2768\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__2765\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__622\ : ClkMux
    port map (
            O => \N__2762\,
            I => \N__2702\
        );

    \I__621\ : ClkMux
    port map (
            O => \N__2761\,
            I => \N__2702\
        );

    \I__620\ : ClkMux
    port map (
            O => \N__2760\,
            I => \N__2702\
        );

    \I__619\ : ClkMux
    port map (
            O => \N__2759\,
            I => \N__2702\
        );

    \I__618\ : ClkMux
    port map (
            O => \N__2758\,
            I => \N__2702\
        );

    \I__617\ : ClkMux
    port map (
            O => \N__2757\,
            I => \N__2702\
        );

    \I__616\ : ClkMux
    port map (
            O => \N__2756\,
            I => \N__2702\
        );

    \I__615\ : ClkMux
    port map (
            O => \N__2755\,
            I => \N__2702\
        );

    \I__614\ : ClkMux
    port map (
            O => \N__2754\,
            I => \N__2702\
        );

    \I__613\ : ClkMux
    port map (
            O => \N__2753\,
            I => \N__2702\
        );

    \I__612\ : ClkMux
    port map (
            O => \N__2752\,
            I => \N__2702\
        );

    \I__611\ : ClkMux
    port map (
            O => \N__2751\,
            I => \N__2702\
        );

    \I__610\ : ClkMux
    port map (
            O => \N__2750\,
            I => \N__2702\
        );

    \I__609\ : ClkMux
    port map (
            O => \N__2749\,
            I => \N__2702\
        );

    \I__608\ : ClkMux
    port map (
            O => \N__2748\,
            I => \N__2702\
        );

    \I__607\ : ClkMux
    port map (
            O => \N__2747\,
            I => \N__2702\
        );

    \I__606\ : ClkMux
    port map (
            O => \N__2746\,
            I => \N__2702\
        );

    \I__605\ : ClkMux
    port map (
            O => \N__2745\,
            I => \N__2702\
        );

    \I__604\ : ClkMux
    port map (
            O => \N__2744\,
            I => \N__2702\
        );

    \I__603\ : ClkMux
    port map (
            O => \N__2743\,
            I => \N__2702\
        );

    \I__602\ : GlobalMux
    port map (
            O => \N__2702\,
            I => \N__2699\
        );

    \I__601\ : gio2CtrlBuf
    port map (
            O => \N__2699\,
            I => clk_system_c_g
        );

    \I__600\ : CEMux
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__598\ : Span4Mux_h
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__2687\,
            I => \uart.N_43_0\
        );

    \I__596\ : SRMux
    port map (
            O => \N__2684\,
            I => \N__2680\
        );

    \I__595\ : SRMux
    port map (
            O => \N__2683\,
            I => \N__2677\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__2680\,
            I => \N__2670\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__2677\,
            I => \N__2670\
        );

    \I__592\ : SRMux
    port map (
            O => \N__2676\,
            I => \N__2667\
        );

    \I__591\ : SRMux
    port map (
            O => \N__2675\,
            I => \N__2664\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__2670\,
            I => \N__2654\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__2667\,
            I => \N__2654\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2664\,
            I => \N__2651\
        );

    \I__587\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2640\
        );

    \I__586\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2640\
        );

    \I__585\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2635\
        );

    \I__584\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2635\
        );

    \I__583\ : SRMux
    port map (
            O => \N__2659\,
            I => \N__2632\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__2654\,
            I => \N__2627\
        );

    \I__581\ : Span4Mux_h
    port map (
            O => \N__2651\,
            I => \N__2627\
        );

    \I__580\ : SRMux
    port map (
            O => \N__2650\,
            I => \N__2624\
        );

    \I__579\ : SRMux
    port map (
            O => \N__2649\,
            I => \N__2621\
        );

    \I__578\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2616\
        );

    \I__577\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2616\
        );

    \I__576\ : SRMux
    port map (
            O => \N__2646\,
            I => \N__2611\
        );

    \I__575\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2611\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2640\,
            I => \N__2606\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__2635\,
            I => \N__2606\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__2632\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__2627\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__2624\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2621\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2616\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__2611\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__2606\,
            I => \uart.un1_state_4_0_a2_iso\
        );

    \I__565\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__2588\,
            I => \N__2582\
        );

    \I__563\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2577\
        );

    \I__562\ : InMux
    port map (
            O => \N__2586\,
            I => \N__2567\
        );

    \I__561\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2564\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__2582\,
            I => \N__2561\
        );

    \I__559\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2556\
        );

    \I__558\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2556\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__2577\,
            I => \N__2553\
        );

    \I__556\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2546\
        );

    \I__555\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2546\
        );

    \I__554\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2546\
        );

    \I__553\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2541\
        );

    \I__552\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2541\
        );

    \I__551\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2536\
        );

    \I__550\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2536\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2567\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2564\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__2561\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2556\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__2553\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2546\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2541\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__2536\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__2519\,
            I => \N__2514\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__2518\,
            I => \N__2511\
        );

    \I__539\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2503\
        );

    \I__538\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2503\
        );

    \I__537\ : InMux
    port map (
            O => \N__2511\,
            I => \N__2500\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__2510\,
            I => \N__2497\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__2509\,
            I => \N__2494\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__2508\,
            I => \N__2491\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2503\,
            I => \N__2485\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2500\,
            I => \N__2482\
        );

    \I__531\ : InMux
    port map (
            O => \N__2497\,
            I => \N__2479\
        );

    \I__530\ : InMux
    port map (
            O => \N__2494\,
            I => \N__2472\
        );

    \I__529\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2472\
        );

    \I__528\ : InMux
    port map (
            O => \N__2490\,
            I => \N__2472\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__2489\,
            I => \N__2469\
        );

    \I__526\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2465\
        );

    \I__525\ : Span4Mux_h
    port map (
            O => \N__2485\,
            I => \N__2462\
        );

    \I__524\ : Span4Mux_v
    port map (
            O => \N__2482\,
            I => \N__2455\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__2479\,
            I => \N__2455\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2472\,
            I => \N__2455\
        );

    \I__521\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2452\
        );

    \I__520\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2449\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2465\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__2462\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__2455\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__2452\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2449\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__2438\,
            I => \N__2430\
        );

    \I__513\ : InMux
    port map (
            O => \N__2437\,
            I => \N__2426\
        );

    \I__512\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2423\
        );

    \I__511\ : InMux
    port map (
            O => \N__2435\,
            I => \N__2418\
        );

    \I__510\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2418\
        );

    \I__509\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2415\
        );

    \I__508\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2410\
        );

    \I__507\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2410\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2426\,
            I => \uart.N_175\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__2423\,
            I => \uart.N_175\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2418\,
            I => \uart.N_175\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2415\,
            I => \uart.N_175\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2410\,
            I => \uart.N_175\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__2399\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_5_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__2396\,
            I => \N__2393\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2393\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_6\
        );

    \I__498\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2387\,
            I => \uart.state_1_sqmuxa\
        );

    \I__496\ : CEMux
    port map (
            O => \N__2384\,
            I => \N__2381\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__2381\,
            I => \uart.N_42_0\
        );

    \I__494\ : CEMux
    port map (
            O => \N__2378\,
            I => \N__2375\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2375\,
            I => \N__2372\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__2372\,
            I => \uart.N_41_0\
        );

    \I__491\ : CEMux
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2366\,
            I => \uart.N_37_0\
        );

    \I__489\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2360\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2360\,
            I => \uart.data_AuxZ0Z_0\
        );

    \I__487\ : IoInMux
    port map (
            O => \N__2357\,
            I => \N__2354\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2354\,
            I => \N__2351\
        );

    \I__485\ : Span12Mux_s5_v
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__484\ : Span12Mux_v
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__483\ : Odrv12
    port map (
            O => \N__2345\,
            I => data_c_0
        );

    \I__482\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2339\,
            I => \N__2336\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__479\ : Odrv4
    port map (
            O => \N__2333\,
            I => \uart.data_AuxZ0Z_1\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2324\
        );

    \I__476\ : IoSpan4Mux
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__475\ : Span4Mux_s3_v
    port map (
            O => \N__2321\,
            I => \N__2318\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__2318\,
            I => \N__2315\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__2315\,
            I => \N__2312\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__2312\,
            I => data_c_1
        );

    \I__471\ : IoInMux
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2306\,
            I => \N__2303\
        );

    \I__469\ : IoSpan4Mux
    port map (
            O => \N__2303\,
            I => \N__2300\
        );

    \I__468\ : Span4Mux_s3_v
    port map (
            O => \N__2300\,
            I => \N__2297\
        );

    \I__467\ : Sp12to4
    port map (
            O => \N__2297\,
            I => \N__2294\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__2294\,
            I => data_rdy_c
        );

    \I__465\ : InMux
    port map (
            O => \N__2291\,
            I => \N__2288\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2288\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_0\
        );

    \I__463\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2282\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2282\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_4\
        );

    \I__461\ : CEMux
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__2273\,
            I => \uart.N_39_0\
        );

    \I__458\ : CEMux
    port map (
            O => \N__2270\,
            I => \N__2267\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__2264\,
            I => \uart.N_40_0\
        );

    \I__455\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2258\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2258\,
            I => \uart.timer_Count_6_rep1_RNI1B4SZ0\
        );

    \I__453\ : InMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2252\,
            I => \uart.timer_Count_6_rep1_RNI02QZ0Z61\
        );

    \I__451\ : InMux
    port map (
            O => \N__2249\,
            I => \N__2245\
        );

    \I__450\ : InMux
    port map (
            O => \N__2248\,
            I => \N__2242\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2245\,
            I => \uart.N_145_0\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2242\,
            I => \uart.N_145_0\
        );

    \I__447\ : InMux
    port map (
            O => \N__2237\,
            I => \N__2232\
        );

    \I__446\ : InMux
    port map (
            O => \N__2236\,
            I => \N__2229\
        );

    \I__445\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2226\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2232\,
            I => \N__2223\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2229\,
            I => \N__2220\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2226\,
            I => \uart.timer_Count28\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__2223\,
            I => \uart.timer_Count28\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__2220\,
            I => \uart.timer_Count28\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__2213\,
            I => \uart.timer_Count28_cascade_\
        );

    \I__438\ : InMux
    port map (
            O => \N__2210\,
            I => \N__2206\
        );

    \I__437\ : InMux
    port map (
            O => \N__2209\,
            I => \N__2196\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2206\,
            I => \N__2193\
        );

    \I__435\ : InMux
    port map (
            O => \N__2205\,
            I => \N__2186\
        );

    \I__434\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2186\
        );

    \I__433\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2186\
        );

    \I__432\ : InMux
    port map (
            O => \N__2202\,
            I => \N__2179\
        );

    \I__431\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2179\
        );

    \I__430\ : InMux
    port map (
            O => \N__2200\,
            I => \N__2179\
        );

    \I__429\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2171\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2196\,
            I => \N__2168\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__2193\,
            I => \N__2161\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2186\,
            I => \N__2161\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2179\,
            I => \N__2161\
        );

    \I__424\ : InMux
    port map (
            O => \N__2178\,
            I => \N__2158\
        );

    \I__423\ : InMux
    port map (
            O => \N__2177\,
            I => \N__2155\
        );

    \I__422\ : InMux
    port map (
            O => \N__2176\,
            I => \N__2148\
        );

    \I__421\ : InMux
    port map (
            O => \N__2175\,
            I => \N__2148\
        );

    \I__420\ : InMux
    port map (
            O => \N__2174\,
            I => \N__2148\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2171\,
            I => \uart.stateZ0Z_4\
        );

    \I__418\ : Odrv12
    port map (
            O => \N__2168\,
            I => \uart.stateZ0Z_4\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__2161\,
            I => \uart.stateZ0Z_4\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2158\,
            I => \uart.stateZ0Z_4\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2155\,
            I => \uart.stateZ0Z_4\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2148\,
            I => \uart.stateZ0Z_4\
        );

    \I__413\ : InMux
    port map (
            O => \N__2135\,
            I => \N__2127\
        );

    \I__412\ : InMux
    port map (
            O => \N__2134\,
            I => \N__2124\
        );

    \I__411\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2117\
        );

    \I__410\ : InMux
    port map (
            O => \N__2132\,
            I => \N__2117\
        );

    \I__409\ : InMux
    port map (
            O => \N__2131\,
            I => \N__2117\
        );

    \I__408\ : InMux
    port map (
            O => \N__2130\,
            I => \N__2111\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2127\,
            I => \N__2104\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2124\,
            I => \N__2104\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2117\,
            I => \N__2104\
        );

    \I__404\ : InMux
    port map (
            O => \N__2116\,
            I => \N__2099\
        );

    \I__403\ : InMux
    port map (
            O => \N__2115\,
            I => \N__2099\
        );

    \I__402\ : InMux
    port map (
            O => \N__2114\,
            I => \N__2093\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2111\,
            I => \N__2086\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__2104\,
            I => \N__2086\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2099\,
            I => \N__2086\
        );

    \I__398\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2081\
        );

    \I__397\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2081\
        );

    \I__396\ : InMux
    port map (
            O => \N__2096\,
            I => \N__2078\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2093\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__394\ : Odrv4
    port map (
            O => \N__2086\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2081\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2078\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__2069\,
            I => \N__2065\
        );

    \I__390\ : InMux
    port map (
            O => \N__2068\,
            I => \N__2057\
        );

    \I__389\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2057\
        );

    \I__388\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2057\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2057\,
            I => \uart.un4_timer_Count_1_c2\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__2054\,
            I => \uart.timer_Count_RNIMLMA1Z0Z_1_cascade_\
        );

    \I__385\ : InMux
    port map (
            O => \N__2051\,
            I => \N__2039\
        );

    \I__384\ : InMux
    port map (
            O => \N__2050\,
            I => \N__2039\
        );

    \I__383\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2039\
        );

    \I__382\ : InMux
    port map (
            O => \N__2048\,
            I => \N__2039\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2039\,
            I => \uart.un4_timer_Count_1_c5\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__2036\,
            I => \uart.un4_timer_Count_1_c5_cascade_\
        );

    \I__379\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2028\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2032\,
            I => \N__2024\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__2031\,
            I => \N__2019\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2028\,
            I => \N__2014\
        );

    \I__375\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2009\
        );

    \I__374\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2009\
        );

    \I__373\ : InMux
    port map (
            O => \N__2023\,
            I => \N__2006\
        );

    \I__372\ : InMux
    port map (
            O => \N__2022\,
            I => \N__2003\
        );

    \I__371\ : InMux
    port map (
            O => \N__2019\,
            I => \N__1996\
        );

    \I__370\ : InMux
    port map (
            O => \N__2018\,
            I => \N__1996\
        );

    \I__369\ : InMux
    port map (
            O => \N__2017\,
            I => \N__1996\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__2014\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2009\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2006\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2003\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__1996\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__363\ : InMux
    port map (
            O => \N__1985\,
            I => \N__1982\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__1982\,
            I => \N__1971\
        );

    \I__361\ : InMux
    port map (
            O => \N__1981\,
            I => \N__1966\
        );

    \I__360\ : InMux
    port map (
            O => \N__1980\,
            I => \N__1966\
        );

    \I__359\ : InMux
    port map (
            O => \N__1979\,
            I => \N__1963\
        );

    \I__358\ : InMux
    port map (
            O => \N__1978\,
            I => \N__1960\
        );

    \I__357\ : InMux
    port map (
            O => \N__1977\,
            I => \N__1951\
        );

    \I__356\ : InMux
    port map (
            O => \N__1976\,
            I => \N__1951\
        );

    \I__355\ : InMux
    port map (
            O => \N__1975\,
            I => \N__1951\
        );

    \I__354\ : InMux
    port map (
            O => \N__1974\,
            I => \N__1951\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__1971\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__1966\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__1963\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__1960\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1951\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__1940\,
            I => \N__1928\
        );

    \I__347\ : InMux
    port map (
            O => \N__1939\,
            I => \N__1924\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__1938\,
            I => \N__1920\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__1937\,
            I => \N__1917\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__1936\,
            I => \N__1914\
        );

    \I__343\ : InMux
    port map (
            O => \N__1935\,
            I => \N__1911\
        );

    \I__342\ : InMux
    port map (
            O => \N__1934\,
            I => \N__1904\
        );

    \I__341\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1904\
        );

    \I__340\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1904\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__1931\,
            I => \N__1901\
        );

    \I__338\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1897\
        );

    \I__337\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1894\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1924\,
            I => \N__1891\
        );

    \I__335\ : InMux
    port map (
            O => \N__1923\,
            I => \N__1884\
        );

    \I__334\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1884\
        );

    \I__333\ : InMux
    port map (
            O => \N__1917\,
            I => \N__1884\
        );

    \I__332\ : InMux
    port map (
            O => \N__1914\,
            I => \N__1881\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1911\,
            I => \N__1876\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__1904\,
            I => \N__1876\
        );

    \I__329\ : InMux
    port map (
            O => \N__1901\,
            I => \N__1871\
        );

    \I__328\ : InMux
    port map (
            O => \N__1900\,
            I => \N__1871\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__1897\,
            I => \uart.stateZ0Z_3\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1894\,
            I => \uart.stateZ0Z_3\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__1891\,
            I => \uart.stateZ0Z_3\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1884\,
            I => \uart.stateZ0Z_3\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1881\,
            I => \uart.stateZ0Z_3\
        );

    \I__322\ : Odrv4
    port map (
            O => \N__1876\,
            I => \uart.stateZ0Z_3\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__1871\,
            I => \uart.stateZ0Z_3\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__1856\,
            I => \uart.timer_Count_RNIHJ661Z0Z_3_cascade_\
        );

    \I__319\ : InMux
    port map (
            O => \N__1853\,
            I => \N__1847\
        );

    \I__318\ : InMux
    port map (
            O => \N__1852\,
            I => \N__1847\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1847\,
            I => \N__1839\
        );

    \I__316\ : InMux
    port map (
            O => \N__1846\,
            I => \N__1833\
        );

    \I__315\ : InMux
    port map (
            O => \N__1845\,
            I => \N__1819\
        );

    \I__314\ : InMux
    port map (
            O => \N__1844\,
            I => \N__1819\
        );

    \I__313\ : InMux
    port map (
            O => \N__1843\,
            I => \N__1819\
        );

    \I__312\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1819\
        );

    \I__311\ : Span4Mux_h
    port map (
            O => \N__1839\,
            I => \N__1816\
        );

    \I__310\ : InMux
    port map (
            O => \N__1838\,
            I => \N__1809\
        );

    \I__309\ : InMux
    port map (
            O => \N__1837\,
            I => \N__1809\
        );

    \I__308\ : InMux
    port map (
            O => \N__1836\,
            I => \N__1809\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1833\,
            I => \N__1806\
        );

    \I__306\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1799\
        );

    \I__305\ : InMux
    port map (
            O => \N__1831\,
            I => \N__1799\
        );

    \I__304\ : InMux
    port map (
            O => \N__1830\,
            I => \N__1799\
        );

    \I__303\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1794\
        );

    \I__302\ : InMux
    port map (
            O => \N__1828\,
            I => \N__1794\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1819\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__300\ : Odrv4
    port map (
            O => \N__1816\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1809\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__298\ : Odrv4
    port map (
            O => \N__1806\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1799\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1794\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__295\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1776\
        );

    \I__294\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1773\
        );

    \I__293\ : InMux
    port map (
            O => \N__1779\,
            I => \N__1770\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1776\,
            I => \N__1767\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1773\,
            I => \N__1762\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1770\,
            I => \N__1762\
        );

    \I__289\ : Span4Mux_h
    port map (
            O => \N__1767\,
            I => \N__1759\
        );

    \I__288\ : Span4Mux_v
    port map (
            O => \N__1762\,
            I => \N__1756\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__1759\,
            I => \uart.state_0_sqmuxa_1_d\
        );

    \I__286\ : Odrv4
    port map (
            O => \N__1756\,
            I => \uart.state_0_sqmuxa_1_d\
        );

    \I__285\ : InMux
    port map (
            O => \N__1751\,
            I => \N__1744\
        );

    \I__284\ : InMux
    port map (
            O => \N__1750\,
            I => \N__1739\
        );

    \I__283\ : InMux
    port map (
            O => \N__1749\,
            I => \N__1739\
        );

    \I__282\ : InMux
    port map (
            O => \N__1748\,
            I => \N__1734\
        );

    \I__281\ : InMux
    port map (
            O => \N__1747\,
            I => \N__1734\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1744\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1739\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1734\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__277\ : InMux
    port map (
            O => \N__1727\,
            I => \N__1718\
        );

    \I__276\ : InMux
    port map (
            O => \N__1726\,
            I => \N__1718\
        );

    \I__275\ : InMux
    port map (
            O => \N__1725\,
            I => \N__1713\
        );

    \I__274\ : InMux
    port map (
            O => \N__1724\,
            I => \N__1713\
        );

    \I__273\ : InMux
    port map (
            O => \N__1723\,
            I => \N__1710\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1718\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1713\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1710\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__269\ : SRMux
    port map (
            O => \N__1703\,
            I => \N__1699\
        );

    \I__268\ : SRMux
    port map (
            O => \N__1702\,
            I => \N__1696\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1699\,
            I => \N__1693\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1696\,
            I => \N__1689\
        );

    \I__265\ : Span4Mux_h
    port map (
            O => \N__1693\,
            I => \N__1686\
        );

    \I__264\ : SRMux
    port map (
            O => \N__1692\,
            I => \N__1683\
        );

    \I__263\ : Span4Mux_v
    port map (
            O => \N__1689\,
            I => \N__1680\
        );

    \I__262\ : Sp12to4
    port map (
            O => \N__1686\,
            I => \N__1675\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1683\,
            I => \N__1675\
        );

    \I__260\ : Odrv4
    port map (
            O => \N__1680\,
            I => \uart.un1_timer_Count_0_sqmuxa_0\
        );

    \I__259\ : Odrv12
    port map (
            O => \N__1675\,
            I => \uart.un1_timer_Count_0_sqmuxa_0\
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__1670\,
            I => \N__1667\
        );

    \I__257\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1661\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__1666\,
            I => \N__1654\
        );

    \I__255\ : CascadeMux
    port map (
            O => \N__1665\,
            I => \N__1651\
        );

    \I__254\ : InMux
    port map (
            O => \N__1664\,
            I => \N__1648\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1661\,
            I => \N__1645\
        );

    \I__252\ : InMux
    port map (
            O => \N__1660\,
            I => \N__1638\
        );

    \I__251\ : InMux
    port map (
            O => \N__1659\,
            I => \N__1638\
        );

    \I__250\ : InMux
    port map (
            O => \N__1658\,
            I => \N__1638\
        );

    \I__249\ : InMux
    port map (
            O => \N__1657\,
            I => \N__1635\
        );

    \I__248\ : InMux
    port map (
            O => \N__1654\,
            I => \N__1632\
        );

    \I__247\ : InMux
    port map (
            O => \N__1651\,
            I => \N__1629\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1648\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__245\ : Odrv12
    port map (
            O => \N__1645\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1638\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1635\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1632\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1629\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__1616\,
            I => \N__1612\
        );

    \I__239\ : InMux
    port map (
            O => \N__1615\,
            I => \N__1599\
        );

    \I__238\ : InMux
    port map (
            O => \N__1612\,
            I => \N__1599\
        );

    \I__237\ : InMux
    port map (
            O => \N__1611\,
            I => \N__1592\
        );

    \I__236\ : InMux
    port map (
            O => \N__1610\,
            I => \N__1592\
        );

    \I__235\ : InMux
    port map (
            O => \N__1609\,
            I => \N__1592\
        );

    \I__234\ : InMux
    port map (
            O => \N__1608\,
            I => \N__1585\
        );

    \I__233\ : InMux
    port map (
            O => \N__1607\,
            I => \N__1582\
        );

    \I__232\ : InMux
    port map (
            O => \N__1606\,
            I => \N__1575\
        );

    \I__231\ : InMux
    port map (
            O => \N__1605\,
            I => \N__1575\
        );

    \I__230\ : InMux
    port map (
            O => \N__1604\,
            I => \N__1575\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__1599\,
            I => \N__1570\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1592\,
            I => \N__1570\
        );

    \I__227\ : InMux
    port map (
            O => \N__1591\,
            I => \N__1565\
        );

    \I__226\ : InMux
    port map (
            O => \N__1590\,
            I => \N__1565\
        );

    \I__225\ : InMux
    port map (
            O => \N__1589\,
            I => \N__1560\
        );

    \I__224\ : InMux
    port map (
            O => \N__1588\,
            I => \N__1560\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1585\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1582\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1575\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__220\ : Odrv4
    port map (
            O => \N__1570\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1565\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1560\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__1547\,
            I => \N__1544\
        );

    \I__216\ : InMux
    port map (
            O => \N__1544\,
            I => \N__1541\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1541\,
            I => \uart.N_28_mux_i_i_0\
        );

    \I__214\ : InMux
    port map (
            O => \N__1538\,
            I => \N__1535\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1535\,
            I => \uart.N_22_mux\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__1532\,
            I => \uart.N_175_cascade_\
        );

    \I__211\ : InMux
    port map (
            O => \N__1529\,
            I => \N__1526\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1526\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_1\
        );

    \I__209\ : CascadeMux
    port map (
            O => \N__1523\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__1520\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__207\ : InMux
    port map (
            O => \N__1517\,
            I => \N__1512\
        );

    \I__206\ : InMux
    port map (
            O => \N__1516\,
            I => \N__1509\
        );

    \I__205\ : InMux
    port map (
            O => \N__1515\,
            I => \N__1503\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1512\,
            I => \N__1500\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1509\,
            I => \N__1497\
        );

    \I__202\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1494\
        );

    \I__201\ : InMux
    port map (
            O => \N__1507\,
            I => \N__1489\
        );

    \I__200\ : InMux
    port map (
            O => \N__1506\,
            I => \N__1489\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1503\,
            I => \uart.timer_Count_6_repZ0Z1\
        );

    \I__198\ : Odrv4
    port map (
            O => \N__1500\,
            I => \uart.timer_Count_6_repZ0Z1\
        );

    \I__197\ : Odrv4
    port map (
            O => \N__1497\,
            I => \uart.timer_Count_6_repZ0Z1\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1494\,
            I => \uart.timer_Count_6_repZ0Z1\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1489\,
            I => \uart.timer_Count_6_repZ0Z1\
        );

    \I__194\ : CascadeMux
    port map (
            O => \N__1478\,
            I => \N__1473\
        );

    \I__193\ : InMux
    port map (
            O => \N__1477\,
            I => \N__1470\
        );

    \I__192\ : InMux
    port map (
            O => \N__1476\,
            I => \N__1467\
        );

    \I__191\ : InMux
    port map (
            O => \N__1473\,
            I => \N__1464\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1470\,
            I => \uart.timer_Count_fastZ0Z_6\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1467\,
            I => \uart.timer_Count_fastZ0Z_6\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1464\,
            I => \uart.timer_Count_fastZ0Z_6\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__1457\,
            I => \uart.un1_state_4_0_a2_iso_cascade_\
        );

    \I__186\ : CEMux
    port map (
            O => \N__1454\,
            I => \N__1451\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1451\,
            I => \N__1448\
        );

    \I__184\ : Span4Mux_h
    port map (
            O => \N__1448\,
            I => \N__1445\
        );

    \I__183\ : Odrv4
    port map (
            O => \N__1445\,
            I => \uart.N_38_0\
        );

    \I__182\ : InMux
    port map (
            O => \N__1442\,
            I => \N__1438\
        );

    \I__181\ : InMux
    port map (
            O => \N__1441\,
            I => \N__1435\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1438\,
            I => \uart.N_165_1\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1435\,
            I => \uart.N_165_1\
        );

    \I__178\ : InMux
    port map (
            O => \N__1430\,
            I => \N__1427\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1427\,
            I => \uart.timer_Count_RNIICSG1Z0Z_6\
        );

    \I__176\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1421\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1421\,
            I => \uart.state_RNO_0Z0Z_3\
        );

    \I__174\ : CascadeMux
    port map (
            O => \N__1418\,
            I => \N__1415\
        );

    \I__173\ : InMux
    port map (
            O => \N__1415\,
            I => \N__1412\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1412\,
            I => \N__1409\
        );

    \I__171\ : Odrv4
    port map (
            O => \N__1409\,
            I => \uart.state_RNO_1Z0Z_3\
        );

    \I__170\ : CascadeMux
    port map (
            O => \N__1406\,
            I => \N__1403\
        );

    \I__169\ : InMux
    port map (
            O => \N__1403\,
            I => \N__1399\
        );

    \I__168\ : InMux
    port map (
            O => \N__1402\,
            I => \N__1396\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1399\,
            I => \N__1393\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1396\,
            I => \uart.N_147_0\
        );

    \I__165\ : Odrv4
    port map (
            O => \N__1393\,
            I => \uart.N_147_0\
        );

    \I__164\ : InMux
    port map (
            O => \N__1388\,
            I => \N__1385\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1385\,
            I => \N__1382\
        );

    \I__162\ : Odrv4
    port map (
            O => \N__1382\,
            I => \uart.N_159\
        );

    \I__161\ : CascadeMux
    port map (
            O => \N__1379\,
            I => \uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_\
        );

    \I__160\ : CascadeMux
    port map (
            O => \N__1376\,
            I => \uart.un1_state_2_0_a3_0_cascade_\
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__1373\,
            I => \N__1367\
        );

    \I__158\ : InMux
    port map (
            O => \N__1372\,
            I => \N__1361\
        );

    \I__157\ : InMux
    port map (
            O => \N__1371\,
            I => \N__1356\
        );

    \I__156\ : InMux
    port map (
            O => \N__1370\,
            I => \N__1356\
        );

    \I__155\ : InMux
    port map (
            O => \N__1367\,
            I => \N__1350\
        );

    \I__154\ : InMux
    port map (
            O => \N__1366\,
            I => \N__1350\
        );

    \I__153\ : InMux
    port map (
            O => \N__1365\,
            I => \N__1345\
        );

    \I__152\ : InMux
    port map (
            O => \N__1364\,
            I => \N__1345\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__1361\,
            I => \N__1340\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1356\,
            I => \N__1340\
        );

    \I__149\ : InMux
    port map (
            O => \N__1355\,
            I => \N__1337\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1350\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1345\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__146\ : Odrv4
    port map (
            O => \N__1340\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1337\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__144\ : CEMux
    port map (
            O => \N__1328\,
            I => \N__1325\
        );

    \I__143\ : LocalMux
    port map (
            O => \N__1325\,
            I => \N__1322\
        );

    \I__142\ : Odrv4
    port map (
            O => \N__1322\,
            I => \uart.N_44_0\
        );

    \I__141\ : CascadeMux
    port map (
            O => \N__1319\,
            I => \uart.N_147_0_cascade_\
        );

    \I__140\ : InMux
    port map (
            O => \N__1316\,
            I => \N__1313\
        );

    \I__139\ : LocalMux
    port map (
            O => \N__1313\,
            I => \uart.timer_Count_RNITC202Z0Z_6\
        );

    \I__138\ : CascadeMux
    port map (
            O => \N__1310\,
            I => \uart.timer_Count_RNIGLM11Z0Z_6_cascade_\
        );

    \I__137\ : InMux
    port map (
            O => \N__1307\,
            I => \N__1303\
        );

    \I__136\ : InMux
    port map (
            O => \N__1306\,
            I => \N__1300\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1303\,
            I => \uart.un1_state_7_0_0\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1300\,
            I => \uart.un1_state_7_0_0\
        );

    \I__133\ : CascadeMux
    port map (
            O => \N__1295\,
            I => \uart.un1_state_7_0_0_cascade_\
        );

    \I__132\ : InMux
    port map (
            O => \N__1292\,
            I => \N__1286\
        );

    \I__131\ : InMux
    port map (
            O => \N__1291\,
            I => \N__1286\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1286\,
            I => \uart.N_177\
        );

    \I__129\ : InMux
    port map (
            O => \N__1283\,
            I => \N__1280\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__1280\,
            I => \N__1277\
        );

    \I__127\ : Odrv4
    port map (
            O => \N__1277\,
            I => \uart.un1_state_5\
        );

    \I__126\ : CascadeMux
    port map (
            O => \N__1274\,
            I => \uart.state_RNO_1Z0Z_2_cascade_\
        );

    \I__125\ : InMux
    port map (
            O => \N__1271\,
            I => \N__1268\
        );

    \I__124\ : LocalMux
    port map (
            O => \N__1268\,
            I => \uart.state_RNO_2Z0Z_2\
        );

    \I__123\ : CascadeMux
    port map (
            O => \N__1265\,
            I => \uart.N_170_cascade_\
        );

    \I__122\ : CascadeMux
    port map (
            O => \N__1262\,
            I => \N__1257\
        );

    \I__121\ : CascadeMux
    port map (
            O => \N__1261\,
            I => \N__1254\
        );

    \I__120\ : InMux
    port map (
            O => \N__1260\,
            I => \N__1244\
        );

    \I__119\ : InMux
    port map (
            O => \N__1257\,
            I => \N__1244\
        );

    \I__118\ : InMux
    port map (
            O => \N__1254\,
            I => \N__1244\
        );

    \I__117\ : InMux
    port map (
            O => \N__1253\,
            I => \N__1244\
        );

    \I__116\ : LocalMux
    port map (
            O => \N__1244\,
            I => \uart.stateZ0Z_2\
        );

    \I__115\ : CascadeMux
    port map (
            O => \N__1241\,
            I => \N__1237\
        );

    \I__114\ : InMux
    port map (
            O => \N__1240\,
            I => \N__1229\
        );

    \I__113\ : InMux
    port map (
            O => \N__1237\,
            I => \N__1229\
        );

    \I__112\ : InMux
    port map (
            O => \N__1236\,
            I => \N__1229\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1229\,
            I => \uart.stateZ0Z_1\
        );

    \I__110\ : CascadeMux
    port map (
            O => \N__1226\,
            I => \uart.data_Aux_esr_RNO_0Z0Z_7_cascade_\
        );

    \I__109\ : CascadeMux
    port map (
            O => \N__1223\,
            I => \uart.CO0_0_cascade_\
        );

    \I__108\ : CascadeMux
    port map (
            O => \N__1220\,
            I => \uart.bit_Count_RNO_1Z0Z_2_cascade_\
        );

    \I__107\ : CascadeMux
    port map (
            O => \N__1217\,
            I => \uart.CO1_1_cascade_\
        );

    \I__106\ : InMux
    port map (
            O => \N__1214\,
            I => \N__1211\
        );

    \I__105\ : LocalMux
    port map (
            O => \N__1211\,
            I => \uart.bit_Count_RNO_2Z0Z_2\
        );

    \I__104\ : InMux
    port map (
            O => \N__1208\,
            I => \N__1205\
        );

    \I__103\ : LocalMux
    port map (
            O => \N__1205\,
            I => \uart.bit_Count_RNO_1Z0Z_1\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart.bit_Count_RNO_0_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1208\,
            in2 => \_gnd_net_\,
            in3 => \N__2586\,
            lcout => OPEN,
            ltout => \uart.CO0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_1_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__1779\,
            in1 => \N__1307\,
            in2 => \N__1223\,
            in3 => \N__2114\,
            lcout => \uart.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_1_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2202\,
            in1 => \N__2098\,
            in2 => \N__1931\,
            in3 => \N__2573\,
            lcout => OPEN,
            ltout => \uart.bit_Count_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_0_2_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__1615\,
            in1 => \N__1214\,
            in2 => \N__1220\,
            in3 => \N__1517\,
            lcout => OPEN,
            ltout => \uart.CO1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_2_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__1780\,
            in1 => \N__1306\,
            in2 => \N__1217\,
            in3 => \N__2488\,
            lcout => \uart.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_2_2_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__2200\,
            in1 => \N__2097\,
            in2 => \_gnd_net_\,
            in3 => \N__2572\,
            lcout => \uart.bit_Count_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_1_1_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110011"
        )
    port map (
            in0 => \N__1372\,
            in1 => \N__1900\,
            in2 => \N__1616\,
            in3 => \N__2201\,
            lcout => \uart.bit_Count_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_1_3_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__1933\,
            in1 => \N__1476\,
            in2 => \N__1261\,
            in3 => \N__1606\,
            lcout => \uart.state_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIB0BC_2_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1253\,
            in2 => \_gnd_net_\,
            in3 => \N__1932\,
            lcout => \uart.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_2_2_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__1364\,
            in1 => \N__1236\,
            in2 => \_gnd_net_\,
            in3 => \N__1604\,
            lcout => \uart.state_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_1_2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__1605\,
            in1 => \N__1365\,
            in2 => \N__1241\,
            in3 => \N__1853\,
            lcout => OPEN,
            ltout => \uart.state_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_2_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1402\,
            in2 => \N__1274\,
            in3 => \N__1271\,
            lcout => OPEN,
            ltout => \uart.N_170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_2_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__1240\,
            in1 => \N__2902\,
            in2 => \N__1265\,
            in3 => \N__1260\,
            lcout => \uart.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_1_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__1934\,
            in1 => \N__2901\,
            in2 => \N__1262\,
            in3 => \N__2210\,
            lcout => \uart.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_3_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__2033\,
            in1 => \N__1985\,
            in2 => \N__1670\,
            in3 => \N__1852\,
            lcout => \uart.state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_7_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2130\,
            in1 => \N__2585\,
            in2 => \N__2489\,
            in3 => \N__2437\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_7_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1226\,
            in3 => \N__2645\,
            lcout => \uart.N_44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_7_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2753\,
            ce => \N__1328\,
            sr => \N__2646\
        );

    \uart.timer_Count_RNIBAKE2_6_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1291\,
            in2 => \_gnd_net_\,
            in3 => \N__1316\,
            lcout => \uart.N_165_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIQ1101_3_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2022\,
            in1 => \N__1978\,
            in2 => \_gnd_net_\,
            in3 => \N__1657\,
            lcout => \uart.N_147_0\,
            ltout => \uart.N_147_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNITC202_6_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__1609\,
            in1 => \N__1370\,
            in2 => \N__1319\,
            in3 => \N__1846\,
            lcout => \uart.timer_Count_RNITC202Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIGLM11_6_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__1371\,
            in1 => \N__1610\,
            in2 => \N__1937\,
            in3 => \N__2203\,
            lcout => OPEN,
            ltout => \uart.timer_Count_RNIGLM11Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIBLJS1_3_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__2204\,
            in1 => \N__1923\,
            in2 => \N__1310\,
            in3 => \N__1292\,
            lcout => \uart.un1_state_7_0_0\,
            ltout => \uart.un1_state_7_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_0_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011000101010"
        )
    port map (
            in0 => \N__2571\,
            in1 => \N__1781\,
            in2 => \N__1295\,
            in3 => \N__1283\,
            lcout => \uart.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNIETHE_2_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2096\,
            in1 => \N__2468\,
            in2 => \_gnd_net_\,
            in3 => \N__2570\,
            lcout => \uart.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNO_0_0_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__1516\,
            in1 => \N__1611\,
            in2 => \N__1938\,
            in3 => \N__2205\,
            lcout => \uart.un1_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNINU001_0_1_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2023\,
            in1 => \N__1979\,
            in2 => \_gnd_net_\,
            in3 => \N__1724\,
            lcout => \uart.N_22_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_3_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100000101"
        )
    port map (
            in0 => \N__1424\,
            in1 => \N__1441\,
            in2 => \N__1418\,
            in3 => \N__1935\,
            lcout => \uart.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_6_rep1_RNIRC5S1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__1832\,
            in1 => \N__1508\,
            in2 => \N__1406\,
            in3 => \N__1591\,
            lcout => OPEN,
            ltout => \uart.timer_Count_6_rep1_RNIRC5SZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNILALH5_4_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__1388\,
            in1 => \N__2236\,
            in2 => \N__1379\,
            in3 => \N__2176\,
            lcout => \uart.un1_timer_Count_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIQ9BL_0_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1665\,
            in3 => \N__1747\,
            lcout => OPEN,
            ltout => \uart.un1_state_2_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIICSG1_6_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1355\,
            in1 => \N__2174\,
            in2 => \N__1376\,
            in3 => \N__1830\,
            lcout => \uart.timer_Count_RNIICSG1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIN6BL_0_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1725\,
            in2 => \_gnd_net_\,
            in3 => \N__1748\,
            lcout => \uart.un4_timer_Count_1_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_fast_RNI7MEA1_6_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111111111"
        )
    port map (
            in0 => \N__1590\,
            in1 => \N__1831\,
            in2 => \N__1478\,
            in3 => \N__2175\,
            lcout => \uart.N_28_mux_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_7_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__1842\,
            in1 => \N__2051\,
            in2 => \N__1373\,
            in3 => \N__1608\,
            lcout => \uart.timer_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2744\,
            ce => 'H',
            sr => \N__1692\
        );

    \uart.timer_Count_6_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2048\,
            in1 => \N__1366\,
            in2 => \_gnd_net_\,
            in3 => \N__1844\,
            lcout => \uart.timer_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2744\,
            ce => 'H',
            sr => \N__1692\
        );

    \uart.timer_Count_fast_6_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__1843\,
            in1 => \N__2050\,
            in2 => \_gnd_net_\,
            in3 => \N__1477\,
            lcout => \uart.timer_Count_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2744\,
            ce => 'H',
            sr => \N__1692\
        );

    \uart.timer_Count_6_rep1_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2049\,
            in1 => \N__1515\,
            in2 => \_gnd_net_\,
            in3 => \N__1845\,
            lcout => \uart.timer_Count_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2744\,
            ce => 'H',
            sr => \N__1692\
        );

    \uart.timer_Count_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1751\,
            lcout => \uart.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2744\,
            ce => 'H',
            sr => \N__1692\
        );

    \uart.data_Aux_esr_1_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2758\,
            ce => \N__1454\,
            sr => \N__2649\
        );

    \uart.data_Aux_esr_RNO_0_4_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2581\,
            in1 => \N__2517\,
            in2 => \N__2438\,
            in3 => \N__2116\,
            lcout => \uart.data_Aux_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_0_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__2115\,
            in1 => \N__2580\,
            in2 => \N__2519\,
            in3 => \N__2429\,
            lcout => \uart.data_Aux_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNID2BC_3_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1939\,
            in2 => \_gnd_net_\,
            in3 => \N__2177\,
            lcout => \uart.un1_state_4_0_a2_iso\,
            ltout => \uart.un1_state_4_0_a2_iso_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_1_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1457\,
            in3 => \N__1529\,
            lcout => \uart.N_38_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_4_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__2235\,
            in1 => \N__1442\,
            in2 => \N__1940\,
            in3 => \N__2199\,
            lcout => \uart.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNI9BTG2_6_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2248\,
            in2 => \_gnd_net_\,
            in3 => \N__1430\,
            lcout => \uart.N_175\,
            ltout => \uart.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_1_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2131\,
            in1 => \N__2490\,
            in2 => \N__1532\,
            in3 => \N__2574\,
            lcout => \uart.data_Aux_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_3_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2576\,
            in1 => \N__2133\,
            in2 => \N__2509\,
            in3 => \N__2435\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_3_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1523\,
            in3 => \N__2661\,
            lcout => \uart.N_40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_2_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2575\,
            in1 => \N__2132\,
            in2 => \N__2508\,
            in3 => \N__2434\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_2_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1520\,
            in3 => \N__2660\,
            lcout => \uart.N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_4_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1664\,
            in1 => \N__2068\,
            in2 => \N__2031\,
            in3 => \N__1977\,
            lcout => \uart.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2751\,
            ce => 'H',
            sr => \N__1703\
        );

    \uart.timer_Count_6_rep1_RNI1B4S_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__1589\,
            in1 => \N__1506\,
            in2 => \_gnd_net_\,
            in3 => \N__1828\,
            lcout => \uart.timer_Count_6_rep1_RNI1B4SZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_6_rep1_RNI02Q61_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__1588\,
            in1 => \N__1507\,
            in2 => \N__1666\,
            in3 => \N__1829\,
            lcout => \uart.timer_Count_6_rep1_RNI02QZ0Z61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNINU001_1_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2017\,
            in1 => \N__1974\,
            in2 => \_gnd_net_\,
            in3 => \N__1723\,
            lcout => \uart.N_145_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_3_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__1976\,
            in1 => \_gnd_net_\,
            in2 => \N__2069\,
            in3 => \N__2018\,
            lcout => \uart.timer_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2751\,
            ce => 'H',
            sr => \N__1703\
        );

    \uart.timer_Count_2_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2064\,
            in2 => \_gnd_net_\,
            in3 => \N__1975\,
            lcout => \uart.timer_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2751\,
            ce => 'H',
            sr => \N__1703\
        );

    \uart.timer_Count_RNIMLMA1_1_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1980\,
            in1 => \N__1660\,
            in2 => \N__2032\,
            in3 => \N__1726\,
            lcout => OPEN,
            ltout => \uart.timer_Count_RNIMLMA1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIH8CL1_0_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2054\,
            in3 => \N__1749\,
            lcout => \uart.un4_timer_Count_1_c5\,
            ltout => \uart.un4_timer_Count_1_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_5_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2036\,
            in3 => \N__1838\,
            lcout => \uart.timer_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2748\,
            ce => 'H',
            sr => \N__1702\
        );

    \uart.timer_Count_RNIHJ661_3_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__1836\,
            in1 => \N__2027\,
            in2 => \N__1936\,
            in3 => \N__1981\,
            lcout => OPEN,
            ltout => \uart.timer_Count_RNIHJ661Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNI6JN12_4_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111010001"
        )
    port map (
            in0 => \N__1927\,
            in1 => \N__1659\,
            in2 => \N__1856\,
            in3 => \N__1837\,
            lcout => \uart.state_0_sqmuxa_1_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_1_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__1727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1750\,
            lcout => \uart.timer_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2748\,
            ce => 'H',
            sr => \N__1702\
        );

    \uart.timer_Count_RNIV5RV2_4_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__1658\,
            in1 => \N__1607\,
            in2 => \N__1547\,
            in3 => \N__1538\,
            lcout => \uart.state_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_rdy_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__2866\,
            in1 => \N__2237\,
            in2 => \_gnd_net_\,
            in3 => \N__2209\,
            lcout => data_rdy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2647\,
            in2 => \_gnd_net_\,
            in3 => \N__2291\,
            lcout => \uart.N_37_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_4_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__2648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2285\,
            lcout => \uart.N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2759\,
            ce => \N__2279\,
            sr => \N__2650\
        );

    \uart.data_Aux_esr_3_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2756\,
            ce => \N__2270\,
            sr => \N__2659\
        );

    \uart.data_Aux_esr_RNO_0_6_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2134\,
            in1 => \N__2587\,
            in2 => \N__2510\,
            in3 => \N__2433\,
            lcout => \uart.data_Aux_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_6_rep1_RNIOBV23_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__2261\,
            in1 => \N__2255\,
            in2 => \_gnd_net_\,
            in3 => \N__2249\,
            lcout => \uart.timer_Count28\,
            ltout => \uart.timer_Count28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIVF8I3_4_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__2909\,
            in1 => \_gnd_net_\,
            in2 => \N__2213\,
            in3 => \N__2178\,
            lcout => \uart.state_RNIVF8I3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_0_5_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2135\,
            in1 => \N__2591\,
            in2 => \N__2518\,
            in3 => \N__2436\,
            lcout => OPEN,
            ltout => \uart.data_Aux_esr_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_5_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2399\,
            in3 => \N__2662\,
            lcout => \uart.N_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_RNO_6_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__2663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2396\,
            lcout => \uart.N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIUL3I6_4_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2390\,
            in2 => \_gnd_net_\,
            in3 => \N__2922\,
            lcout => \uart.state_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_esr_5_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2907\,
            lcout => \uart.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2752\,
            ce => \N__2384\,
            sr => \N__2683\
        );

    \uart.data_Aux_esr_4_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2762\,
            ce => \N__2378\,
            sr => \N__2676\
        );

    \uart.data_Aux_esr_0_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2761\,
            ce => \N__2369\,
            sr => \N__2675\
        );

    \uart.data_esr_0_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2363\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => data_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => data_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_2_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3113\,
            lcout => data_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_3_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3086\,
            lcout => data_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_5_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3056\,
            lcout => data_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_6_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => data_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_7_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3011\,
            lcout => data_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2760\,
            ce => \N__2954\,
            sr => \N__2936\
        );

    \uart.data_esr_4_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2981\,
            lcout => data_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2757\,
            ce => \N__2953\,
            sr => \N__2929\
        );

    \uart.data_Aux_esr_6_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2755\,
            ce => \N__2696\,
            sr => \N__2684\
        );
end \INTERFACE\;
